module fake_jpeg_2827_n_442 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_8),
.B1(n_13),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_46),
.A2(n_41),
.B1(n_18),
.B2(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_53),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_60),
.Y(n_110)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_82),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_0),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_17),
.Y(n_78)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_39),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_41),
.B1(n_18),
.B2(n_36),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_32),
.B1(n_29),
.B2(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_100),
.A2(n_63),
.B1(n_59),
.B2(n_56),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_33),
.B1(n_16),
.B2(n_21),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_25),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_25),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_29),
.B1(n_42),
.B2(n_15),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_29),
.B1(n_42),
.B2(n_15),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_54),
.A2(n_23),
.B1(n_33),
.B2(n_15),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_20),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_42),
.B1(n_16),
.B2(n_27),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_20),
.B1(n_81),
.B2(n_65),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_138),
.A2(n_131),
.B1(n_127),
.B2(n_137),
.Y(n_209)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_140),
.B(n_161),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_46),
.B1(n_72),
.B2(n_86),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_141),
.A2(n_180),
.B1(n_125),
.B2(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_49),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_121),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_61),
.B1(n_60),
.B2(n_67),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_149),
.Y(n_216)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_69),
.B(n_57),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_152),
.A2(n_166),
.B(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_27),
.B1(n_21),
.B2(n_16),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_75),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_64),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_97),
.B(n_82),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_169),
.B(n_181),
.Y(n_214)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_82),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_173),
.Y(n_217)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_176),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_120),
.A2(n_73),
.B1(n_77),
.B2(n_62),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_40),
.B(n_30),
.C(n_107),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_79),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_118),
.Y(n_177)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_177),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_92),
.A2(n_79),
.B1(n_70),
.B2(n_68),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_94),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_91),
.B1(n_121),
.B2(n_130),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_185),
.A2(n_201),
.B1(n_203),
.B2(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_166),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_91),
.B1(n_55),
.B2(n_51),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_98),
.B1(n_102),
.B2(n_92),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_211),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_152),
.A2(n_130),
.B1(n_125),
.B2(n_102),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_159),
.B(n_164),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_162),
.B1(n_174),
.B2(n_145),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_98),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_37),
.A3(n_108),
.B1(n_103),
.B2(n_124),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_167),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_147),
.A2(n_124),
.B1(n_108),
.B2(n_103),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_222),
.B(n_158),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_144),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_223),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_138),
.B(n_153),
.Y(n_224)
);

OAI31xp33_ASAP7_75t_L g282 ( 
.A1(n_224),
.A2(n_232),
.A3(n_236),
.B(n_237),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_150),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_224),
.C(n_223),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_147),
.B1(n_175),
.B2(n_151),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_245),
.B1(n_230),
.B2(n_246),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_179),
.B1(n_178),
.B2(n_173),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_227),
.A2(n_235),
.B1(n_218),
.B2(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_147),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_229),
.B(n_231),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_167),
.B(n_159),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_164),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_218),
.C(n_200),
.Y(n_265)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_160),
.B1(n_169),
.B2(n_178),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_SL g237 ( 
.A(n_184),
.B(n_140),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_248),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_170),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_241),
.B(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_161),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_214),
.B(n_165),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_252),
.Y(n_262)
);

AO21x2_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_148),
.B(n_142),
.Y(n_250)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_139),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_154),
.Y(n_255)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_259),
.Y(n_288)
);

AO21x2_ASAP7_75t_L g257 ( 
.A1(n_203),
.A2(n_149),
.B(n_1),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_194),
.B1(n_189),
.B2(n_183),
.Y(n_289)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_207),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_10),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_261),
.A2(n_216),
.B(n_188),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_285),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_251),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_269),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_246),
.B1(n_250),
.B2(n_230),
.Y(n_299)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_231),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_281),
.C(n_233),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_218),
.B(n_202),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_274),
.A2(n_190),
.B(n_198),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_225),
.B(n_229),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_202),
.B1(n_201),
.B2(n_185),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_284),
.B1(n_250),
.B2(n_257),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_195),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_200),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_202),
.B1(n_213),
.B2(n_222),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_228),
.B(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_190),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_194),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_282),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_232),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_297),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_306),
.B1(n_307),
.B2(n_311),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_308),
.B1(n_286),
.B2(n_289),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_248),
.B(n_254),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_301),
.A2(n_309),
.B(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_243),
.C(n_238),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_313),
.C(n_320),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_291),
.B(n_293),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_282),
.B(n_279),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_250),
.B1(n_257),
.B2(n_258),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_250),
.B1(n_257),
.B2(n_253),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_270),
.A2(n_257),
.B1(n_212),
.B2(n_252),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_277),
.A2(n_216),
.B1(n_186),
.B2(n_206),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_186),
.Y(n_312)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_205),
.B(n_188),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_316),
.A2(n_322),
.B(n_309),
.Y(n_327)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_285),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_267),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_205),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_286),
.A2(n_188),
.B1(n_206),
.B2(n_40),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_292),
.B1(n_268),
.B2(n_287),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_291),
.A2(n_40),
.B1(n_37),
.B2(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_334),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_327),
.A2(n_343),
.B(n_301),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_329),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_339),
.B1(n_340),
.B2(n_342),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_273),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_344),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_318),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_289),
.B1(n_283),
.B2(n_268),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_288),
.B1(n_262),
.B2(n_271),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_297),
.A2(n_287),
.B(n_271),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_263),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_319),
.A2(n_263),
.B1(n_260),
.B2(n_1),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_295),
.B1(n_317),
.B2(n_323),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_260),
.B1(n_1),
.B2(n_37),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_348),
.A2(n_321),
.B1(n_310),
.B2(n_322),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_298),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_349)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_351),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_298),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_352),
.B(n_356),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_302),
.C(n_320),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_361),
.C(n_367),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_354),
.A2(n_360),
.B(n_363),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_344),
.B(n_314),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_297),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_365),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_324),
.A2(n_315),
.B(n_307),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_294),
.C(n_295),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_312),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_362),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_324),
.A2(n_303),
.B(n_316),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_294),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_330),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_383),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_346),
.Y(n_376)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_369),
.A2(n_332),
.B1(n_339),
.B2(n_345),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_378),
.A2(n_380),
.B1(n_382),
.B2(n_326),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_359),
.A2(n_335),
.B1(n_328),
.B2(n_331),
.Y(n_380)
);

AOI322xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_337),
.A3(n_329),
.B1(n_341),
.B2(n_331),
.C1(n_327),
.C2(n_328),
.Y(n_381)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_381),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_357),
.C(n_358),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_364),
.A2(n_360),
.B1(n_326),
.B2(n_341),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_367),
.B1(n_363),
.B2(n_311),
.Y(n_397)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_389),
.Y(n_398)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_388),
.B(n_370),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_391),
.B(n_392),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_372),
.B(n_370),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_364),
.B1(n_337),
.B2(n_371),
.Y(n_394)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_400),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_372),
.B(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

OAI321xp33_ASAP7_75t_L g410 ( 
.A1(n_401),
.A2(n_403),
.A3(n_373),
.B1(n_384),
.B2(n_374),
.C(n_377),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_354),
.B(n_355),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_393),
.B(n_389),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_348),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_383),
.C(n_385),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_411),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_403),
.B(n_387),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_410),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_385),
.C(n_357),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_379),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_365),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_374),
.C(n_379),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_415),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_373),
.C(n_384),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_416),
.A2(n_421),
.B(n_424),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_387),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_420),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_380),
.C(n_394),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_406),
.A2(n_368),
.B(n_308),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_423),
.B(n_8),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_413),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_1),
.C(n_6),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_425),
.B(n_6),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g426 ( 
.A1(n_424),
.A2(n_407),
.B(n_409),
.C(n_9),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_427),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_428),
.A2(n_429),
.B(n_430),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_417),
.A2(n_11),
.B(n_12),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_11),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_R g435 ( 
.A(n_431),
.B(n_421),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_432),
.B(n_425),
.C(n_13),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_12),
.C(n_13),
.Y(n_437)
);

NAND4xp25_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_434),
.C(n_433),
.D(n_14),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_R g441 ( 
.A1(n_440),
.A2(n_12),
.B1(n_438),
.B2(n_393),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_441),
.Y(n_442)
);


endmodule