module fake_jpeg_780_n_455 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_74),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_36),
.B1(n_25),
.B2(n_34),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_23),
.B(n_0),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_23),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_17),
.Y(n_120)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_1),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_28),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_28),
.Y(n_85)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_95),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_90),
.B(n_99),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_22),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_17),
.B1(n_41),
.B2(n_36),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_122),
.B1(n_127),
.B2(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_27),
.B1(n_39),
.B2(n_42),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_49),
.A2(n_81),
.B1(n_85),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_143),
.B1(n_59),
.B2(n_86),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_120),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_41),
.B1(n_25),
.B2(n_36),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_51),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_59),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_37),
.B1(n_25),
.B2(n_40),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_46),
.B(n_21),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_21),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_91),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_42),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_4),
.B(n_5),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_63),
.B(n_40),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_52),
.B(n_40),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_45),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_50),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_27),
.B1(n_66),
.B2(n_28),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_56),
.A2(n_38),
.B1(n_35),
.B2(n_39),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_38),
.B1(n_44),
.B2(n_42),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_82),
.A2(n_44),
.B1(n_38),
.B2(n_39),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_147),
.A2(n_161),
.B1(n_184),
.B2(n_185),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_88),
.A2(n_133),
.B(n_109),
.C(n_89),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_149),
.B(n_151),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_78),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_173),
.C(n_178),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_107),
.A2(n_44),
.B1(n_22),
.B2(n_27),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_154),
.B(n_155),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_157),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_197),
.B1(n_4),
.B2(n_6),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_170),
.Y(n_200)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_77),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_167),
.B(n_180),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_172),
.Y(n_203)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_67),
.B1(n_84),
.B2(n_26),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_91),
.B(n_26),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_98),
.B(n_79),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_79),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_187),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_128),
.A2(n_26),
.B1(n_61),
.B2(n_47),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_26),
.C(n_75),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_182),
.Y(n_242)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_98),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_98),
.A2(n_73),
.B1(n_26),
.B2(n_18),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_26),
.B1(n_18),
.B2(n_5),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_3),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_4),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_190),
.Y(n_220)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_4),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_125),
.B(n_93),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_114),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_114),
.A2(n_26),
.B(n_5),
.C(n_6),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_18),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_112),
.B1(n_105),
.B2(n_113),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_199),
.A2(n_232),
.B1(n_200),
.B2(n_211),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_96),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_213),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_136),
.B1(n_106),
.B2(n_101),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_211),
.B1(n_215),
.B2(n_218),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_209),
.A2(n_13),
.B(n_165),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_136),
.B1(n_96),
.B2(n_123),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_216),
.B1(n_221),
.B2(n_229),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_106),
.B1(n_101),
.B2(n_93),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_121),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_161),
.A2(n_100),
.B1(n_125),
.B2(n_108),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_100),
.B1(n_108),
.B2(n_119),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_108),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_166),
.A2(n_119),
.B1(n_111),
.B2(n_18),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_226),
.B1(n_245),
.B2(n_174),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_146),
.A2(n_111),
.B1(n_8),
.B2(n_9),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_111),
.B1(n_8),
.B2(n_10),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_164),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_144),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_158),
.B(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_12),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_159),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_183),
.C(n_175),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_249),
.C(n_256),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_183),
.C(n_175),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_149),
.B(n_196),
.C(n_178),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_250),
.B(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_207),
.B(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_259),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_231),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_184),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_256),
.B(n_239),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_186),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_184),
.B(n_171),
.C(n_181),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_258),
.B(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_169),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_205),
.A2(n_170),
.B(n_177),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_195),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_179),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_283),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_163),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_267),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_272),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_235),
.A2(n_185),
.B(n_192),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_182),
.C(n_148),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_190),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_278),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_198),
.B(n_188),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_277),
.B(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_204),
.A2(n_233),
.B(n_200),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_200),
.B(n_232),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_204),
.A2(n_232),
.B(n_234),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_233),
.B(n_234),
.C(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_288),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_241),
.B(n_231),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_242),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_283),
.A2(n_201),
.B1(n_218),
.B2(n_239),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_292),
.A2(n_269),
.B(n_260),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_208),
.B1(n_239),
.B2(n_210),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_321),
.B1(n_254),
.B2(n_264),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_325),
.C(n_249),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_299),
.B(n_307),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_267),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_302),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_267),
.Y(n_302)
);

OAI32xp33_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_216),
.A3(n_245),
.B1(n_221),
.B2(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_312),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_243),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_253),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_315),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_263),
.A2(n_206),
.B1(n_243),
.B2(n_222),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_247),
.B1(n_254),
.B2(n_287),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_252),
.A2(n_206),
.A3(n_223),
.B1(n_230),
.B2(n_227),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_246),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_275),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_250),
.A2(n_227),
.B1(n_223),
.B2(n_246),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_261),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_281),
.B(n_248),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_327),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_332),
.Y(n_372)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_283),
.B(n_276),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_329),
.A2(n_330),
.B(n_339),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_304),
.B1(n_295),
.B2(n_324),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_299),
.C(n_307),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_261),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_349),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_272),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_337),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_319),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_311),
.A2(n_291),
.B(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_291),
.A2(n_285),
.B(n_284),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_348),
.B(n_351),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_271),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_350),
.Y(n_357)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_346),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_301),
.B1(n_326),
.B2(n_305),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_318),
.A2(n_255),
.B(n_262),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_288),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_313),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_316),
.A2(n_279),
.B(n_268),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_313),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_354),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_270),
.B(n_273),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_353),
.A2(n_293),
.B(n_323),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_309),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_309),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_326),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_367),
.B1(n_368),
.B2(n_373),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_380),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_290),
.B1(n_304),
.B2(n_324),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_366),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_334),
.A2(n_304),
.B1(n_321),
.B2(n_292),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_294),
.B1(n_322),
.B2(n_308),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_322),
.B1(n_323),
.B2(n_247),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_332),
.B(n_296),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_374),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_333),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_375),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_312),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_368),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_347),
.A2(n_306),
.B1(n_320),
.B2(n_273),
.Y(n_378)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_329),
.A2(n_320),
.B(n_286),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_354),
.B1(n_355),
.B2(n_352),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_382),
.A2(n_378),
.B1(n_381),
.B2(n_348),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_383),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_338),
.C(n_343),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_385),
.C(n_392),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_338),
.C(n_343),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_375),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_391),
.Y(n_406)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_349),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_365),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_375),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_336),
.C(n_339),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_356),
.C(n_335),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_401),
.C(n_402),
.Y(n_409)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_377),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_358),
.B(n_337),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_361),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_356),
.C(n_350),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_341),
.C(n_345),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_407),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_405),
.B(n_414),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_371),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_392),
.A2(n_397),
.B(n_393),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_416),
.B1(n_418),
.B2(n_387),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_415),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_371),
.C(n_360),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_360),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_380),
.C(n_353),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_398),
.C(n_402),
.Y(n_426)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_396),
.B1(n_400),
.B2(n_376),
.Y(n_428)
);

OAI321xp33_ASAP7_75t_L g420 ( 
.A1(n_406),
.A2(n_357),
.A3(n_400),
.B1(n_386),
.B2(n_387),
.C(n_383),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_376),
.B1(n_379),
.B2(n_364),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_413),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_421),
.B(n_424),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_384),
.C(n_385),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_428),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_423),
.B(n_411),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g424 ( 
.A(n_415),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_431),
.Y(n_439)
);

OAI322xp33_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_407),
.A3(n_412),
.B1(n_414),
.B2(n_417),
.C1(n_404),
.C2(n_393),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_430),
.A2(n_330),
.B(n_351),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_366),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_434),
.B1(n_436),
.B2(n_438),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_433),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_426),
.A2(n_340),
.B1(n_346),
.B2(n_342),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_438),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_403),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_278),
.B(n_303),
.Y(n_443)
);

OAI221xp5_ASAP7_75t_L g441 ( 
.A1(n_435),
.A2(n_425),
.B1(n_429),
.B2(n_280),
.C(n_274),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_441),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_444),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_439),
.A2(n_303),
.B(n_289),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_432),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_445),
.B(n_442),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_450),
.Y(n_452)
);

BUFx24_ASAP7_75t_SL g453 ( 
.A(n_452),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_451),
.B(n_447),
.C(n_437),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_442),
.Y(n_455)
);


endmodule