module fake_jpeg_20802_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_16),
.B1(n_6),
.B2(n_11),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_6),
.A2(n_4),
.B1(n_11),
.B2(n_9),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_13),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_25),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_21),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_24),
.C(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_20),
.B1(n_28),
.B2(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_9),
.Y(n_32)
);


endmodule