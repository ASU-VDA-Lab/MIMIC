module fake_jpeg_3940_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_23),
.B(n_6),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_31),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_53),
.B(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_55),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_59),
.Y(n_118)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_62),
.Y(n_122)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_17),
.B1(n_30),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_17),
.B1(n_30),
.B2(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_73),
.Y(n_102)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_17),
.B1(n_32),
.B2(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_29),
.CI(n_33),
.CON(n_84),
.SN(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_89),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_26),
.C(n_32),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_19),
.Y(n_116)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_18),
.B1(n_22),
.B2(n_28),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_27),
.B1(n_24),
.B2(n_31),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_36),
.B(n_33),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_31),
.B1(n_25),
.B2(n_19),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_125),
.B1(n_8),
.B2(n_10),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_25),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_29),
.B1(n_31),
.B2(n_25),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_68),
.A3(n_80),
.B1(n_77),
.B2(n_57),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_77),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_25),
.B1(n_15),
.B2(n_2),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_84),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_128),
.CON(n_173),
.SN(n_173)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_130),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_71),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_144),
.B1(n_153),
.B2(n_106),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_136),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_125),
.B1(n_110),
.B2(n_116),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_60),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_83),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_90),
.B(n_70),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_116),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_56),
.A3(n_50),
.B1(n_82),
.B2(n_65),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_51),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_50),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_82),
.B1(n_72),
.B2(n_64),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_15),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_155),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_15),
.B1(n_60),
.B2(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_51),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_102),
.B(n_6),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_180),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_111),
.B1(n_106),
.B2(n_102),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_167),
.B1(n_175),
.B2(n_143),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_176),
.B1(n_132),
.B2(n_136),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_112),
.B1(n_119),
.B2(n_100),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_144),
.C(n_150),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_156),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_112),
.B1(n_119),
.B2(n_124),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_117),
.B1(n_124),
.B2(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_121),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_130),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_192),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_131),
.B1(n_139),
.B2(n_145),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_162),
.C(n_163),
.Y(n_212)
);

AOI321xp33_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_204),
.A3(n_205),
.B1(n_206),
.B2(n_207),
.C(n_186),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_152),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_128),
.B1(n_140),
.B2(n_147),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_173),
.B1(n_168),
.B2(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_128),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_139),
.B(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_0),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_172),
.C(n_161),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_210),
.B(n_213),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_216),
.C(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_165),
.C(n_184),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_165),
.C(n_171),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_171),
.C(n_174),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_221),
.C(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_174),
.C(n_170),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_178),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_177),
.C(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_230),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_194),
.B1(n_203),
.B2(n_190),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_235),
.B1(n_207),
.B2(n_188),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_201),
.B(n_197),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_219),
.B(n_189),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_233),
.B1(n_206),
.B2(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_203),
.B1(n_191),
.B2(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_191),
.B1(n_208),
.B2(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_216),
.C(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_207),
.C(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_209),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_234),
.C(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_166),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_244),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_240),
.B1(n_227),
.B2(n_248),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_158),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_247),
.C(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_187),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_228),
.B(n_233),
.Y(n_252)
);

NAND4xp25_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_192),
.C(n_207),
.D(n_202),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_198),
.B1(n_238),
.B2(n_200),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_247),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_255),
.A3(n_245),
.B1(n_254),
.B2(n_232),
.C1(n_251),
.C2(n_159),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_246),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_230),
.C(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_246),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_259),
.B(n_261),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_262),
.C(n_5),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_232),
.A3(n_158),
.B1(n_176),
.B2(n_10),
.C1(n_4),
.C2(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_265),
.B(n_6),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_12),
.C(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_266),
.B(n_4),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_268),
.A3(n_269),
.B1(n_14),
.B2(n_1),
.C1(n_2),
.C2(n_3),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_263),
.C2(n_257),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_0),
.Y(n_273)
);


endmodule