module real_jpeg_5728_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_145),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_1),
.A2(n_30),
.B1(n_218),
.B2(n_277),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_66),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_2),
.A2(n_66),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_3),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_6),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_6),
.Y(n_224)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_6),
.B(n_10),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_7),
.A2(n_98),
.B1(n_99),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_7),
.A2(n_98),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_7),
.A2(n_98),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_56),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_10),
.A2(n_56),
.B1(n_192),
.B2(n_196),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_56),
.B1(n_172),
.B2(n_241),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_10),
.A2(n_268),
.B(n_269),
.C(n_273),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_10),
.B(n_109),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_10),
.B(n_303),
.C(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_10),
.B(n_96),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_10),
.B(n_91),
.C(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_10),
.B(n_32),
.Y(n_340)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_12),
.Y(n_389)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_387),
.B(n_390),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_199),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_198),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_19),
.B(n_148),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_139),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_137),
.B2(n_138),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_58),
.B2(n_59),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_23),
.A2(n_24),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_23),
.A2(n_24),
.B1(n_160),
.B2(n_341),
.Y(n_366)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_24),
.B(n_206),
.C(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_24),
.B(n_160),
.C(n_266),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_54),
.B2(n_57),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_25),
.A2(n_31),
.B1(n_54),
.B2(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_29),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_31),
.A2(n_54),
.B(n_57),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_44),
.Y(n_31)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_34),
.Y(n_145)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_35),
.Y(n_268)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_56),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_106),
.B2(n_136),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_69),
.B1(n_96),
.B2(n_97),
.Y(n_61)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_68),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_69),
.B(n_143),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_69),
.A2(n_96),
.B1(n_143),
.B2(n_162),
.Y(n_226)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_70),
.A2(n_71),
.B1(n_161),
.B2(n_167),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_70),
.B(n_71),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_88),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_81),
.B2(n_84),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_75),
.Y(n_301)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g323 ( 
.A(n_90),
.Y(n_323)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_137),
.C(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_136),
.B1(n_140),
.B2(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_133),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_121),
.Y(n_107)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_108),
.A2(n_121),
.B1(n_191),
.B2(n_210),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_108),
.A2(n_121),
.B1(n_191),
.B2(n_210),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_108),
.A2(n_121),
.B(n_191),
.Y(n_352)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_115),
.B2(n_119),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_191),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_137),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_138),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_232),
.C(n_242),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_137),
.A2(n_138),
.B1(n_242),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_137),
.A2(n_138),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_138),
.B(n_226),
.C(n_352),
.Y(n_370)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_143),
.B(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_168),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_149),
.Y(n_384)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_154),
.A2(n_155),
.B(n_160),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_159),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_160),
.A2(n_337),
.B1(n_338),
.B2(n_341),
.Y(n_336)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_168),
.B(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B(n_197),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_189),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_170),
.A2(n_189),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_170),
.A2(n_197),
.B1(n_230),
.B2(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_178),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_179),
.B(n_240),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_181),
.A2(n_240),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_181),
.A2(n_240),
.B1(n_276),
.B2(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_186),
.Y(n_292)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx5_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_381),
.B(n_386),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI211xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_280),
.B(n_376),
.C(n_380),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_255),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_203),
.A2(n_255),
.B(n_377),
.C(n_379),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_244),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_204),
.B(n_244),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_228),
.C(n_231),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_228),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_225),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_207),
.A2(n_215),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_207),
.A2(n_264),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_208),
.A2(n_209),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_236),
.B(n_239),
.Y(n_235)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_226),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_226),
.B(n_233),
.C(n_320),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_226),
.A2(n_227),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_233),
.A2(n_234),
.B1(n_299),
.B2(n_307),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_233),
.B(n_307),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_235),
.Y(n_368)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_253),
.B2(n_254),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_250),
.B(n_252),
.C(n_254),
.Y(n_385)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_256),
.B(n_258),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_265),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_259),
.B(n_262),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_275),
.C(n_313),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_264),
.B(n_333),
.C(n_335),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_265),
.B(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_266),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_267),
.A2(n_274),
.B1(n_275),
.B2(n_358),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_275),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_294),
.Y(n_295)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_360),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_345),
.B(n_359),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_330),
.B(n_344),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_317),
.B(n_329),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_309),
.B(n_316),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_296),
.B(n_308),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_293),
.B(n_295),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_291),
.A2(n_297),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_339),
.C(n_341),
.Y(n_355)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_326),
.B2(n_327),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_327),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_343),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_343),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_335),
.B1(n_336),
.B2(n_342),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_347),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_355),
.C(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_363),
.B(n_371),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_363),
.C(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.C(n_369),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_367),
.A2(n_369),
.B1(n_370),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_373),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_385),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_388),
.Y(n_391)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);


endmodule