module fake_jpeg_1632_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_9),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_49),
.B(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_9),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_62),
.Y(n_115)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_56),
.Y(n_133)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_8),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_10),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_10),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_85),
.Y(n_146)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_69),
.Y(n_144)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_79),
.B(n_92),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_5),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_87),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_11),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_0),
.Y(n_145)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_42),
.B1(n_20),
.B2(n_26),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_26),
.B1(n_42),
.B2(n_20),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_35),
.B1(n_43),
.B2(n_27),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_109),
.B1(n_136),
.B2(n_80),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_23),
.B1(n_29),
.B2(n_41),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_54),
.A2(n_23),
.B1(n_29),
.B2(n_41),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_120),
.A2(n_128),
.B1(n_113),
.B2(n_99),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_121)
);

AOI22x1_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_142),
.B1(n_90),
.B2(n_85),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_49),
.B(n_38),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_138),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_27),
.B1(n_24),
.B2(n_46),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_50),
.A2(n_24),
.B1(n_46),
.B2(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_51),
.B(n_12),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_16),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_68),
.A2(n_46),
.B1(n_11),
.B2(n_15),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_63),
.A2(n_16),
.B1(n_1),
.B2(n_3),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_108),
.B1(n_137),
.B2(n_100),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_113),
.Y(n_174)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_151),
.A2(n_179),
.B1(n_187),
.B2(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_65),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_159),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_140),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_167),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_172),
.B1(n_132),
.B2(n_114),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_16),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_162),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_56),
.B(n_55),
.C(n_67),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_184),
.B(n_134),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_55),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_67),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_72),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_72),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_118),
.Y(n_171)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_80),
.B1(n_56),
.B2(n_86),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_119),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_177),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_126),
.C(n_111),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_180),
.C(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_104),
.B(n_98),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_181),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_143),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_124),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_132),
.B(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_121),
.B(n_133),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_130),
.Y(n_184)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_121),
.A2(n_129),
.B1(n_128),
.B2(n_97),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_188),
.B1(n_129),
.B2(n_100),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_133),
.C(n_120),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_105),
.A3(n_125),
.B1(n_134),
.B2(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_147),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_198),
.B1(n_206),
.B2(n_207),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_179),
.A2(n_125),
.B1(n_105),
.B2(n_114),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_213),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_193),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_168),
.B1(n_154),
.B2(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_219),
.B1(n_171),
.B2(n_165),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_151),
.B1(n_185),
.B2(n_173),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_186),
.B1(n_185),
.B2(n_187),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_217),
.B1(n_150),
.B2(n_157),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_163),
.B(n_174),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_203),
.B(n_215),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_174),
.B1(n_162),
.B2(n_172),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_175),
.A2(n_149),
.B1(n_188),
.B2(n_178),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_205),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_228),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_167),
.B(n_171),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_240),
.B(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_158),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_226),
.A2(n_212),
.B1(n_200),
.B2(n_195),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_233),
.B1(n_236),
.B2(n_196),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_148),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_216),
.C(n_206),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_199),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_238),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_242),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_189),
.B1(n_203),
.B2(n_204),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_221),
.B1(n_228),
.B2(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_243),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_250),
.B1(n_257),
.B2(n_236),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_240),
.B(n_237),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_237),
.C(n_240),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_219),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_256),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_212),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_274),
.B1(n_258),
.B2(n_253),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_238),
.A3(n_237),
.B1(n_231),
.B2(n_232),
.C1(n_226),
.C2(n_221),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_259),
.A3(n_256),
.B1(n_257),
.B2(n_260),
.C1(n_252),
.C2(n_190),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_231),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_272),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_273),
.B(n_245),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_211),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_271),
.C(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_251),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_235),
.C(n_190),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_222),
.B(n_233),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_233),
.B1(n_227),
.B2(n_239),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_250),
.B1(n_255),
.B2(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_264),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_244),
.B1(n_255),
.B2(n_251),
.Y(n_277)
);

AOI31xp67_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_282),
.A3(n_252),
.B(n_225),
.Y(n_293)
);

OA21x2_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_283),
.B(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_285),
.A2(n_233),
.B1(n_249),
.B2(n_243),
.Y(n_294)
);

FAx1_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_265),
.CI(n_273),
.CON(n_287),
.SN(n_287)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_293),
.B(n_197),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_263),
.C(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_292),
.B1(n_294),
.B2(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_271),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_270),
.B(n_269),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_247),
.B(n_242),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_257),
.B1(n_268),
.B2(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_299),
.B1(n_290),
.B2(n_197),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_279),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_298),
.B(n_287),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_275),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_301),
.C(n_286),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_198),
.B1(n_208),
.B2(n_209),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_301),
.B(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_306),
.C(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_306),
.B(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_191),
.B(n_312),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_209),
.C(n_218),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_191),
.C(n_210),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);


endmodule