module fake_ibex_303_n_1084 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_132, n_174, n_210, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1084);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_132;
input n_174;
input n_210;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1084;

wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1079;
wire n_1031;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_1018;
wire n_258;
wire n_861;
wire n_930;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_1070;
wire n_454;
wire n_980;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_506;
wire n_562;
wire n_444;
wire n_564;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_1073;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_912;
wire n_1058;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_231;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_87),
.B(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_104),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_29),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_156),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_55),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_151),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_114),
.B(n_93),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_122),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_18),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_74),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_148),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_52),
.B(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_83),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_47),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_45),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_177),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_61),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_103),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_77),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_90),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_63),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_70),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_60),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_175),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_27),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_138),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_127),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_180),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_14),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_95),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_120),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_178),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_82),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_20),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_123),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_102),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_24),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_97),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_66),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_186),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_118),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_135),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_196),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_36),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_206),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_9),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_88),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_98),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_80),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_183),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_179),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_165),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_112),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_157),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_28),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_59),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_105),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_48),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_57),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_75),
.B(n_86),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_47),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_10),
.B(n_143),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_73),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_68),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_24),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_115),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_109),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_113),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_202),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_15),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_65),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_130),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_194),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_94),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_23),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_31),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_108),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_81),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_192),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_188),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_42),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_205),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_257),
.B(n_0),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_328),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_217),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_278),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_4),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_227),
.Y(n_360)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_217),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_5),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_220),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_282),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_239),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_369)
);

INVx6_ASAP7_75t_L g370 ( 
.A(n_307),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_216),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_286),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_R g376 ( 
.A1(n_287),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_12),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_224),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_232),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_13),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_227),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_234),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_236),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_246),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_288),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_251),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_253),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_227),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_254),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_260),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_267),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_293),
.B(n_16),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_226),
.B(n_16),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_268),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_226),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_227),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_239),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_273),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_273),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_274),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_250),
.B(n_19),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_293),
.B(n_326),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_281),
.B(n_21),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_275),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_281),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

XNOR2x2_ASAP7_75t_L g412 ( 
.A(n_294),
.B(n_21),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_262),
.B(n_22),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_228),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_215),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_252),
.B(n_50),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_277),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_235),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_265),
.B(n_22),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_279),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_256),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_346),
.B(n_26),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_346),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_290),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_284),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_237),
.B(n_30),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_291),
.A2(n_297),
.B(n_295),
.Y(n_431)
);

AND3x2_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_365),
.C(n_356),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_351),
.C(n_247),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_357),
.B(n_229),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g441 ( 
.A(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

AND3x2_ASAP7_75t_L g443 ( 
.A(n_365),
.B(n_331),
.C(n_248),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_406),
.B(n_357),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_378),
.B(n_238),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_431),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_357),
.B(n_351),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_230),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_375),
.B(n_299),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_230),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_361),
.B(n_301),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_231),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_361),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_390),
.B(n_416),
.Y(n_461)
);

AO21x2_ASAP7_75t_L g462 ( 
.A1(n_420),
.A2(n_305),
.B(n_303),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_358),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_231),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_374),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_361),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_354),
.B(n_340),
.C(n_241),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_370),
.B(n_416),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_370),
.B(n_309),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_370),
.B(n_353),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_372),
.B(n_373),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_430),
.A2(n_270),
.B1(n_308),
.B2(n_310),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_368),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_233),
.Y(n_484)
);

AND3x4_ASAP7_75t_L g485 ( 
.A(n_376),
.B(n_332),
.C(n_218),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_372),
.B(n_240),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_292),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_379),
.B(n_292),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_379),
.B(n_343),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_377),
.B(n_259),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_364),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_364),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_423),
.B(n_343),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_380),
.B(n_349),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_380),
.B(n_349),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_386),
.B(n_352),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_383),
.B(n_313),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_383),
.B(n_352),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_384),
.B(n_221),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_384),
.B(n_315),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_L g507 ( 
.A(n_369),
.B(n_283),
.C(n_276),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_430),
.A2(n_289),
.B1(n_345),
.B2(n_320),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_364),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_385),
.B(n_223),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_374),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_386),
.B(n_285),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_417),
.A2(n_300),
.B1(n_335),
.B2(n_347),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_355),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_414),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_L g522 ( 
.A(n_385),
.B(n_284),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_389),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_389),
.B(n_225),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_355),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_381),
.B(n_317),
.C(n_316),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_386),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_391),
.A2(n_319),
.B1(n_334),
.B2(n_339),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_391),
.B(n_244),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_393),
.B(n_284),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_400),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_414),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_393),
.A2(n_228),
.B1(n_243),
.B2(n_338),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_363),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_394),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_363),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_394),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_395),
.B(n_245),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_395),
.B(n_249),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_523),
.B(n_398),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_537),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_478),
.B(n_387),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_398),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_442),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_445),
.B(n_426),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_404),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_441),
.A2(n_426),
.B1(n_405),
.B2(n_413),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_461),
.B(n_426),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_452),
.B(n_408),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_408),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_481),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_418),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_490),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_490),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_454),
.B(n_418),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_497),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_537),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_527),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_438),
.B(n_243),
.Y(n_565)
);

A2O1A1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_463),
.A2(n_421),
.B(n_428),
.C(n_427),
.Y(n_566)
);

NOR4xp25_ASAP7_75t_SL g567 ( 
.A(n_534),
.B(n_376),
.C(n_329),
.D(n_304),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_457),
.B(n_421),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_467),
.A2(n_403),
.B(n_427),
.C(n_425),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_451),
.A2(n_403),
.B(n_425),
.C(n_367),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_520),
.B(n_401),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_527),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_470),
.B(n_517),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_464),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_439),
.B(n_359),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_462),
.B(n_367),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_462),
.B(n_388),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_451),
.A2(n_402),
.B(n_388),
.C(n_409),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_492),
.B(n_359),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_485),
.A2(n_422),
.B1(n_256),
.B2(n_272),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_450),
.B(n_464),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_447),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_462),
.B(n_399),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_447),
.B(n_362),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_495),
.A2(n_424),
.B(n_411),
.C(n_409),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_333),
.C(n_269),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_459),
.A2(n_321),
.B1(n_314),
.B2(n_255),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_473),
.B(n_272),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_447),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_470),
.B(n_263),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_484),
.A2(n_321),
.B1(n_338),
.B2(n_255),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_470),
.B(n_264),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_528),
.A2(n_415),
.B1(n_411),
.B2(n_402),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_517),
.B(n_480),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

O2A1O1Ixp5_ASAP7_75t_L g600 ( 
.A1(n_442),
.A2(n_415),
.B(n_399),
.C(n_371),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_456),
.B(n_371),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_479),
.B(n_266),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_508),
.B(n_494),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_449),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_495),
.A2(n_261),
.B(n_314),
.C(n_302),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_455),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_311),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_494),
.B(n_271),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_455),
.B(n_330),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_491),
.A2(n_261),
.B1(n_330),
.B2(n_342),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_491),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_493),
.B(n_296),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_513),
.B(n_306),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_516),
.B(n_242),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_489),
.B(n_322),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_468),
.B(n_323),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_468),
.B(n_336),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_514),
.B(n_337),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_514),
.B(n_312),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_465),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_535),
.B(n_412),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_515),
.A2(n_341),
.B1(n_284),
.B2(n_412),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_432),
.B(n_504),
.Y(n_627)
);

AO22x1_ASAP7_75t_L g628 ( 
.A1(n_513),
.A2(n_341),
.B1(n_31),
.B2(n_32),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_512),
.B(n_341),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_534),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_515),
.B(n_341),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_487),
.B(n_51),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_501),
.B(n_477),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_477),
.A2(n_488),
.B1(n_501),
.B2(n_509),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_536),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_524),
.B(n_429),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_443),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_496),
.B(n_429),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_496),
.B(n_429),
.Y(n_639)
);

OAI221xp5_ASAP7_75t_L g640 ( 
.A1(n_529),
.A2(n_507),
.B1(n_506),
.B2(n_503),
.C(n_526),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_496),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_53),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_498),
.B(n_35),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_610),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_606),
.Y(n_646)
);

O2A1O1Ixp5_ASAP7_75t_L g647 ( 
.A1(n_598),
.A2(n_476),
.B(n_458),
.C(n_474),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_633),
.A2(n_449),
.B(n_544),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_546),
.A2(n_466),
.B(n_500),
.Y(n_649)
);

O2A1O1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_589),
.A2(n_466),
.B(n_510),
.C(n_545),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_562),
.A2(n_510),
.B(n_505),
.C(n_531),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_510),
.B(n_460),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_642),
.A2(n_542),
.B(n_433),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_556),
.B(n_460),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_549),
.A2(n_552),
.B(n_577),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_558),
.B(n_469),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_612),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_614),
.B(n_469),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_610),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_610),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_555),
.B(n_542),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_557),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_37),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_568),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_603),
.A2(n_625),
.B(n_640),
.C(n_560),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_563),
.B(n_530),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_550),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_595),
.B(n_485),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_583),
.A2(n_522),
.B1(n_532),
.B2(n_533),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_37),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_SL g671 ( 
.A1(n_642),
.A2(n_453),
.B(n_533),
.C(n_471),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_575),
.A2(n_522),
.B(n_434),
.C(n_433),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_601),
.A2(n_434),
.B(n_435),
.C(n_521),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_624),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_563),
.B(n_530),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_565),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_577),
.A2(n_435),
.B(n_446),
.C(n_521),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_578),
.A2(n_440),
.B(n_448),
.C(n_511),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_621),
.B(n_532),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_578),
.A2(n_440),
.B(n_444),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_607),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_581),
.B(n_444),
.C(n_446),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_585),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_SL g684 ( 
.A1(n_554),
.A2(n_483),
.B(n_453),
.C(n_471),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_592),
.B(n_630),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_548),
.A2(n_532),
.B1(n_486),
.B2(n_483),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_600),
.A2(n_499),
.B(n_486),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_551),
.B(n_38),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_587),
.A2(n_499),
.B(n_448),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_593),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_602),
.B(n_532),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_584),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_572),
.A2(n_511),
.B(n_482),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_587),
.A2(n_530),
.B(n_541),
.C(n_482),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_588),
.A2(n_530),
.B(n_541),
.C(n_482),
.Y(n_695)
);

OR2x6_ASAP7_75t_SL g696 ( 
.A(n_591),
.B(n_38),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_572),
.A2(n_482),
.B(n_475),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_631),
.A2(n_532),
.B(n_541),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_548),
.A2(n_541),
.B1(n_475),
.B2(n_41),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_611),
.A2(n_541),
.B1(n_40),
.B2(n_41),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_609),
.B(n_39),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_553),
.B(n_40),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_616),
.A2(n_475),
.B1(n_43),
.B2(n_44),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_570),
.A2(n_137),
.B(n_214),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_634),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_627),
.B(n_46),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_616),
.B(n_46),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_580),
.B(n_48),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_608),
.B(n_49),
.Y(n_709)
);

NOR2x1_ASAP7_75t_L g710 ( 
.A(n_590),
.B(n_49),
.Y(n_710)
);

AO22x1_ASAP7_75t_L g711 ( 
.A1(n_567),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_597),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_638),
.A2(n_639),
.B(n_550),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_626),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_615),
.B(n_79),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_607),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_628),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_613),
.B(n_84),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_643),
.B(n_85),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_SL g721 ( 
.A1(n_579),
.A2(n_89),
.B(n_91),
.C(n_92),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_605),
.B(n_99),
.Y(n_722)
);

BUFx12f_ASAP7_75t_L g723 ( 
.A(n_637),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_550),
.B(n_106),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_620),
.B(n_107),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_571),
.B(n_213),
.Y(n_726)
);

BUFx8_ASAP7_75t_L g727 ( 
.A(n_564),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_623),
.A2(n_116),
.B(n_117),
.C(n_121),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_571),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_604),
.B(n_128),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_547),
.B(n_129),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_635),
.A2(n_132),
.B1(n_134),
.B2(n_140),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_639),
.A2(n_141),
.B(n_142),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_566),
.A2(n_145),
.B(n_150),
.C(n_152),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_636),
.A2(n_203),
.B(n_155),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_617),
.B(n_201),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_604),
.B(n_153),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_569),
.A2(n_158),
.B(n_159),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_641),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_604),
.B(n_163),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_571),
.B(n_164),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_632),
.A2(n_167),
.B(n_168),
.C(n_169),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_667),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_727),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_655),
.A2(n_629),
.B(n_586),
.Y(n_747)
);

AOI21x1_ASAP7_75t_L g748 ( 
.A1(n_653),
.A2(n_573),
.B(n_596),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_660),
.B(n_594),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_700),
.A2(n_619),
.B(n_618),
.C(n_181),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_644),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_685),
.B(n_172),
.Y(n_752)
);

OA21x2_ASAP7_75t_L g753 ( 
.A1(n_677),
.A2(n_173),
.B(n_182),
.Y(n_753)
);

INVx3_ASAP7_75t_SL g754 ( 
.A(n_674),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_645),
.B(n_193),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_649),
.A2(n_650),
.B(n_688),
.C(n_652),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_662),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_668),
.B(n_195),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_659),
.B(n_663),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_714),
.A2(n_671),
.B(n_697),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_727),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_661),
.A2(n_699),
.B1(n_708),
.B2(n_663),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_692),
.B(n_683),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_696),
.B(n_726),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_690),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_693),
.A2(n_689),
.B(n_680),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_689),
.A2(n_678),
.B(n_691),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_694),
.A2(n_673),
.A3(n_739),
.B(n_734),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_723),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_704),
.A2(n_739),
.B(n_735),
.Y(n_770)
);

CKINVDCx11_ASAP7_75t_R g771 ( 
.A(n_718),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_670),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_654),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_702),
.A2(n_676),
.B1(n_682),
.B2(n_706),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_681),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_728),
.A2(n_735),
.A3(n_744),
.B(n_740),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_743),
.B(n_722),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_707),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_713),
.B(n_656),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_701),
.B(n_709),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_733),
.A2(n_712),
.A3(n_732),
.B(n_672),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_724),
.A2(n_742),
.B(n_730),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_646),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_651),
.B(n_741),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_667),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_720),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_647),
.A2(n_705),
.B(n_725),
.C(n_710),
.Y(n_787)
);

AO31x2_ASAP7_75t_L g788 ( 
.A1(n_733),
.A2(n_695),
.A3(n_716),
.B(n_679),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_711),
.B(n_729),
.C(n_658),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_720),
.B(n_657),
.Y(n_790)
);

INVx6_ASAP7_75t_L g791 ( 
.A(n_667),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_686),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_717),
.B(n_738),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_738),
.B(n_703),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_684),
.A2(n_666),
.B(n_675),
.Y(n_795)
);

OAI22x1_ASAP7_75t_L g796 ( 
.A1(n_715),
.A2(n_669),
.B1(n_736),
.B2(n_737),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_721),
.A2(n_655),
.B(n_604),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_698),
.A2(n_664),
.B1(n_518),
.B2(n_441),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_722),
.B(n_426),
.C(n_554),
.Y(n_799)
);

OAI21xp33_ASAP7_75t_L g800 ( 
.A1(n_664),
.A2(n_438),
.B(n_583),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_664),
.B(n_665),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_664),
.A2(n_665),
.B(n_700),
.C(n_562),
.Y(n_802)
);

NAND2x1p5_ASAP7_75t_L g803 ( 
.A(n_674),
.B(n_599),
.Y(n_803)
);

CKINVDCx11_ASAP7_75t_R g804 ( 
.A(n_723),
.Y(n_804)
);

OA21x2_ASAP7_75t_L g805 ( 
.A1(n_677),
.A2(n_678),
.B(n_704),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_664),
.A2(n_665),
.B(n_700),
.C(n_562),
.Y(n_806)
);

AO31x2_ASAP7_75t_L g807 ( 
.A1(n_655),
.A2(n_677),
.A3(n_678),
.B(n_694),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_665),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_SL g809 ( 
.A1(n_744),
.A2(n_655),
.B(n_719),
.C(n_684),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_664),
.A2(n_534),
.B(n_630),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_655),
.A2(n_648),
.B(n_664),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_655),
.A2(n_648),
.B(n_664),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_692),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_664),
.A2(n_665),
.B(n_700),
.C(n_562),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_655),
.A2(n_677),
.A3(n_678),
.B(n_694),
.Y(n_815)
);

AO31x2_ASAP7_75t_L g816 ( 
.A1(n_655),
.A2(n_677),
.A3(n_678),
.B(n_694),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_727),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_655),
.A2(n_677),
.A3(n_678),
.B(n_694),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_653),
.A2(n_687),
.B(n_680),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_655),
.A2(n_604),
.B(n_550),
.Y(n_820)
);

AO21x1_ASAP7_75t_L g821 ( 
.A1(n_655),
.A2(n_731),
.B(n_739),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_664),
.B(n_665),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_674),
.B(n_614),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_645),
.B(n_723),
.Y(n_824)
);

AO31x2_ASAP7_75t_L g825 ( 
.A1(n_655),
.A2(n_677),
.A3(n_678),
.B(n_694),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_718),
.B(n_535),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_664),
.B(n_665),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_644),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_664),
.A2(n_655),
.B(n_665),
.C(n_568),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_SL g830 ( 
.A1(n_744),
.A2(n_655),
.B(n_719),
.C(n_684),
.Y(n_830)
);

CKINVDCx11_ASAP7_75t_R g831 ( 
.A(n_723),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_685),
.B(n_490),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_664),
.A2(n_655),
.B(n_665),
.C(n_568),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_665),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_664),
.B(n_665),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_653),
.A2(n_687),
.B(n_680),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_664),
.A2(n_655),
.B(n_665),
.C(n_568),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_664),
.A2(n_655),
.B(n_665),
.C(n_568),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_655),
.A2(n_648),
.B(n_664),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_664),
.A2(n_655),
.B(n_665),
.C(n_568),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_655),
.A2(n_648),
.B(n_664),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_692),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_801),
.B(n_808),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_822),
.B(n_827),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_813),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_773),
.B(n_786),
.Y(n_846)
);

AO21x2_ASAP7_75t_L g847 ( 
.A1(n_797),
.A2(n_836),
.B(n_819),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_754),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_834),
.B(n_835),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_SL g850 ( 
.A1(n_829),
.A2(n_840),
.B(n_838),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_832),
.B(n_764),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_785),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_837),
.A2(n_766),
.B(n_760),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_765),
.B(n_811),
.Y(n_854)
);

AO21x2_ASAP7_75t_L g855 ( 
.A1(n_821),
.A2(n_767),
.B(n_839),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_800),
.B(n_779),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_810),
.B(n_826),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

NOR2x1_ASAP7_75t_L g859 ( 
.A(n_817),
.B(n_761),
.Y(n_859)
);

AOI221xp5_ASAP7_75t_L g860 ( 
.A1(n_802),
.A2(n_814),
.B1(n_806),
.B2(n_812),
.C(n_841),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_792),
.A2(n_828),
.B1(n_751),
.B2(n_771),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_785),
.B(n_745),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_758),
.B(n_759),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_780),
.A2(n_750),
.B(n_787),
.C(n_789),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_SL g866 ( 
.A1(n_746),
.A2(n_769),
.B(n_823),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_763),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_770),
.A2(n_796),
.B(n_782),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_791),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_804),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_805),
.A2(n_795),
.B(n_799),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_774),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_784),
.B(n_762),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_778),
.B(n_749),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_756),
.A2(n_820),
.B(n_747),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_790),
.A2(n_794),
.B(n_748),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_798),
.A2(n_783),
.B1(n_791),
.B2(n_755),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_793),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_772),
.B(n_775),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_772),
.B(n_775),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_807),
.A2(n_815),
.A3(n_825),
.B(n_818),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_757),
.B(n_777),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_824),
.B(n_815),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_831),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_815),
.B(n_825),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_753),
.A2(n_816),
.B(n_818),
.Y(n_886)
);

OAI221xp5_ASAP7_75t_L g887 ( 
.A1(n_781),
.A2(n_776),
.B1(n_816),
.B2(n_818),
.C(n_768),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_776),
.A2(n_781),
.B(n_768),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_788),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_781),
.B(n_776),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_768),
.A2(n_833),
.B(n_829),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_788),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_801),
.B(n_808),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_842),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_754),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_801),
.B(n_808),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_773),
.B(n_786),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_803),
.B(n_645),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_801),
.B(n_808),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_801),
.B(n_808),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_761),
.B(n_645),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_SL g902 ( 
.A(n_777),
.B(n_718),
.Y(n_902)
);

AO31x2_ASAP7_75t_L g903 ( 
.A1(n_821),
.A2(n_766),
.A3(n_756),
.B(n_767),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_801),
.B(n_808),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_832),
.B(n_685),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_809),
.A2(n_830),
.B(n_655),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_829),
.A2(n_837),
.B(n_833),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_832),
.B(n_685),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_801),
.B(n_808),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_802),
.A2(n_814),
.B(n_806),
.C(n_808),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_829),
.A2(n_837),
.B(n_833),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_854),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_870),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_854),
.B(n_867),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_857),
.B(n_858),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_846),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_SL g917 ( 
.A1(n_873),
.A2(n_883),
.B(n_860),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_SL g918 ( 
.A1(n_877),
.A2(n_873),
.B(n_865),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_894),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_852),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_846),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_897),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_906),
.A2(n_853),
.B(n_886),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_907),
.B(n_911),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_843),
.B(n_844),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_849),
.B(n_893),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_897),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_872),
.A2(n_856),
.B1(n_851),
.B2(n_863),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_845),
.B(n_849),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_877),
.B(n_850),
.Y(n_932)
);

OAI21x1_ASAP7_75t_SL g933 ( 
.A1(n_907),
.A2(n_911),
.B(n_909),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_893),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_896),
.B(n_909),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_896),
.B(n_900),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_899),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_910),
.B(n_852),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_869),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_892),
.B(n_875),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_900),
.B(n_904),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_889),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_848),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_885),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_878),
.B(n_908),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_891),
.A2(n_888),
.B(n_887),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_855),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_905),
.B(n_890),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_890),
.B(n_881),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_859),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_903),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_869),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_890),
.B(n_881),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_895),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_875),
.B(n_903),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_903),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_895),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_942),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_922),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_882),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_926),
.B(n_892),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_938),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_938),
.Y(n_963)
);

OAI22xp33_ASAP7_75t_L g964 ( 
.A1(n_932),
.A2(n_902),
.B1(n_901),
.B2(n_884),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_948),
.B(n_861),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_940),
.B(n_847),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_926),
.B(n_949),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_932),
.A2(n_902),
.B1(n_874),
.B2(n_901),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_944),
.B(n_876),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_944),
.B(n_879),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_949),
.B(n_868),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_953),
.B(n_956),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_953),
.B(n_871),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_913),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_914),
.B(n_880),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_914),
.B(n_898),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_946),
.B(n_866),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_936),
.B(n_901),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_912),
.B(n_928),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_922),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_951),
.B(n_884),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_941),
.B(n_934),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_916),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_947),
.B(n_955),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_972),
.B(n_932),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_972),
.B(n_932),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_932),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_966),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_982),
.B(n_931),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_931),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_959),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_958),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_958),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_979),
.B(n_941),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_967),
.B(n_925),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_966),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_967),
.B(n_925),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_967),
.B(n_961),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_961),
.B(n_925),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_961),
.B(n_925),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_979),
.B(n_937),
.Y(n_1001)
);

NAND2xp67_ASAP7_75t_L g1002 ( 
.A(n_981),
.B(n_977),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_975),
.B(n_937),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_992),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_995),
.B(n_973),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_995),
.B(n_973),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_969),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_997),
.B(n_999),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_973),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_985),
.A2(n_964),
.B1(n_977),
.B2(n_981),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_989),
.B(n_981),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_994),
.B(n_984),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_990),
.B(n_977),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1000),
.B(n_971),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_992),
.Y(n_1015)
);

AOI32xp33_ASAP7_75t_L g1016 ( 
.A1(n_998),
.A2(n_964),
.A3(n_968),
.B1(n_954),
.B2(n_957),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_993),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_998),
.B(n_984),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_988),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1000),
.B(n_984),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_985),
.B(n_986),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_985),
.B(n_971),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_1013),
.B(n_943),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_1016),
.A2(n_950),
.B(n_915),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1004),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1004),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_1020),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1010),
.A2(n_983),
.B1(n_1018),
.B2(n_978),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1020),
.B(n_988),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_1007),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1008),
.B(n_1014),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1015),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1008),
.B(n_988),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_1001),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1014),
.B(n_996),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1012),
.B(n_917),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1036),
.B(n_1005),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_1028),
.A2(n_930),
.B1(n_917),
.B2(n_978),
.C(n_1003),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_1030),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1040)
);

OR4x1_ASAP7_75t_L g1041 ( 
.A(n_1027),
.B(n_991),
.C(n_950),
.D(n_1017),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_1027),
.A2(n_1002),
.B(n_1022),
.Y(n_1042)
);

AOI322xp5_ASAP7_75t_L g1043 ( 
.A1(n_1031),
.A2(n_1006),
.A3(n_1005),
.B1(n_1009),
.B2(n_1022),
.C1(n_983),
.C2(n_1021),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1024),
.A2(n_986),
.B1(n_987),
.B2(n_1021),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1029),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1032),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_1033),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1029),
.A2(n_991),
.B(n_918),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_1039),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1038),
.A2(n_1044),
.B1(n_1042),
.B2(n_1037),
.Y(n_1050)
);

OAI211xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1043),
.A2(n_1023),
.B(n_918),
.C(n_965),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_1038),
.A2(n_1034),
.B1(n_1035),
.B2(n_1033),
.C(n_1032),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1037),
.B(n_1009),
.Y(n_1054)
);

AOI221x1_ASAP7_75t_L g1055 ( 
.A1(n_1048),
.A2(n_1025),
.B1(n_1026),
.B2(n_1019),
.C(n_933),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_1051),
.A2(n_976),
.B(n_965),
.C(n_1047),
.Y(n_1056)
);

OAI211xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1052),
.A2(n_1050),
.B(n_1053),
.C(n_1054),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1049),
.B(n_1041),
.Y(n_1058)
);

AOI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_1057),
.A2(n_1045),
.B1(n_1035),
.B2(n_1026),
.C(n_962),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1056),
.B(n_1055),
.C(n_963),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_1060),
.B(n_1058),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_974),
.C(n_921),
.Y(n_1062)
);

XNOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1061),
.B(n_976),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1062),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_1064),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1065),
.Y(n_1068)
);

XNOR2xp5_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_945),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1067),
.A2(n_963),
.B1(n_962),
.B2(n_1019),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1068),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_1006),
.Y(n_1072)
);

NAND2x1_ASAP7_75t_L g1073 ( 
.A(n_1067),
.B(n_921),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1071),
.A2(n_1073),
.B(n_1070),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1072),
.A2(n_924),
.B(n_929),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1071),
.Y(n_1076)
);

OAI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1071),
.A2(n_923),
.B(n_945),
.C(n_952),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1071),
.A2(n_952),
.B1(n_939),
.B2(n_919),
.C(n_920),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1071),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1076),
.A2(n_927),
.B(n_935),
.Y(n_1080)
);

OAI222xp33_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_980),
.B1(n_960),
.B2(n_975),
.C1(n_970),
.C2(n_928),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1074),
.A2(n_927),
.B(n_935),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_1078),
.B1(n_1077),
.B2(n_1075),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_SL g1084 ( 
.A1(n_1083),
.A2(n_1080),
.B1(n_1081),
.B2(n_952),
.Y(n_1084)
);


endmodule