module fake_jpeg_30830_n_451 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_51),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_53),
.B(n_94),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_55),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_8),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_8),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_8),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_20),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_91),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_95),
.Y(n_122)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_97),
.B1(n_33),
.B2(n_41),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_110),
.B1(n_118),
.B2(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_24),
.C(n_35),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_105),
.B(n_142),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_47),
.B1(n_45),
.B2(n_42),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_69),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_33),
.B1(n_36),
.B2(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_129),
.B1(n_133),
.B2(n_135),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_36),
.B1(n_40),
.B2(n_35),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_84),
.A2(n_47),
.B1(n_45),
.B2(n_42),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_22),
.B1(n_21),
.B2(n_27),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_54),
.A2(n_29),
.B(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_94),
.B1(n_41),
.B2(n_55),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_34),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_43),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_153),
.B(n_162),
.Y(n_232)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_76),
.B1(n_66),
.B2(n_74),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_100),
.B1(n_147),
.B2(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_36),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_34),
.B1(n_24),
.B2(n_19),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_172),
.B1(n_173),
.B2(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_170),
.Y(n_209)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_33),
.B1(n_62),
.B2(n_85),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_183),
.B1(n_188),
.B2(n_191),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_32),
.B1(n_43),
.B2(n_57),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_43),
.B1(n_95),
.B2(n_51),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_104),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_190),
.Y(n_213)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_103),
.A2(n_93),
.B1(n_91),
.B2(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_108),
.A2(n_43),
.B1(n_97),
.B2(n_96),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_195),
.B(n_196),
.Y(n_221)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_116),
.A2(n_146),
.A3(n_124),
.B1(n_128),
.B2(n_151),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_43),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_104),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_41),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_194),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_197),
.B1(n_140),
.B2(n_132),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_198),
.A2(n_224),
.B1(n_174),
.B2(n_196),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_147),
.B(n_150),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_206),
.B(n_220),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_118),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_165),
.C(n_192),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_127),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_163),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_112),
.B(n_123),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_153),
.B(n_138),
.CI(n_102),
.CON(n_207),
.SN(n_207)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_178),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_125),
.B1(n_119),
.B2(n_144),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_218),
.B1(n_160),
.B2(n_154),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_125),
.B1(n_144),
.B2(n_132),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_112),
.B(n_138),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_138),
.B(n_140),
.C(n_115),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_230),
.B(n_174),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_162),
.A2(n_9),
.B(n_14),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_187),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_236),
.Y(n_268)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_182),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_237),
.B(n_245),
.C(n_253),
.Y(n_289)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_252),
.B(n_256),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_175),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_216),
.B1(n_228),
.B2(n_217),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_178),
.B1(n_197),
.B2(n_188),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_259),
.B1(n_220),
.B2(n_208),
.Y(n_272)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_177),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_250),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_191),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_176),
.C(n_156),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_215),
.Y(n_255)
);

AO21x2_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_215),
.B(n_231),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_191),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_264),
.B(n_199),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_169),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_221),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_164),
.B1(n_157),
.B2(n_158),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_0),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_223),
.B(n_203),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_199),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_218),
.A3(n_207),
.B1(n_229),
.B2(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_274),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_246),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_276),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_205),
.B1(n_203),
.B2(n_207),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_205),
.B1(n_203),
.B2(n_229),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_283),
.B1(n_286),
.B2(n_288),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_284),
.B(n_287),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_237),
.A2(n_209),
.B1(n_227),
.B2(n_210),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_212),
.B(n_222),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_227),
.B1(n_201),
.B2(n_233),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_242),
.A2(n_233),
.B1(n_225),
.B2(n_201),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_252),
.A2(n_215),
.B(n_212),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_225),
.B1(n_219),
.B2(n_222),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_219),
.B1(n_212),
.B2(n_215),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_246),
.Y(n_304)
);

XOR2x2_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_253),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_295),
.B(n_282),
.Y(n_342)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_264),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_311),
.B(n_9),
.Y(n_348)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_307),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_241),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_308),
.A2(n_267),
.B1(n_272),
.B2(n_273),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_280),
.A2(n_246),
.B1(n_262),
.B2(n_260),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_309),
.A2(n_319),
.B1(n_291),
.B2(n_285),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_258),
.B(n_257),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_313),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_268),
.B(n_250),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_236),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_316),
.B(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_318),
.Y(n_347)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_263),
.B1(n_244),
.B2(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_261),
.B1(n_238),
.B2(n_249),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_289),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_334),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_324),
.A2(n_327),
.B1(n_340),
.B2(n_305),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_289),
.C(n_283),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_332),
.C(n_339),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_310),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_328),
.A2(n_344),
.B1(n_298),
.B2(n_311),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_348),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_296),
.A2(n_287),
.B1(n_290),
.B2(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_276),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_342),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_290),
.C(n_263),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_263),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_298),
.A2(n_308),
.B(n_310),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_335),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_288),
.B1(n_282),
.B2(n_279),
.Y(n_336)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_279),
.C(n_235),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_282),
.B1(n_248),
.B2(n_235),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_282),
.B1(n_248),
.B2(n_255),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_282),
.C(n_1),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_319),
.C(n_297),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g351 ( 
.A1(n_338),
.A2(n_303),
.B(n_307),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_364),
.Y(n_378)
);

XOR2x2_ASAP7_75t_SL g352 ( 
.A(n_331),
.B(n_303),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_357),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_341),
.B(n_314),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_365),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_367),
.B1(n_340),
.B2(n_324),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_294),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_362),
.C(n_366),
.Y(n_377)
);

XOR2x2_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_309),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_294),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_321),
.B1(n_320),
.B2(n_302),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_327),
.A2(n_317),
.B1(n_315),
.B2(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_371),
.B(n_346),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_348),
.B1(n_343),
.B2(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_342),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_387),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_339),
.C(n_347),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_385),
.C(n_388),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_384),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_347),
.C(n_335),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_351),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_389),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_344),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_337),
.C(n_333),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_360),
.B(n_333),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_337),
.Y(n_390)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_L g391 ( 
.A1(n_373),
.A2(n_358),
.B1(n_354),
.B2(n_371),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_391),
.A2(n_7),
.B1(n_14),
.B2(n_3),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_393),
.B(n_12),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_367),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_402),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_361),
.C(n_366),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_400),
.C(n_405),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_364),
.C(n_362),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_352),
.B1(n_370),
.B2(n_3),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_377),
.A2(n_370),
.B(n_9),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_404),
.B(n_3),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_387),
.C(n_375),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_405),
.B(n_375),
.CI(n_379),
.CON(n_408),
.SN(n_408)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_404),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_394),
.A2(n_378),
.B(n_12),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_409),
.B(n_410),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_0),
.C(n_1),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_414),
.B1(n_14),
.B2(n_15),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_395),
.C(n_400),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_416),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_0),
.C(n_1),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_418),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_397),
.B(n_3),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_403),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_419),
.A2(n_421),
.B(n_408),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_425),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_401),
.Y(n_422)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_422),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_412),
.A2(n_396),
.B1(n_399),
.B2(n_391),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_390),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_426),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_392),
.Y(n_427)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_411),
.A2(n_396),
.B1(n_6),
.B2(n_13),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_417),
.C(n_418),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_429),
.C(n_424),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_407),
.B(n_410),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_436),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_422),
.A2(n_408),
.B(n_416),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_435),
.B(n_0),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_427),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_439),
.A2(n_441),
.B(n_431),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_442),
.B(n_436),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_433),
.A2(n_423),
.B(n_15),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_443),
.A2(n_0),
.B(n_1),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_432),
.C(n_437),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_444),
.B(n_445),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_447),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_446),
.C(n_1),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);


endmodule