module fake_netlist_6_4435_n_1192 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1192);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1192;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_208;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_168;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_1101;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_1119;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_167;
wire n_631;
wire n_174;
wire n_720;
wire n_758;
wire n_153;
wire n_842;
wire n_525;
wire n_1163;
wire n_516;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_156;
wire n_1168;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_953;
wire n_448;
wire n_1017;
wire n_1094;
wire n_1004;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_196;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_1084;
wire n_929;
wire n_460;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_163;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_265;
wire n_260;
wire n_313;
wire n_624;
wire n_451;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_556;
wire n_159;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_1053;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_195;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_834;
wire n_207;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_165;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_663;
wire n_508;
wire n_856;
wire n_1050;
wire n_379;
wire n_170;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_169;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

INVx1_ASAP7_75t_L g153 ( 
.A(n_10),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_85),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_27),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_53),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_23),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_55),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_67),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_65),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_48),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_25),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_101),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_103),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_89),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_113),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_75),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_50),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_59),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_2),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_63),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_116),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_73),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_31),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_12),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_152),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_45),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_155),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_174),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_154),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_176),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_234),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_214),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_231),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_219),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_232),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_215),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_224),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_224),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_216),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_216),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_226),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_251),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_257),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_246),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_291),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

BUFx2_ASAP7_75t_SL g322 ( 
.A(n_292),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_286),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_246),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_291),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_248),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_248),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_254),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_300),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_303),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_324),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_309),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_267),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_311),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_320),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_320),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_268),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_266),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_317),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_337),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_306),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_310),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_322),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_332),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_314),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_336),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_260),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_367),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_335),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_354),
.A2(n_319),
.B1(n_336),
.B2(n_339),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_339),
.B1(n_271),
.B2(n_274),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_339),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_312),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_289),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_289),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_349),
.B(n_266),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_376),
.A2(n_307),
.B(n_305),
.Y(n_416)
);

AOI22x1_ASAP7_75t_SL g417 ( 
.A1(n_350),
.A2(n_260),
.B1(n_164),
.B2(n_352),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_304),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_354),
.B(n_288),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_368),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_354),
.B(n_288),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

CKINVDCx6p67_ASAP7_75t_R g434 ( 
.A(n_356),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_354),
.A2(n_166),
.B1(n_169),
.B2(n_284),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_289),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_350),
.A2(n_270),
.B1(n_169),
.B2(n_166),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_312),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_354),
.B(n_313),
.Y(n_444)
);

BUFx8_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_304),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_340),
.B(n_313),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

CKINVDCx6p67_ASAP7_75t_R g449 ( 
.A(n_356),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_347),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_340),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_318),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_340),
.A2(n_307),
.B(n_305),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_344),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_354),
.B(n_318),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_453),
.Y(n_464)
);

BUFx8_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_455),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_386),
.B(n_414),
.Y(n_467)
);

AND3x2_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_157),
.C(n_282),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_283),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_321),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_321),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_297),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_436),
.C(n_438),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_297),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_285),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_308),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_270),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

NAND2x1_ASAP7_75t_L g495 ( 
.A(n_388),
.B(n_293),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_308),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_457),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_380),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_294),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_163),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

AND3x2_ASAP7_75t_L g504 ( 
.A(n_415),
.B(n_204),
.C(n_180),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_407),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_315),
.Y(n_509)
);

AND3x2_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_204),
.C(n_187),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_432),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_407),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_R g520 ( 
.A(n_506),
.B(n_450),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_484),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_465),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_506),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_484),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_518),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_465),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_518),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_465),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_503),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_471),
.B(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_503),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_503),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_467),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_492),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_515),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_486),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_499),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_492),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_507),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_471),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_511),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_515),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_515),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_474),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_464),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_502),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_496),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_485),
.B(n_434),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_474),
.B(n_480),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_546),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_525),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_548),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_549),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_556),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_534),
.B(n_481),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_521),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_542),
.B(n_400),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_551),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_530),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_550),
.B(n_392),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_522),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_390),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

INVx4_ASAP7_75t_SL g578 ( 
.A(n_528),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_521),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_532),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_539),
.Y(n_583)
);

XOR2x2_ASAP7_75t_SL g584 ( 
.A(n_547),
.B(n_441),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_520),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_522),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_R g589 ( 
.A(n_524),
.B(n_417),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_547),
.A2(n_410),
.B1(n_423),
.B2(n_445),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_554),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_544),
.Y(n_593)
);

AOI22x1_ASAP7_75t_L g594 ( 
.A1(n_557),
.A2(n_397),
.B1(n_395),
.B2(n_512),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_522),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_525),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_527),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_554),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_472),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_560),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_540),
.A2(n_414),
.B1(n_418),
.B2(n_421),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_541),
.B(n_483),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_540),
.B(n_422),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_462),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_545),
.B(n_418),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_553),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_545),
.B(n_391),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_528),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_528),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_523),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_537),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_559),
.B(n_463),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_536),
.B(n_390),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_469),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_549),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g623 ( 
.A1(n_534),
.A2(n_410),
.B1(n_423),
.B2(n_445),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_534),
.B(n_404),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_549),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_534),
.B(n_404),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_534),
.B(n_404),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_534),
.A2(n_421),
.B1(n_408),
.B2(n_412),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_546),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_534),
.B(n_404),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_534),
.B(n_411),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_473),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_534),
.B(n_411),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_534),
.B(n_458),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_546),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_534),
.B(n_405),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_546),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_534),
.B(n_405),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_540),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_549),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_633),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_567),
.B(n_458),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_598),
.Y(n_644)
);

AO22x2_ASAP7_75t_L g645 ( 
.A1(n_567),
.A2(n_412),
.B1(n_421),
.B2(n_475),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_561),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_564),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_416),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_571),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_607),
.B(n_416),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_624),
.B(n_426),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_635),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_637),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_613),
.B(n_505),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_573),
.A2(n_468),
.B1(n_163),
.B2(n_206),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_632),
.Y(n_659)
);

AND3x1_ASAP7_75t_L g660 ( 
.A(n_618),
.B(n_424),
.C(n_402),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_574),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_634),
.B(n_476),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_582),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_572),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_570),
.B(n_405),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_598),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_634),
.B(n_476),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_563),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_626),
.B(n_482),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_SL g672 ( 
.A1(n_627),
.A2(n_416),
.B1(n_420),
.B2(n_424),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_613),
.B(n_612),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_612),
.B(n_505),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_572),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_563),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_569),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_569),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_578),
.B(n_479),
.Y(n_679)
);

AOI22x1_ASAP7_75t_L g680 ( 
.A1(n_617),
.A2(n_425),
.B1(n_409),
.B2(n_406),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_565),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_580),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_578),
.B(n_488),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_579),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_579),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_581),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_621),
.B(n_426),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_570),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_610),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_578),
.B(n_491),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_630),
.B(n_482),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_636),
.B(n_426),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_580),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_566),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_574),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_568),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_638),
.B(n_623),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_640),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_573),
.A2(n_519),
.B1(n_517),
.B2(n_501),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_588),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_609),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_SL g705 ( 
.A(n_614),
.B(n_405),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_587),
.B(n_406),
.Y(n_706)
);

AND2x2_ASAP7_75t_SL g707 ( 
.A(n_575),
.B(n_406),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_568),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_602),
.B(n_493),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_605),
.B(n_406),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_612),
.B(n_426),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_611),
.A2(n_489),
.B1(n_480),
.B2(n_474),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_588),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_588),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_439),
.B1(n_443),
.B2(n_440),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_625),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_602),
.B(n_494),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_625),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_581),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_601),
.B(n_498),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_587),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_679),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_647),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_653),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_654),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_646),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_657),
.B(n_590),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_649),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_659),
.B(n_599),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_689),
.B(n_599),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_663),
.B(n_640),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_643),
.B(n_705),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_666),
.Y(n_734)
);

AO21x2_ASAP7_75t_L g735 ( 
.A1(n_702),
.A2(n_611),
.B(n_597),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_643),
.B(n_705),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_690),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_652),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_658),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_697),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_663),
.B(n_585),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_675),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_642),
.B(n_609),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_669),
.B(n_585),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_656),
.A2(n_575),
.B1(n_606),
.B2(n_608),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_662),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_651),
.B(n_423),
.Y(n_747)
);

OAI221xp5_ASAP7_75t_L g748 ( 
.A1(n_656),
.A2(n_603),
.B1(n_591),
.B2(n_600),
.C(n_639),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_698),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_700),
.A2(n_615),
.B1(n_619),
.B2(n_618),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_697),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_593),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_667),
.B(n_604),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_665),
.Y(n_754)
);

CKINVDCx14_ASAP7_75t_R g755 ( 
.A(n_644),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_651),
.A2(n_620),
.B1(n_617),
.B2(n_615),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_695),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_695),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_704),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_669),
.B(n_583),
.Y(n_760)
);

BUFx4f_ASAP7_75t_L g761 ( 
.A(n_697),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_677),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_679),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_701),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_668),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_684),
.B(n_595),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_703),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_688),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_703),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_703),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_667),
.B(n_596),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_667),
.B(n_616),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_701),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_693),
.A2(n_620),
.B1(n_396),
.B2(n_618),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_702),
.B(n_680),
.C(n_660),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_672),
.B(n_594),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_671),
.B(n_586),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_670),
.Y(n_779)
);

INVx4_ASAP7_75t_SL g780 ( 
.A(n_673),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_685),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_715),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_668),
.Y(n_783)
);

INVx5_ASAP7_75t_L g784 ( 
.A(n_711),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_686),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_676),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_681),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_722),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_693),
.B(n_423),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_671),
.B(n_562),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_683),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_687),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_696),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_715),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_743),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_783),
.B(n_710),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_769),
.B(n_682),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_753),
.B(n_694),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_724),
.B(n_672),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_745),
.B(n_660),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_788),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_727),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_748),
.B(n_706),
.C(n_396),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_745),
.B(n_707),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_729),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_776),
.B(n_413),
.Y(n_807)
);

NOR2x1p5_ASAP7_75t_L g808 ( 
.A(n_776),
.B(n_616),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_738),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_725),
.B(n_648),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_739),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_765),
.B(n_756),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_726),
.B(n_650),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_756),
.B(n_584),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_752),
.B(n_692),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_748),
.A2(n_419),
.B1(n_645),
.B2(n_711),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_752),
.B(n_692),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_777),
.B(n_645),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_749),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_759),
.B(n_419),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_764),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_754),
.Y(n_824)
);

OAI221xp5_ASAP7_75t_L g825 ( 
.A1(n_750),
.A2(n_712),
.B1(n_711),
.B2(n_589),
.C(n_459),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_779),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_733),
.A2(n_614),
.B1(n_390),
.B2(n_712),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_723),
.B(n_763),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_728),
.B(n_708),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_786),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_766),
.B(n_413),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_728),
.B(n_713),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_773),
.B(n_614),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_777),
.A2(n_775),
.B1(n_736),
.B2(n_747),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_787),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_740),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_731),
.B(n_790),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_723),
.B(n_584),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_766),
.B(n_413),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_740),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_734),
.B(n_383),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_789),
.B(n_383),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_763),
.B(n_684),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_791),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_790),
.B(n_717),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_773),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_730),
.B(n_719),
.Y(n_848)
);

CKINVDCx11_ASAP7_75t_R g849 ( 
.A(n_742),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_793),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_775),
.A2(n_167),
.B(n_189),
.C(n_188),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_780),
.B(n_691),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_730),
.B(n_720),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_753),
.B(n_641),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_SL g855 ( 
.A(n_735),
.B(n_413),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_778),
.B(n_721),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_778),
.B(n_721),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_795),
.B(n_760),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_762),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_784),
.A2(n_201),
.B(n_203),
.C(n_198),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_757),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_780),
.B(n_691),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_755),
.B(n_434),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_768),
.B(n_449),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_760),
.B(n_673),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_758),
.B(n_641),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_740),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_751),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_751),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_768),
.B(n_449),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_751),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_784),
.B(n_766),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_774),
.B(n_673),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_834),
.B(n_784),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_829),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_835),
.B(n_772),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_867),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_849),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_796),
.B(n_393),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_835),
.B(n_772),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_803),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_867),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_838),
.B(n_735),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_801),
.A2(n_741),
.B(n_732),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_802),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_804),
.A2(n_766),
.B1(n_673),
.B2(n_674),
.Y(n_886)
);

AND2x6_ASAP7_75t_SL g887 ( 
.A(n_863),
.B(n_842),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_823),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_806),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_814),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_816),
.B(n_767),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_815),
.A2(n_761),
.B(n_782),
.C(n_393),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_818),
.B(n_856),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_857),
.B(n_781),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_809),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_858),
.B(n_865),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_826),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_800),
.B(n_853),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_805),
.A2(n_782),
.B1(n_761),
.B2(n_741),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_845),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_861),
.B(n_732),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_847),
.B(n_785),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_847),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_848),
.B(n_792),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_808),
.A2(n_183),
.B1(n_206),
.B2(n_163),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_821),
.B(n_872),
.Y(n_906)
);

NOR2x1_ASAP7_75t_R g907 ( 
.A(n_839),
.B(n_454),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_850),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_812),
.A2(n_744),
.B(n_718),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_817),
.A2(n_744),
.B1(n_709),
.B2(n_718),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_811),
.B(n_794),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_819),
.B(n_770),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_831),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_846),
.B(n_770),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_802),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_802),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_807),
.A2(n_709),
.B(n_716),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_872),
.B(n_771),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_797),
.B(n_771),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_854),
.B(n_799),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_828),
.B(n_715),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_798),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_836),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_866),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_874),
.A2(n_840),
.B(n_832),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_888),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_899),
.A2(n_825),
.B1(n_820),
.B2(n_855),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_884),
.A2(n_851),
.B(n_860),
.C(n_864),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_899),
.A2(n_862),
.B(n_852),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_906),
.A2(n_820),
.B(n_844),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_884),
.B(n_885),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_886),
.A2(n_827),
.B1(n_820),
.B2(n_843),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_881),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_898),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_876),
.A2(n_880),
.B(n_918),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_896),
.B(n_859),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_917),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_918),
.A2(n_873),
.B(n_833),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_905),
.A2(n_830),
.B(n_870),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_919),
.A2(n_813),
.B(n_810),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_907),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_883),
.B(n_837),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_892),
.A2(n_822),
.B(n_868),
.C(n_841),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_878),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_902),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_910),
.A2(n_871),
.B1(n_869),
.B2(n_867),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_875),
.B(n_661),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_893),
.B(n_661),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_885),
.B(n_871),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_922),
.A2(n_716),
.B(n_592),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_920),
.A2(n_674),
.B1(n_183),
.B2(n_206),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_910),
.A2(n_714),
.B(n_664),
.C(n_195),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_903),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_916),
.B(n_674),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_925),
.B(n_664),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_909),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_901),
.A2(n_592),
.B(n_401),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_894),
.B(n_911),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_901),
.A2(n_904),
.B(n_891),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_921),
.B(n_923),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_915),
.B(n_895),
.Y(n_962)
);

AOI21xp33_ASAP7_75t_L g963 ( 
.A1(n_879),
.A2(n_445),
.B(n_0),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_897),
.B(n_655),
.Y(n_964)
);

CKINVDCx10_ASAP7_75t_R g965 ( 
.A(n_887),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_900),
.B(n_655),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_890),
.B(n_588),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_908),
.B(n_655),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_912),
.A2(n_914),
.B(n_889),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_902),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_877),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_877),
.B(n_882),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_903),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_877),
.A2(n_882),
.B1(n_913),
.B2(n_924),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_899),
.A2(n_674),
.B1(n_655),
.B2(n_510),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_877),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_874),
.B(n_454),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_884),
.B(n_403),
.Y(n_978)
);

INVx11_ASAP7_75t_L g979 ( 
.A(n_878),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_936),
.A2(n_403),
.B(n_184),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_929),
.A2(n_158),
.B(n_480),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_976),
.Y(n_982)
);

OA22x2_ASAP7_75t_L g983 ( 
.A1(n_932),
.A2(n_504),
.B1(n_158),
.B2(n_178),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_928),
.A2(n_975),
.B1(n_930),
.B2(n_935),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_976),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_953),
.A2(n_399),
.B1(n_489),
.B2(n_496),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_927),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_965),
.B(n_0),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_976),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_926),
.B(n_496),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_960),
.B(n_1),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_939),
.B(n_1),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_938),
.Y(n_993)
);

AO31x2_ASAP7_75t_L g994 ( 
.A1(n_931),
.A2(n_2),
.A3(n_3),
.B(n_4),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_963),
.A2(n_447),
.B(n_489),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_959),
.B(n_3),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_978),
.A2(n_181),
.B(n_177),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_941),
.B(n_5),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_947),
.A2(n_495),
.B(n_514),
.C(n_448),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_934),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_1000),
.B(n_957),
.Y(n_1001)
);

INVx3_ASAP7_75t_SL g1002 ( 
.A(n_993),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_992),
.A2(n_944),
.B(n_942),
.C(n_933),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_984),
.B(n_977),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_980),
.A2(n_950),
.B(n_940),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_983),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_991),
.A2(n_969),
.B(n_970),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_998),
.A2(n_977),
.B1(n_952),
.B2(n_951),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_987),
.B(n_943),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_985),
.A2(n_954),
.B(n_973),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_985),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_981),
.A2(n_974),
.B1(n_958),
.B2(n_971),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_982),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_994),
.B(n_962),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_988),
.B(n_979),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_989),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_990),
.A2(n_972),
.B(n_948),
.C(n_966),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_994),
.B(n_946),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_996),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_994),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_997),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_997),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_986),
.A2(n_967),
.B(n_956),
.C(n_954),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_999),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_986),
.A2(n_972),
.B(n_968),
.C(n_964),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1022),
.A2(n_995),
.B(n_945),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_1002),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1005),
.A2(n_949),
.B(n_937),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_1006),
.B(n_961),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1011),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1016),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1013),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_1032),
.A2(n_1007),
.B(n_1010),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1033),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1033),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_1034),
.A2(n_1026),
.B(n_1020),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_1037),
.A2(n_1026),
.B(n_1031),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_1027),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1040),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1039),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_1042),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1041),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1043),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1044),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_1045),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1046),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_1048),
.A2(n_1039),
.B(n_1038),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_1047),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_1049),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1051),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1052),
.A2(n_1011),
.B1(n_1006),
.B2(n_1029),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_1051),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_1019),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_1019),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1058),
.B(n_1019),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_SL g1061 ( 
.A1(n_1059),
.A2(n_1057),
.B(n_1015),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_1060),
.B(n_1011),
.C(n_1003),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1061),
.B(n_1001),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1062),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1064),
.B(n_1001),
.C(n_1024),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1063),
.A2(n_1023),
.B1(n_1004),
.B2(n_1021),
.C(n_1014),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1065),
.B(n_1009),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1066),
.B(n_1018),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1068),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1070),
.A2(n_1008),
.B1(n_1028),
.B2(n_1012),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1070),
.B(n_1017),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1073),
.B(n_1025),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1072),
.B(n_5),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1071),
.B(n_1012),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1076),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1075),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_1074),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1078),
.A2(n_1008),
.B(n_6),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1079),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1080),
.B(n_7),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_7),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_1084),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1083),
.B(n_8),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_182),
.B(n_185),
.C(n_186),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1086),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1088),
.B(n_8),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1087),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1088),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_SL g1092 ( 
.A1(n_1091),
.A2(n_191),
.B(n_190),
.Y(n_1092)
);

AOI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_1090),
.A2(n_192),
.B(n_196),
.C(n_197),
.Y(n_1093)
);

AOI211xp5_ASAP7_75t_L g1094 ( 
.A1(n_1089),
.A2(n_200),
.B(n_202),
.C(n_207),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

BUFx4_ASAP7_75t_R g1096 ( 
.A(n_1092),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_1093),
.C(n_208),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_9),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_1097),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1098),
.A2(n_9),
.B(n_10),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1100),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1102),
.B(n_11),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_330),
.B(n_11),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1104),
.B(n_12),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_1103),
.B(n_509),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1106),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_13),
.C(n_14),
.Y(n_1108)
);

AO22x1_ASAP7_75t_L g1109 ( 
.A1(n_1105),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_1107),
.B(n_15),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1108),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_17),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_1111),
.B(n_18),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_1110),
.Y(n_1115)
);

NAND4xp75_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_19),
.C(n_20),
.D(n_21),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_1115),
.B(n_19),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_L g1119 ( 
.A(n_1117),
.B(n_20),
.C(n_21),
.Y(n_1119)
);

AOI211xp5_ASAP7_75t_SL g1120 ( 
.A1(n_1118),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_1119),
.B(n_1120),
.C(n_22),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_24),
.B(n_25),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_1121),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1123),
.B(n_26),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_1126)
);

NAND2x1_ASAP7_75t_L g1127 ( 
.A(n_1123),
.B(n_30),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1126),
.B(n_509),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1125),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1130),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1128),
.A2(n_456),
.B1(n_451),
.B2(n_509),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_SL g1135 ( 
.A1(n_1133),
.A2(n_1129),
.B1(n_33),
.B2(n_34),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1134),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1136),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1135),
.A2(n_508),
.B1(n_487),
.B2(n_478),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1137),
.A2(n_461),
.B1(n_508),
.B2(n_487),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1140),
.B(n_461),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

XNOR2xp5_ASAP7_75t_L g1143 ( 
.A(n_1140),
.B(n_32),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1141),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_35),
.B(n_36),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1142),
.A2(n_37),
.B(n_38),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1144),
.A2(n_39),
.B(n_41),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1145),
.B(n_477),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1146),
.A2(n_42),
.B(n_43),
.Y(n_1150)
);

AOI22x1_ASAP7_75t_L g1151 ( 
.A1(n_1147),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1150),
.A2(n_49),
.B(n_51),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

AOI222xp33_ASAP7_75t_L g1154 ( 
.A1(n_1149),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.C1(n_57),
.C2(n_58),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1148),
.A2(n_61),
.B(n_62),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1150),
.A2(n_508),
.B1(n_487),
.B2(n_478),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1150),
.A2(n_64),
.B(n_66),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1150),
.A2(n_508),
.B1(n_487),
.B2(n_478),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1150),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1150),
.B(n_68),
.Y(n_1160)
);

OAI22x1_ASAP7_75t_SL g1161 ( 
.A1(n_1150),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_1161)
);

AOI222xp33_ASAP7_75t_L g1162 ( 
.A1(n_1150),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.C1(n_80),
.C2(n_81),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1150),
.B(n_82),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1159),
.A2(n_83),
.B(n_84),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1153),
.A2(n_86),
.B(n_88),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1153),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1163),
.B(n_91),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1156),
.A2(n_955),
.B1(n_478),
.B2(n_477),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1158),
.A2(n_92),
.B(n_93),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1160),
.A2(n_94),
.B(n_95),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_L g1171 ( 
.A(n_1152),
.B(n_96),
.C(n_97),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1157),
.A2(n_98),
.B(n_100),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1166),
.A2(n_1155),
.B1(n_1161),
.B2(n_1162),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1171),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1167),
.B(n_1154),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1172),
.A2(n_1169),
.B1(n_1164),
.B2(n_1170),
.Y(n_1176)
);

XNOR2xp5_ASAP7_75t_L g1177 ( 
.A(n_1165),
.B(n_102),
.Y(n_1177)
);

XNOR2xp5_ASAP7_75t_L g1178 ( 
.A(n_1168),
.B(n_104),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1166),
.A2(n_477),
.B1(n_106),
.B2(n_107),
.Y(n_1179)
);

AOI222xp33_ASAP7_75t_L g1180 ( 
.A1(n_1174),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.C1(n_111),
.C2(n_112),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1175),
.A2(n_955),
.B1(n_477),
.B2(n_516),
.Y(n_1181)
);

XOR2x2_ASAP7_75t_L g1182 ( 
.A(n_1173),
.B(n_114),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1176),
.A2(n_115),
.B(n_118),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1182),
.B(n_1177),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_1178),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1185),
.A2(n_1183),
.B1(n_1179),
.B2(n_1180),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1186),
.B(n_1181),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1187),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.C(n_122),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1188),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.C(n_128),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1189),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1190)
);

AOI211xp5_ASAP7_75t_L g1191 ( 
.A1(n_1190),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_1191)
);

AOI211xp5_ASAP7_75t_L g1192 ( 
.A1(n_1191),
.A2(n_136),
.B(n_137),
.C(n_139),
.Y(n_1192)
);


endmodule