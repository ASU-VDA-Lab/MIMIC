module fake_netlist_1_397_n_31 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
CKINVDCx8_ASAP7_75t_R g16 ( .A(n_5), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_13), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_11), .B(n_0), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_6), .B(n_8), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_0), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_1), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_17), .B1(n_16), .B2(n_19), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_20), .B(n_24), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_27), .B(n_1), .Y(n_29) );
AO22x2_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_2), .B1(n_3), .B2(n_7), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_18), .B1(n_28), .B2(n_10), .Y(n_31) );
endmodule