module fake_ibex_1206_n_906 (n_85, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_63, n_98, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_116, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_112, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_24, n_52, n_99, n_105, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_906);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_24;
input n_52;
input n_99;
input n_105;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_906;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_130;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_125;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_470;
wire n_339;
wire n_276;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_598;
wire n_825;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_127;
wire n_121;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_120;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_136;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_141;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_506;
wire n_562;
wire n_444;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_135;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_148;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_159;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_118),
.Y(n_123)
);

INVxp33_ASAP7_75t_SL g124 ( 
.A(n_19),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVxp33_ASAP7_75t_SL g126 ( 
.A(n_64),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVxp33_ASAP7_75t_SL g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_38),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_25),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_47),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_77),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_27),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_7),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_26),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_39),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_15),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_107),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_44),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_24),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_33),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_45),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_67),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_29),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_5),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_34),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_22),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_49),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_24),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_68),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_23),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_36),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_73),
.B(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_19),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_48),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_54),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_1),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_97),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_74),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

OR2x6_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_1),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_139),
.B(n_2),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_136),
.B(n_3),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_4),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_7),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_137),
.B(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_9),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_143),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_15),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_122),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_145),
.A2(n_62),
.B(n_115),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_160),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_132),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_142),
.B(n_16),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g259 ( 
.A(n_189),
.B(n_61),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_142),
.B(n_16),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_160),
.B(n_18),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_165),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_171),
.B(n_20),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_202),
.B(n_20),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_170),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_167),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_205),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_134),
.B(n_21),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_124),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_146),
.B(n_26),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_203),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_178),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_182),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_196),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_204),
.B(n_28),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_197),
.Y(n_291)
);

CKINVDCx6p67_ASAP7_75t_R g292 ( 
.A(n_167),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_200),
.B(n_131),
.Y(n_293)
);

OR2x2_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_150),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_274),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_214),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_281),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_214),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_238),
.B(n_120),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_214),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_213),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_159),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_259),
.B(n_181),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

NOR2x1p5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_127),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_180),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_213),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_213),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_210),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_211),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_219),
.B(n_120),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_168),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_224),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_247),
.B(n_148),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_212),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_240),
.A2(n_174),
.B1(n_207),
.B2(n_153),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_211),
.A2(n_181),
.B1(n_198),
.B2(n_169),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_253),
.B(n_140),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_283),
.B(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_212),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_217),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_259),
.B(n_187),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_259),
.A2(n_129),
.B1(n_126),
.B2(n_198),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_229),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_216),
.B(n_190),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_257),
.B(n_161),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_217),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_211),
.B(n_194),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_226),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_215),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_215),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_211),
.B(n_191),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_226),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_260),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_290),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_233),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_237),
.B(n_244),
.Y(n_357)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_279),
.B(n_239),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_218),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_229),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_218),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_293),
.B(n_195),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_222),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_243),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_222),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_237),
.B(n_209),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_225),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_229),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_229),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_256),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_262),
.B(n_199),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_244),
.B(n_173),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_240),
.A2(n_179),
.B1(n_162),
.B2(n_184),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_221),
.B(n_140),
.Y(n_374)
);

BUFx4f_ASAP7_75t_L g375 ( 
.A(n_287),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_256),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_283),
.B(n_149),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_221),
.B(n_161),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_221),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_223),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_221),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_245),
.B(n_201),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_231),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_265),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_256),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_245),
.B(n_129),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_246),
.B(n_149),
.Y(n_389)
);

AO21x2_ASAP7_75t_L g390 ( 
.A1(n_220),
.A2(n_206),
.B(n_155),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_246),
.B(n_166),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_265),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_262),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_270),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_262),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_248),
.B(n_126),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_270),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_249),
.B(n_151),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_275),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_287),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_275),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_283),
.B(n_154),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_249),
.Y(n_406)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g408 ( 
.A(n_353),
.B(n_248),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_353),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_R g413 ( 
.A(n_312),
.B(n_248),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_301),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_346),
.B(n_251),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_330),
.B(n_251),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_283),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_346),
.B(n_254),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_329),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_350),
.B(n_254),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

AND3x2_ASAP7_75t_SL g425 ( 
.A(n_315),
.B(n_174),
.C(n_207),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_310),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_310),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_284),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_356),
.B(n_284),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_337),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_329),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_327),
.Y(n_439)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_305),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_388),
.B(n_284),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_307),
.B(n_267),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_305),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_296),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_388),
.B(n_266),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_374),
.B(n_266),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_397),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_354),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_267),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_396),
.A2(n_248),
.B(n_241),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_297),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_297),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_396),
.A2(n_234),
.B(n_230),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_389),
.B(n_268),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_324),
.B(n_278),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_318),
.A2(n_268),
.B1(n_258),
.B2(n_288),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_362),
.B(n_258),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_306),
.B(n_264),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_317),
.B(n_277),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_311),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_311),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_333),
.B(n_280),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_318),
.B(n_255),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_357),
.B(n_255),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_362),
.B(n_285),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_344),
.B(n_278),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_325),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_325),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_373),
.B(n_289),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_309),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_352),
.B(n_273),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_295),
.B(n_264),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_273),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_325),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_364),
.B(n_343),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_298),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_391),
.B(n_285),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_298),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_340),
.A2(n_288),
.B1(n_286),
.B2(n_289),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_384),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_364),
.B(n_391),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_390),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

O2A1O1Ixp5_ASAP7_75t_L g494 ( 
.A1(n_402),
.A2(n_286),
.B(n_228),
.C(n_242),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_328),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_366),
.B(n_242),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_366),
.B(n_241),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_340),
.A2(n_291),
.B1(n_287),
.B2(n_250),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_299),
.Y(n_499)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_372),
.A2(n_398),
.B(n_313),
.Y(n_500)
);

CKINVDCx6p67_ASAP7_75t_R g501 ( 
.A(n_304),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_415),
.A2(n_355),
.B1(n_328),
.B2(n_358),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_358),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_420),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_421),
.A2(n_355),
.B1(n_328),
.B2(n_358),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_417),
.B(n_303),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_405),
.B(n_299),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_418),
.B(n_341),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_501),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_412),
.A2(n_410),
.B1(n_438),
.B2(n_421),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_412),
.A2(n_382),
.B1(n_308),
.B2(n_321),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_408),
.A2(n_314),
.B(n_316),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_436),
.B(n_312),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

AO31x2_ASAP7_75t_L g523 ( 
.A1(n_449),
.A2(n_322),
.A3(n_320),
.B(n_228),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_406),
.B(n_328),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_382),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_422),
.Y(n_526)
);

AOI221xp5_ASAP7_75t_L g527 ( 
.A1(n_437),
.A2(n_398),
.B1(n_372),
.B2(n_379),
.C(n_227),
.Y(n_527)
);

BUFx12f_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_429),
.B(n_328),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_479),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_490),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_405),
.B(n_402),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_493),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_437),
.B(n_379),
.Y(n_537)
);

OAI22x1_ASAP7_75t_L g538 ( 
.A1(n_425),
.A2(n_294),
.B1(n_123),
.B2(n_227),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_405),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_429),
.B(n_390),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_408),
.A2(n_395),
.B(n_348),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_412),
.B(n_232),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_232),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_439),
.B(n_491),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_481),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_476),
.A2(n_371),
.B1(n_367),
.B2(n_365),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_405),
.Y(n_550)
);

BUFx2_ASAP7_75t_SL g551 ( 
.A(n_407),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_451),
.B(n_395),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_480),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_481),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_432),
.B(n_371),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_414),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_463),
.B(n_383),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_463),
.B(n_383),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_460),
.B(n_381),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_460),
.B(n_381),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_464),
.A2(n_349),
.B(n_359),
.C(n_376),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_410),
.B(n_287),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_454),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_448),
.Y(n_567)
);

NAND2x2_ASAP7_75t_L g568 ( 
.A(n_425),
.B(n_291),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_407),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_454),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_453),
.A2(n_458),
.B(n_449),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_470),
.B(n_423),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_414),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_481),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_438),
.B(n_381),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_475),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_465),
.B(n_361),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_440),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_500),
.A2(n_230),
.B(n_234),
.C(n_250),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_478),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_489),
.A2(n_291),
.B1(n_363),
.B2(n_345),
.Y(n_585)
);

INVx8_ASAP7_75t_L g586 ( 
.A(n_407),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_488),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_478),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_484),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_452),
.A2(n_339),
.B(n_347),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_432),
.B(n_471),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_442),
.B(n_464),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_473),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_499),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_483),
.A2(n_351),
.B1(n_347),
.B2(n_345),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_407),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_452),
.A2(n_339),
.B(n_351),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_593),
.A2(n_487),
.B1(n_483),
.B2(n_462),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_469),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_522),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_592),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_513),
.A2(n_503),
.B1(n_572),
.B2(n_554),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_511),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_515),
.Y(n_606)
);

BUFx4f_ASAP7_75t_L g607 ( 
.A(n_528),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_469),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_508),
.B(n_469),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_591),
.B(n_473),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_430),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_543),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_503),
.A2(n_476),
.B1(n_447),
.B2(n_492),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_510),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_505),
.B(n_459),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_545),
.B(n_430),
.Y(n_619)
);

OA21x2_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_494),
.B(n_441),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_447),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_536),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_541),
.A2(n_441),
.B(n_487),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_530),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_504),
.A2(n_507),
.B1(n_542),
.B2(n_568),
.Y(n_626)
);

CKINVDCx11_ASAP7_75t_R g627 ( 
.A(n_542),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_524),
.B(n_430),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_459),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_506),
.A2(n_465),
.B1(n_413),
.B2(n_461),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_586),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_586),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_526),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_521),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_532),
.B(n_465),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_540),
.A2(n_472),
.B1(n_409),
.B2(n_411),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_587),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_506),
.A2(n_498),
.B1(n_470),
.B2(n_431),
.Y(n_642)
);

OAI222xp33_ASAP7_75t_L g643 ( 
.A1(n_517),
.A2(n_455),
.B1(n_450),
.B2(n_444),
.C1(n_424),
.C2(n_416),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_544),
.B(n_497),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_527),
.B(n_585),
.C(n_549),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_539),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_575),
.B(n_430),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_567),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_589),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_516),
.A2(n_497),
.B1(n_496),
.B2(n_291),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_537),
.A2(n_496),
.B1(n_291),
.B2(n_433),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_565),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_565),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_538),
.A2(n_494),
.B1(n_477),
.B2(n_443),
.C(n_403),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_581),
.B(n_440),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_546),
.B(n_478),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_539),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_546),
.A2(n_256),
.B1(n_272),
.B2(n_440),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_595),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_520),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_523),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_550),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_558),
.B(n_428),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_520),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_529),
.A2(n_519),
.B1(n_553),
.B2(n_561),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_555),
.A2(n_426),
.B1(n_256),
.B2(n_272),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_558),
.B(n_272),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_272),
.Y(n_670)
);

AOI21xp33_ASAP7_75t_L g671 ( 
.A1(n_556),
.A2(n_564),
.B(n_565),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_547),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_272),
.B1(n_263),
.B2(n_236),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_560),
.A2(n_236),
.B1(n_263),
.B2(n_375),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_523),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_523),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_561),
.A2(n_236),
.B1(n_263),
.B2(n_375),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_551),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_576),
.A2(n_236),
.B1(n_263),
.B2(n_446),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_559),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_531),
.Y(n_682)
);

AND2x2_ASAP7_75t_SL g683 ( 
.A(n_547),
.B(n_319),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_573),
.A2(n_319),
.B1(n_323),
.B2(n_400),
.Y(n_684)
);

OAI222xp33_ASAP7_75t_L g685 ( 
.A1(n_576),
.A2(n_378),
.B1(n_368),
.B2(n_360),
.C1(n_400),
.C2(n_377),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_550),
.B(n_323),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_578),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_585),
.A2(n_457),
.B1(n_456),
.B2(n_445),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_590),
.A2(n_377),
.B(n_378),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_569),
.B(n_319),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_547),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_569),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_598),
.A2(n_276),
.B1(n_282),
.B2(n_319),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_552),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_573),
.A2(n_323),
.B1(n_360),
.B2(n_368),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_531),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_534),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_583),
.A2(n_323),
.B(n_276),
.C(n_282),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_557),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_574),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_509),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_596),
.A2(n_282),
.B1(n_276),
.B2(n_369),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_509),
.A2(n_282),
.B1(n_276),
.B2(n_369),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_534),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_509),
.A2(n_282),
.B1(n_276),
.B2(n_369),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_636),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_646),
.A2(n_512),
.B(n_535),
.Y(n_709)
);

AOI211xp5_ASAP7_75t_L g710 ( 
.A1(n_630),
.A2(n_535),
.B(n_512),
.C(n_582),
.Y(n_710)
);

AND2x4_ASAP7_75t_SL g711 ( 
.A(n_608),
.B(n_566),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_611),
.B(n_621),
.Y(n_712)
);

CKINVDCx8_ASAP7_75t_R g713 ( 
.A(n_634),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_621),
.A2(n_599),
.B1(n_594),
.B2(n_566),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_629),
.A2(n_582),
.B1(n_509),
.B2(n_597),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_SL g716 ( 
.A1(n_608),
.A2(n_597),
.B1(n_552),
.B2(n_570),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_636),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_608),
.A2(n_552),
.B1(n_566),
.B2(n_570),
.Y(n_718)
);

OA21x2_ASAP7_75t_L g719 ( 
.A1(n_700),
.A2(n_387),
.B(n_370),
.Y(n_719)
);

AOI221xp5_ASAP7_75t_L g720 ( 
.A1(n_603),
.A2(n_588),
.B1(n_584),
.B2(n_577),
.C(n_387),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_633),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_629),
.A2(n_588),
.B1(n_584),
.B2(n_577),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_636),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_661),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_604),
.A2(n_588),
.B1(n_584),
.B2(n_577),
.C(n_570),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_618),
.Y(n_726)
);

OAI221xp5_ASAP7_75t_L g727 ( 
.A1(n_604),
.A2(n_387),
.B1(n_370),
.B2(n_369),
.C(n_342),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_630),
.A2(n_601),
.B1(n_610),
.B2(n_615),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_644),
.B(n_387),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_615),
.B(n_370),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_653),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_602),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_627),
.A2(n_370),
.B1(n_342),
.B2(n_331),
.Y(n_733)
);

OAI211xp5_ASAP7_75t_SL g734 ( 
.A1(n_625),
.A2(n_342),
.B(n_331),
.C(n_35),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_616),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_651),
.A2(n_342),
.B1(n_331),
.B2(n_41),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_627),
.A2(n_331),
.B1(n_31),
.B2(n_42),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_638),
.A2(n_30),
.B1(n_43),
.B2(n_50),
.C(n_52),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_637),
.A2(n_53),
.B1(n_57),
.B2(n_59),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_633),
.Y(n_740)
);

OAI211xp5_ASAP7_75t_L g741 ( 
.A1(n_626),
.A2(n_63),
.B(n_69),
.C(n_70),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_614),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_613),
.B(n_641),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_600),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_651),
.A2(n_82),
.B1(n_86),
.B2(n_98),
.C(n_100),
.Y(n_746)
);

OAI33xp33_ASAP7_75t_L g747 ( 
.A1(n_663),
.A2(n_101),
.A3(n_104),
.B1(n_106),
.B2(n_109),
.B3(n_117),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_643),
.A2(n_635),
.B1(n_631),
.B2(n_645),
.C(n_650),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_607),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_640),
.A2(n_642),
.B1(n_622),
.B2(n_606),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_636),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_670),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_676),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_694),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_677),
.B(n_687),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_679),
.A2(n_607),
.B1(n_656),
.B2(n_639),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_640),
.B(n_697),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_605),
.B(n_609),
.Y(n_758)
);

OAI21xp33_ASAP7_75t_L g759 ( 
.A1(n_652),
.A2(n_626),
.B(n_655),
.Y(n_759)
);

OAI211xp5_ASAP7_75t_L g760 ( 
.A1(n_652),
.A2(n_657),
.B(n_678),
.C(n_674),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_681),
.B(n_653),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_624),
.A2(n_671),
.B1(n_667),
.B2(n_649),
.C(n_704),
.Y(n_762)
);

OAI222xp33_ASAP7_75t_L g763 ( 
.A1(n_660),
.A2(n_707),
.B1(n_705),
.B2(n_703),
.C1(n_667),
.C2(n_692),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

OAI221xp5_ASAP7_75t_L g765 ( 
.A1(n_673),
.A2(n_665),
.B1(n_660),
.B2(n_674),
.C(n_678),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_654),
.A2(n_696),
.B1(n_682),
.B2(n_699),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_706),
.A2(n_659),
.B1(n_664),
.B2(n_647),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_647),
.A2(n_664),
.B1(n_659),
.B2(n_692),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_L g769 ( 
.A1(n_623),
.A2(n_632),
.B1(n_675),
.B2(n_612),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_694),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_675),
.A2(n_683),
.B1(n_704),
.B2(n_623),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_700),
.A2(n_693),
.B(n_668),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_632),
.A2(n_683),
.B1(n_658),
.B2(n_628),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_628),
.B(n_619),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_612),
.A2(n_619),
.B1(n_666),
.B2(n_691),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_694),
.Y(n_776)
);

OAI221xp5_ASAP7_75t_L g777 ( 
.A1(n_673),
.A2(n_684),
.B1(n_707),
.B2(n_705),
.C(n_689),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_648),
.A2(n_620),
.B1(n_702),
.B2(n_701),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_620),
.B(n_666),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_620),
.B(n_648),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_780),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_755),
.B(n_698),
.Y(n_782)
);

OAI211xp5_ASAP7_75t_SL g783 ( 
.A1(n_732),
.A2(n_684),
.B(n_695),
.C(n_693),
.Y(n_783)
);

OAI221xp5_ASAP7_75t_L g784 ( 
.A1(n_750),
.A2(n_680),
.B1(n_688),
.B2(n_686),
.C(n_690),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_712),
.A2(n_728),
.B1(n_757),
.B2(n_759),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_SL g786 ( 
.A(n_749),
.B(n_686),
.C(n_690),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_712),
.B(n_662),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_740),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_763),
.A2(n_685),
.B(n_694),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_779),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_765),
.A2(n_662),
.B1(n_672),
.B2(n_691),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_743),
.B(n_672),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_755),
.B(n_658),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_777),
.A2(n_658),
.B1(n_773),
.B2(n_714),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_724),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_719),
.A2(n_658),
.B(n_771),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_724),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_L g798 ( 
.A1(n_748),
.A2(n_658),
.B1(n_726),
.B2(n_762),
.C(n_760),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_SL g799 ( 
.A1(n_756),
.A2(n_718),
.B(n_716),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_745),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_745),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_776),
.B(n_757),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_725),
.A2(n_715),
.B1(n_731),
.B2(n_768),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_779),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_SL g806 ( 
.A(n_749),
.B(n_713),
.C(n_710),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_709),
.B(n_753),
.C(n_738),
.Y(n_807)
);

BUFx2_ASAP7_75t_SL g808 ( 
.A(n_713),
.Y(n_808)
);

AO21x1_ASAP7_75t_L g809 ( 
.A1(n_736),
.A2(n_739),
.B(n_769),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_743),
.B(n_758),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_758),
.B(n_740),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_761),
.B(n_752),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_727),
.A2(n_720),
.B(n_734),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_778),
.B(n_766),
.C(n_741),
.Y(n_814)
);

OAI222xp33_ASAP7_75t_L g815 ( 
.A1(n_731),
.A2(n_746),
.B1(n_744),
.B2(n_761),
.C1(n_721),
.C2(n_775),
.Y(n_815)
);

AOI33xp33_ASAP7_75t_L g816 ( 
.A1(n_767),
.A2(n_730),
.A3(n_711),
.B1(n_737),
.B2(n_722),
.B3(n_764),
.Y(n_816)
);

OA21x2_ASAP7_75t_L g817 ( 
.A1(n_780),
.A2(n_730),
.B(n_751),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_721),
.A2(n_711),
.B1(n_733),
.B2(n_774),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_729),
.C(n_719),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_721),
.B(n_776),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_708),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_781),
.B(n_776),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_803),
.B(n_708),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_788),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_803),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_820),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_814),
.B(n_717),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_810),
.B(n_785),
.Y(n_828)
);

OAI33xp33_ASAP7_75t_L g829 ( 
.A1(n_802),
.A2(n_747),
.A3(n_751),
.B1(n_723),
.B2(n_717),
.B3(n_754),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_781),
.B(n_723),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_819),
.A2(n_772),
.B(n_754),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_790),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_797),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_808),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_800),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_790),
.B(n_805),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_801),
.Y(n_838)
);

NAND4xp25_ASAP7_75t_L g839 ( 
.A(n_785),
.B(n_770),
.C(n_772),
.D(n_719),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_805),
.B(n_770),
.Y(n_840)
);

OAI33xp33_ASAP7_75t_L g841 ( 
.A1(n_794),
.A2(n_772),
.A3(n_811),
.B1(n_812),
.B2(n_804),
.B3(n_787),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_L g842 ( 
.A1(n_799),
.A2(n_798),
.B1(n_807),
.B2(n_784),
.C(n_806),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_810),
.B(n_803),
.Y(n_843)
);

OAI33xp33_ASAP7_75t_L g844 ( 
.A1(n_782),
.A2(n_818),
.A3(n_783),
.B1(n_791),
.B2(n_793),
.B3(n_821),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_817),
.B(n_803),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_782),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_832),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_827),
.B(n_816),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_845),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_845),
.B(n_796),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_832),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_833),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_835),
.B(n_792),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_833),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_842),
.A2(n_793),
.B1(n_789),
.B2(n_792),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_837),
.B(n_817),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_837),
.B(n_817),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_834),
.Y(n_858)
);

OA211x2_ASAP7_75t_L g859 ( 
.A1(n_848),
.A2(n_786),
.B(n_828),
.C(n_841),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_848),
.A2(n_843),
.B1(n_826),
.B2(n_846),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_847),
.B(n_824),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_856),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_849),
.B(n_833),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_851),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_853),
.B(n_822),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_849),
.B(n_831),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_858),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_855),
.A2(n_844),
.B1(n_826),
.B2(n_825),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_852),
.Y(n_869)
);

NAND2x1_ASAP7_75t_L g870 ( 
.A(n_865),
.B(n_849),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_862),
.B(n_825),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_857),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_861),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_860),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_864),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_868),
.B(n_850),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_859),
.A2(n_850),
.B1(n_827),
.B2(n_843),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_867),
.Y(n_878)
);

CKINVDCx14_ASAP7_75t_R g879 ( 
.A(n_873),
.Y(n_879)
);

NOR4xp25_ASAP7_75t_L g880 ( 
.A(n_874),
.B(n_839),
.C(n_836),
.D(n_838),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_875),
.B(n_863),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_876),
.B(n_839),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_872),
.B(n_856),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_871),
.Y(n_884)
);

XNOR2xp5_ASAP7_75t_L g885 ( 
.A(n_877),
.B(n_863),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_878),
.B(n_869),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_SL g887 ( 
.A(n_870),
.B(n_816),
.C(n_809),
.Y(n_887)
);

XOR2x2_ASAP7_75t_L g888 ( 
.A(n_879),
.B(n_871),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_SL g889 ( 
.A1(n_884),
.A2(n_850),
.B1(n_866),
.B2(n_857),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_880),
.A2(n_866),
.B1(n_838),
.B2(n_836),
.C(n_834),
.Y(n_890)
);

AOI221xp5_ASAP7_75t_L g891 ( 
.A1(n_887),
.A2(n_881),
.B1(n_885),
.B2(n_886),
.C(n_883),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_869),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_892),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_891),
.A2(n_882),
.B(n_822),
.Y(n_894)
);

OAI221xp5_ASAP7_75t_L g895 ( 
.A1(n_889),
.A2(n_854),
.B1(n_852),
.B2(n_813),
.C(n_820),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_894),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_897),
.B(n_896),
.C(n_895),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_897),
.A2(n_888),
.B1(n_890),
.B2(n_809),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_SL g900 ( 
.A1(n_899),
.A2(n_898),
.B1(n_823),
.B2(n_815),
.Y(n_900)
);

OA22x2_ASAP7_75t_L g901 ( 
.A1(n_899),
.A2(n_823),
.B1(n_830),
.B2(n_854),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_900),
.A2(n_823),
.B1(n_829),
.B2(n_831),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_901),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_903),
.Y(n_904)
);

XNOR2xp5_ASAP7_75t_L g905 ( 
.A(n_904),
.B(n_902),
.Y(n_905)
);

OAI221xp5_ASAP7_75t_L g906 ( 
.A1(n_905),
.A2(n_821),
.B1(n_830),
.B2(n_840),
.C(n_831),
.Y(n_906)
);


endmodule