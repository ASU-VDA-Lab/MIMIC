module fake_jpeg_12190_n_646 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_646);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_646;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_63),
.B(n_86),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_66),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_8),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_75),
.B(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_31),
.B(n_8),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_77),
.B(n_82),
.Y(n_153)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_31),
.B(n_10),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_85),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_7),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_87),
.B(n_92),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_96),
.B(n_100),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_98),
.B(n_101),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_58),
.Y(n_148)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_117),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_108),
.Y(n_164)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_17),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_6),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_123),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_54),
.Y(n_120)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_32),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_124),
.B(n_126),
.Y(n_224)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_81),
.B1(n_114),
.B2(n_105),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_125),
.A2(n_24),
.B(n_25),
.C(n_36),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_129),
.B(n_131),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_49),
.B1(n_38),
.B2(n_57),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_130),
.A2(n_162),
.B1(n_171),
.B2(n_193),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_SL g131 ( 
.A(n_62),
.B(n_58),
.C(n_53),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_57),
.C(n_38),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_44),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_137),
.B(n_138),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_44),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_83),
.A2(n_28),
.B1(n_52),
.B2(n_19),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_142),
.A2(n_169),
.B1(n_185),
.B2(n_24),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_148),
.B(n_152),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_151),
.B(n_154),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_60),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_21),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_96),
.A2(n_49),
.B1(n_38),
.B2(n_41),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_163),
.B(n_196),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_46),
.B1(n_53),
.B2(n_52),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_100),
.A2(n_49),
.B1(n_52),
.B2(n_19),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_67),
.B(n_18),
.C(n_52),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_61),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_64),
.A2(n_19),
.B1(n_28),
.B2(n_55),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g246 ( 
.A1(n_190),
.A2(n_199),
.B1(n_200),
.B2(n_30),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_100),
.A2(n_28),
.B1(n_22),
.B2(n_55),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_74),
.A2(n_22),
.B1(n_51),
.B2(n_35),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_173),
.B1(n_147),
.B2(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_69),
.B(n_48),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_62),
.B(n_35),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_198),
.B(n_0),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_70),
.A2(n_43),
.B1(n_39),
.B2(n_25),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_71),
.A2(n_43),
.B1(n_39),
.B2(n_25),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_80),
.B(n_39),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_201),
.B(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_88),
.B1(n_123),
.B2(n_118),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_205),
.A2(n_181),
.B(n_139),
.Y(n_341)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_206),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_207),
.A2(n_263),
.B(n_181),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_124),
.A2(n_79),
.A3(n_89),
.B1(n_110),
.B2(n_107),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_212),
.B(n_191),
.CI(n_172),
.CON(n_323),
.SN(n_323)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_78),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_213),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_168),
.B(n_73),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_214),
.B(n_227),
.Y(n_295)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_216),
.Y(n_340)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_217),
.Y(n_339)
);

OR2x2_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_36),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_219),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_223),
.B(n_254),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_226),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_32),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_32),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_230),
.B(n_233),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_129),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_259),
.Y(n_282)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_161),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_234),
.A2(n_240),
.B1(n_241),
.B2(n_251),
.Y(n_293)
);

BUFx12_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_235),
.Y(n_287)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_142),
.A2(n_99),
.B1(n_97),
.B2(n_24),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_36),
.B1(n_89),
.B2(n_79),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

INVx6_ASAP7_75t_SL g245 ( 
.A(n_141),
.Y(n_245)
);

INVx11_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_246),
.A2(n_160),
.B1(n_128),
.B2(n_192),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_164),
.B(n_30),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_247),
.B(n_250),
.C(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_164),
.B(n_30),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_93),
.B1(n_14),
.B2(n_17),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_137),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_253),
.A2(n_156),
.B1(n_146),
.B2(n_172),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_134),
.B(n_6),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_126),
.B(n_13),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_256),
.B(n_265),
.Y(n_317)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_258),
.Y(n_338)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

BUFx16f_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_262),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_165),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_261),
.Y(n_304)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_138),
.A2(n_106),
.B1(n_94),
.B2(n_15),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_151),
.B(n_14),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_178),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_267),
.B(n_268),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_154),
.B(n_125),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_0),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_279),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_273),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_147),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_275),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_167),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_277),
.Y(n_336)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_278),
.Y(n_314)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_210),
.A2(n_128),
.B1(n_160),
.B2(n_192),
.Y(n_280)
);

AO21x2_ASAP7_75t_L g378 ( 
.A1(n_280),
.A2(n_306),
.B(n_307),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_224),
.B(n_132),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_283),
.B(n_312),
.C(n_325),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_182),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_299),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_297),
.A2(n_316),
.B1(n_324),
.B2(n_240),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_199),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_189),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_303),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_149),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_210),
.A2(n_197),
.B1(n_183),
.B2(n_180),
.Y(n_306)
);

AO22x2_ASAP7_75t_L g307 ( 
.A1(n_246),
.A2(n_207),
.B1(n_213),
.B2(n_241),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_186),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_197),
.B1(n_183),
.B2(n_180),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_332),
.B1(n_337),
.B2(n_248),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_341),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_213),
.A2(n_179),
.B1(n_166),
.B2(n_177),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_177),
.C(n_176),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_234),
.A2(n_179),
.B1(n_166),
.B2(n_176),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_250),
.B(n_149),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_343),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_225),
.B(n_139),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_342),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_253),
.B(n_0),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_250),
.B(n_181),
.C(n_15),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_330),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_345),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_348),
.Y(n_434)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_352),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_239),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_353),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_242),
.Y(n_352)
);

AO22x1_ASAP7_75t_SL g353 ( 
.A1(n_285),
.A2(n_307),
.B1(n_293),
.B2(n_303),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_308),
.A2(n_274),
.B1(n_206),
.B2(n_218),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_313),
.B(n_283),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_358),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_385),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_293),
.A2(n_270),
.B1(n_251),
.B2(n_205),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_357),
.A2(n_362),
.B1(n_374),
.B2(n_388),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_245),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_330),
.Y(n_360)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_289),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_364),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_270),
.B1(n_266),
.B2(n_259),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_286),
.B(n_222),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_365),
.B(n_369),
.Y(n_426)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_279),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_370),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_219),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_373),
.C(n_281),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_282),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_286),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_291),
.Y(n_372)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_312),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_285),
.A2(n_258),
.B1(n_238),
.B2(n_232),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_302),
.A2(n_236),
.B(n_235),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_375),
.A2(n_382),
.B(n_345),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_221),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_377),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_292),
.B(n_217),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_292),
.B(n_318),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_386),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_301),
.B(n_278),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_389),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_261),
.B(n_215),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_297),
.A2(n_299),
.B1(n_307),
.B2(n_323),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_390),
.B1(n_393),
.B2(n_379),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_320),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_276),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_294),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_307),
.A2(n_211),
.B1(n_273),
.B2(n_216),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_305),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_307),
.A2(n_209),
.B1(n_262),
.B2(n_277),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_281),
.B(n_1),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_294),
.Y(n_392)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_323),
.A2(n_208),
.B1(n_260),
.B2(n_3),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_396),
.A2(n_406),
.B1(n_284),
.B2(n_314),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_399),
.C(n_409),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_398),
.B(n_403),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_373),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_358),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_384),
.A2(n_321),
.B1(n_341),
.B2(n_325),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_355),
.B(n_334),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_407),
.B(n_317),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_343),
.C(n_333),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_333),
.C(n_328),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_416),
.C(n_418),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_320),
.B(n_304),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_365),
.B(n_389),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_327),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_327),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_421),
.Y(n_444)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_349),
.B(n_311),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_437),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_406),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_374),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_435),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_379),
.A2(n_393),
.B1(n_390),
.B2(n_369),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_433),
.A2(n_326),
.B(n_309),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_370),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_378),
.A2(n_317),
.B1(n_304),
.B2(n_329),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_436),
.A2(n_382),
.B1(n_348),
.B2(n_378),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_287),
.C(n_288),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_440),
.A2(n_466),
.B1(n_427),
.B2(n_420),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_441),
.A2(n_454),
.B(n_475),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_352),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_442),
.B(n_449),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_396),
.A2(n_378),
.B1(n_357),
.B2(n_353),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_446),
.A2(n_453),
.B1(n_455),
.B2(n_464),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_429),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_456),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_361),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_422),
.Y(n_450)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_450),
.Y(n_504)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

AOI322xp5_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_353),
.A3(n_378),
.B1(n_346),
.B2(n_367),
.C1(n_347),
.C2(n_381),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_473),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_434),
.A2(n_378),
.B1(n_388),
.B2(n_356),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_419),
.A2(n_353),
.B(n_346),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_433),
.A2(n_378),
.B1(n_347),
.B2(n_362),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_414),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_391),
.Y(n_458)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_458),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_392),
.Y(n_459)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_459),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_465),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_474),
.B(n_424),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_399),
.B(n_385),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_468),
.C(n_469),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_415),
.A2(n_382),
.B1(n_387),
.B2(n_340),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_400),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_382),
.B1(n_329),
.B2(n_340),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_311),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_397),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_404),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_437),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_472),
.A2(n_413),
.B1(n_395),
.B2(n_394),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_287),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_398),
.B(n_284),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_431),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_476),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_477),
.A2(n_480),
.B1(n_490),
.B2(n_498),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_440),
.A2(n_410),
.B1(n_424),
.B2(n_411),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_481),
.B(n_455),
.Y(n_527)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_484),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_407),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_494),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_412),
.Y(n_487)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_493),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_461),
.A2(n_454),
.B1(n_466),
.B2(n_447),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_491),
.B(n_499),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_412),
.Y(n_492)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_492),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_409),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_448),
.A2(n_410),
.B1(n_424),
.B2(n_427),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_438),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_446),
.A2(n_428),
.B1(n_423),
.B2(n_421),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_509),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_464),
.A2(n_413),
.B1(n_404),
.B2(n_408),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_502),
.A2(n_503),
.B1(n_444),
.B2(n_470),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_439),
.B(n_288),
.C(n_395),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_510),
.C(n_457),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_394),
.Y(n_507)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_507),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_408),
.C(n_338),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_456),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_442),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_514),
.B(n_520),
.C(n_521),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_516),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_462),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_518),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_443),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_443),
.C(n_468),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_471),
.C(n_474),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_522),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_463),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_523),
.B(n_533),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_475),
.B(n_453),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_524),
.A2(n_519),
.B(n_498),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_460),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_526),
.B(n_527),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_495),
.A2(n_465),
.B1(n_445),
.B2(n_444),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_529),
.A2(n_538),
.B1(n_501),
.B2(n_479),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_445),
.C(n_309),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_493),
.C(n_483),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_536),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_478),
.B(n_383),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_495),
.A2(n_502),
.B1(n_500),
.B2(n_505),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_535),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_481),
.B(n_338),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_508),
.A2(n_326),
.B1(n_359),
.B2(n_366),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_505),
.B(n_314),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_539),
.B(n_489),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_488),
.B(n_331),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_541),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_331),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_487),
.Y(n_542)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_542),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_492),
.Y(n_545)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_546),
.B(n_2),
.C(n_567),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_508),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_548),
.B(n_552),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_480),
.C(n_490),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_549),
.B(n_562),
.C(n_567),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_551),
.A2(n_524),
.B(n_531),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_507),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_555),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_483),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_526),
.B(n_489),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_556),
.B(n_563),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_484),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_558),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_560),
.A2(n_561),
.B1(n_564),
.B2(n_548),
.Y(n_572)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_503),
.C(n_504),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_515),
.B(n_504),
.Y(n_563)
);

INVx13_ASAP7_75t_L g564 ( 
.A(n_528),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_513),
.B(n_479),
.C(n_300),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_568),
.A2(n_569),
.B(n_573),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_553),
.A2(n_519),
.B(n_525),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_553),
.A2(n_525),
.B1(n_527),
.B2(n_521),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_570),
.A2(n_576),
.B1(n_584),
.B2(n_564),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_559),
.A2(n_530),
.B1(n_540),
.B2(n_538),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_571),
.A2(n_581),
.B1(n_557),
.B2(n_543),
.Y(n_605)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_572),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_551),
.A2(n_528),
.B(n_517),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_561),
.A2(n_513),
.B(n_518),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_574),
.A2(n_566),
.B(n_562),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_550),
.A2(n_536),
.B1(n_339),
.B2(n_275),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_587),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_560),
.A2(n_339),
.B1(n_260),
.B2(n_235),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_566),
.B(n_1),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_547),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_549),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_581)
);

FAx1_ASAP7_75t_SL g583 ( 
.A(n_554),
.B(n_2),
.CI(n_5),
.CON(n_583),
.SN(n_583)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_583),
.B(n_545),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_563),
.A2(n_2),
.B1(n_555),
.B2(n_558),
.Y(n_584)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_590),
.Y(n_607)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_585),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_591),
.B(n_593),
.Y(n_615)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_585),
.Y(n_593)
);

AOI21x1_ASAP7_75t_L g617 ( 
.A1(n_594),
.A2(n_599),
.B(n_582),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_550),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_595),
.B(n_597),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_546),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_596),
.B(n_604),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_565),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_543),
.C(n_544),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_598),
.B(n_600),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_568),
.A2(n_547),
.B(n_542),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_557),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_602),
.A2(n_571),
.B1(n_588),
.B2(n_581),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_577),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_603),
.A2(n_605),
.B1(n_570),
.B2(n_588),
.Y(n_610)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_578),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_579),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_586),
.C(n_544),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_608),
.B(n_612),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_618),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_610),
.B(n_617),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_574),
.C(n_587),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_616),
.B(n_608),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_602),
.A2(n_582),
.B1(n_577),
.B2(n_583),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_618),
.B(n_619),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_589),
.B(n_601),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_592),
.A2(n_576),
.B(n_583),
.C(n_600),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_620),
.A2(n_599),
.B(n_603),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_605),
.C(n_592),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_621),
.B(n_612),
.Y(n_627)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_622),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_615),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_623),
.B(n_630),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_621),
.A2(n_606),
.B(n_611),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_626),
.A2(n_613),
.B(n_620),
.Y(n_632)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_627),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_628),
.B(n_629),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_607),
.A2(n_614),
.B(n_610),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_632),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g635 ( 
.A(n_624),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g638 ( 
.A1(n_635),
.A2(n_634),
.B(n_625),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_638),
.Y(n_643)
);

AOI31xp67_ASAP7_75t_SL g640 ( 
.A1(n_636),
.A2(n_629),
.A3(n_628),
.B(n_617),
.Y(n_640)
);

BUFx24_ASAP7_75t_SL g642 ( 
.A(n_640),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_637),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_642),
.A2(n_641),
.B(n_639),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_644),
.A2(n_633),
.B(n_643),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_631),
.C(n_609),
.Y(n_646)
);


endmodule