module fake_jpeg_17059_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

AOI22xp33_ASAP7_75t_SL g7 ( 
.A1(n_0),
.A2(n_4),
.B1(n_3),
.B2(n_1),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_4),
.A2(n_0),
.B1(n_2),
.B2(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_0),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_1),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_1),
.C(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_14),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_13),
.B1(n_15),
.B2(n_11),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_7),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_6),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_6),
.B1(n_8),
.B2(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_12),
.B(n_17),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

AOI322xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_20),
.A3(n_22),
.B1(n_21),
.B2(n_18),
.C1(n_16),
.C2(n_19),
.Y(n_24)
);


endmodule