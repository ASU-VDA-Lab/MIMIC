module real_jpeg_16171_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_404),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_0),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

NAND2x1_ASAP7_75t_SL g136 ( 
.A(n_2),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_2),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_2),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_2),
.B(n_318),
.Y(n_317)
);

NAND2x1_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_81),
.Y(n_80)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_128),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_5),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_6),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_234),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_10),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_169),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_10),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_10),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_10),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_10),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_10),
.B(n_24),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_151),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_131),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_19),
.B(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.C(n_98),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_20),
.B(n_75),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_47),
.B1(n_48),
.B2(n_74),
.Y(n_20)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_22),
.B(n_37),
.C(n_41),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.C(n_30),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_23),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_126),
.C(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_23),
.A2(n_77),
.B1(n_78),
.B2(n_124),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_23),
.B(n_56),
.C(n_71),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_23),
.A2(n_124),
.B1(n_129),
.B2(n_147),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_107),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_25),
.A2(n_70),
.B1(n_71),
.B2(n_123),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_25),
.A2(n_71),
.B(n_176),
.C(n_238),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g347 ( 
.A1(n_25),
.A2(n_112),
.B1(n_113),
.B2(n_123),
.Y(n_347)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_33),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_40),
.Y(n_269)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_70),
.C(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_41),
.A2(n_46),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_41),
.A2(n_276),
.B(n_280),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_41),
.B(n_276),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_42),
.B(n_109),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_42),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_64),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_64),
.C(n_74),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_50),
.B(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_50),
.A2(n_127),
.B(n_233),
.Y(n_349)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_55),
.A2(n_56),
.B1(n_168),
.B2(n_172),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_55),
.A2(n_56),
.B1(n_145),
.B2(n_146),
.Y(n_293)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_67),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_70),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_59),
.C(n_141),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_R g231 ( 
.A1(n_56),
.A2(n_168),
.B(n_232),
.C(n_238),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_56),
.B(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_59),
.B(n_108),
.C(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_59),
.A2(n_60),
.B1(n_107),
.B2(n_108),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_59),
.A2(n_60),
.B1(n_267),
.B2(n_270),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_60),
.B(n_66),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_60),
.B(n_89),
.C(n_267),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_60),
.A2(n_65),
.B(n_73),
.Y(n_331)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_71),
.B1(n_80),
.B2(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_70),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_70),
.B(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_84),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_76),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_79),
.A2(n_84),
.B1(n_85),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_79),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_80),
.A2(n_127),
.B(n_171),
.Y(n_170)
);

NAND2x1p5_ASAP7_75t_L g171 ( 
.A(n_80),
.B(n_127),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_80),
.A2(n_105),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_83),
.Y(n_235)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_83),
.Y(n_305)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.C(n_92),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_87),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_86),
.A2(n_87),
.B1(n_191),
.B2(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_86),
.A2(n_87),
.B1(n_170),
.B2(n_173),
.Y(n_344)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_105),
.C(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_87),
.B(n_171),
.C(n_191),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_89),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_89),
.A2(n_119),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_89),
.B(n_129),
.C(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_99),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_120),
.C(n_125),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_101),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_116),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_102),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_106),
.B(n_116),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_107),
.A2(n_108),
.B1(n_191),
.B2(n_194),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_107),
.B(n_194),
.C(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2x2_ASAP7_75t_L g346 ( 
.A(n_108),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_119),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_120),
.B(n_125),
.Y(n_392)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_126),
.B(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_127),
.A2(n_221),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_127),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_127),
.B(n_233),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_127),
.A2(n_227),
.B1(n_233),
.B2(n_236),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_129),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_129),
.B(n_317),
.C(n_319),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_129),
.B(n_299),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_129),
.A2(n_147),
.B1(n_317),
.B2(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_149),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_148),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_143),
.B2(n_144),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_147),
.B(n_299),
.C(n_321),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_396),
.B(n_401),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_385),
.Y(n_152)
);

OAI321xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_311),
.A3(n_373),
.B1(n_378),
.B2(n_379),
.C(n_384),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_283),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_255),
.B(n_282),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_211),
.B(n_254),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_186),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_186),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.C(n_179),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_168),
.B(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_162),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_179),
.B1(n_180),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_176),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_176),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_183),
.A2(n_204),
.B1(n_266),
.B2(n_271),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_189),
.B(n_195),
.C(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_202),
.C(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_204),
.B(n_233),
.C(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_207),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_207),
.A2(n_210),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_207),
.B(n_300),
.C(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_220),
.B(n_221),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_229),
.B(n_253),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_216),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_225),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_225),
.B1(n_226),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_242),
.B(n_252),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_239),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_239),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_236),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_249),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_248),
.B(n_251),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_246),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_257),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_272),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_260),
.C(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_265),
.C(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_264),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_281),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_275),
.C(n_281),
.Y(n_310)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_284),
.B(n_285),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_296),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_297),
.C(n_310),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_292),
.C(n_294),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_310),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_306),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_308),
.C(n_309),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_361),
.Y(n_311)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_350),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_350),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_334),
.C(n_342),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_343),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_327),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_326),
.C(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.C(n_332),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_338),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_346),
.C(n_348),
.Y(n_356)
);

XOR2x1_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_353),
.C(n_355),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_358),
.C(n_360),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

AOI31xp67_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_374),
.A3(n_380),
.B(n_383),
.Y(n_379)
);

NAND2x1p5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_364),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.C(n_370),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_370),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_377),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_386),
.Y(n_385)
);

AND2x4_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_388),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_391),
.C(n_393),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_400),
.Y(n_403)
);


endmodule