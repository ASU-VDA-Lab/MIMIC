module real_aes_7738_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g459 ( .A(n_0), .Y(n_459) );
INVx1_ASAP7_75t_L g492 ( .A(n_1), .Y(n_492) );
INVx1_ASAP7_75t_L g201 ( .A(n_2), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_3), .A2(n_37), .B1(n_162), .B2(n_522), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g169 ( .A1(n_4), .A2(n_143), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_5), .B(n_136), .Y(n_505) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_8), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_8), .B(n_38), .Y(n_460) );
INVx1_ASAP7_75t_L g176 ( .A(n_9), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
INVx1_ASAP7_75t_L g486 ( .A(n_12), .Y(n_486) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_14), .B(n_184), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_15), .B(n_137), .Y(n_563) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_16), .A2(n_136), .A3(n_181), .B1(n_514), .B2(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_17), .A2(n_62), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_17), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_18), .B(n_162), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_19), .B(n_157), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_20), .B(n_137), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_50), .B1(n_162), .B2(n_522), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_22), .B(n_143), .Y(n_213) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_23), .A2(n_77), .B1(n_162), .B2(n_184), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_24), .B(n_162), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_25), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_26), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_28), .B(n_178), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_29), .B(n_174), .Y(n_203) );
INVx1_ASAP7_75t_L g190 ( .A(n_30), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_31), .A2(n_121), .B1(n_122), .B2(n_453), .Y(n_120) );
INVx1_ASAP7_75t_L g453 ( .A(n_31), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_32), .B(n_178), .Y(n_552) );
INVx2_ASAP7_75t_L g146 ( .A(n_33), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_34), .B(n_162), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_35), .B(n_178), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_36), .A2(n_148), .B(n_152), .C(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g109 ( .A(n_38), .Y(n_109) );
INVx1_ASAP7_75t_L g188 ( .A(n_39), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g766 ( .A1(n_40), .A2(n_767), .B1(n_770), .B2(n_771), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_40), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_41), .B(n_174), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_42), .B(n_162), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_43), .A2(n_88), .B1(n_220), .B2(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_44), .B(n_162), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_45), .B(n_162), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_46), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_47), .A2(n_70), .B1(n_768), .B2(n_769), .Y(n_767) );
CKINVDCx16_ASAP7_75t_R g769 ( .A(n_47), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_48), .B(n_491), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_49), .B(n_143), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_51), .A2(n_60), .B1(n_162), .B2(n_184), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_52), .A2(n_152), .B1(n_184), .B2(n_186), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_53), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_54), .B(n_162), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_55), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_56), .B(n_162), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_57), .A2(n_161), .B(n_173), .C(n_175), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_58), .Y(n_233) );
INVx1_ASAP7_75t_L g171 ( .A(n_59), .Y(n_171) );
INVx1_ASAP7_75t_L g149 ( .A(n_61), .Y(n_149) );
INVx1_ASAP7_75t_L g125 ( .A(n_62), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_63), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_64), .B(n_162), .Y(n_493) );
INVx1_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
AO32x2_ASAP7_75t_L g519 ( .A1(n_67), .A2(n_136), .A3(n_237), .B1(n_514), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g512 ( .A(n_68), .Y(n_512) );
INVx1_ASAP7_75t_L g547 ( .A(n_69), .Y(n_547) );
INVx1_ASAP7_75t_L g768 ( .A(n_70), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_SL g156 ( .A1(n_71), .A2(n_157), .B(n_158), .C(n_161), .Y(n_156) );
INVxp67_ASAP7_75t_L g159 ( .A(n_72), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_73), .B(n_184), .Y(n_548) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_75), .Y(n_194) );
INVx1_ASAP7_75t_L g226 ( .A(n_76), .Y(n_226) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_78), .A2(n_465), .B1(n_765), .B2(n_766), .C1(n_772), .C2(n_773), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_79), .A2(n_148), .B(n_152), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_80), .B(n_522), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_81), .B(n_184), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_82), .B(n_202), .Y(n_216) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_84), .B(n_157), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_85), .B(n_184), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_86), .A2(n_148), .B(n_152), .C(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
OR2x2_ASAP7_75t_L g456 ( .A(n_87), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g470 ( .A(n_87), .B(n_458), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_89), .A2(n_102), .B1(n_184), .B2(n_185), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_90), .A2(n_104), .B1(n_115), .B2(n_779), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_91), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_92), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_93), .A2(n_148), .B(n_152), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_94), .Y(n_247) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_96), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_97), .B(n_202), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_98), .B(n_184), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_99), .B(n_136), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_101), .A2(n_143), .B(n_150), .Y(n_142) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g780 ( .A(n_107), .Y(n_780) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g472 ( .A(n_111), .B(n_458), .Y(n_472) );
NOR2x2_ASAP7_75t_L g772 ( .A(n_111), .B(n_457), .Y(n_772) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B(n_463), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g778 ( .A(n_117), .Y(n_778) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_454), .B(n_461), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_127), .B2(n_452), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g452 ( .A(n_127), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_127), .A2(n_467), .B1(n_471), .B2(n_473), .Y(n_466) );
INVx1_ASAP7_75t_SL g775 ( .A(n_127), .Y(n_775) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND4x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_370), .C(n_417), .D(n_437), .Y(n_128) );
NOR3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_300), .C(n_325), .Y(n_129) );
OAI211xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_208), .B(n_260), .C(n_290), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_179), .Y(n_132) );
INVx3_ASAP7_75t_SL g342 ( .A(n_133), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_133), .B(n_273), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_133), .B(n_195), .Y(n_423) );
AND2x2_ASAP7_75t_L g446 ( .A(n_133), .B(n_312), .Y(n_446) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_167), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g264 ( .A(n_135), .B(n_168), .Y(n_264) );
INVx3_ASAP7_75t_L g277 ( .A(n_135), .Y(n_277) );
AND2x2_ASAP7_75t_L g282 ( .A(n_135), .B(n_167), .Y(n_282) );
OR2x2_ASAP7_75t_L g333 ( .A(n_135), .B(n_274), .Y(n_333) );
BUFx2_ASAP7_75t_L g353 ( .A(n_135), .Y(n_353) );
AND2x2_ASAP7_75t_L g363 ( .A(n_135), .B(n_274), .Y(n_363) );
AND2x2_ASAP7_75t_L g369 ( .A(n_135), .B(n_180), .Y(n_369) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_164), .Y(n_135) );
INVx4_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_136), .A2(n_498), .B(n_505), .Y(n_497) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_138), .B(n_139), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx2_ASAP7_75t_L g251 ( .A(n_143), .Y(n_251) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_144), .B(n_148), .Y(n_192) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g491 ( .A(n_145), .Y(n_491) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g153 ( .A(n_146), .Y(n_153) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx1_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
INVx1_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx4_ASAP7_75t_SL g163 ( .A(n_148), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_148), .A2(n_485), .B(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_148), .A2(n_499), .B(n_502), .Y(n_498) );
BUFx3_ASAP7_75t_L g514 ( .A(n_148), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_148), .A2(n_527), .B(n_531), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_148), .A2(n_546), .B(n_549), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B(n_156), .C(n_163), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_163), .B(n_171), .C(n_172), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_151), .A2(n_163), .B(n_253), .C(n_254), .Y(n_252) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
BUFx3_ASAP7_75t_L g220 ( .A(n_153), .Y(n_220) );
INVx1_ASAP7_75t_L g522 ( .A(n_153), .Y(n_522) );
INVx1_ASAP7_75t_L g530 ( .A(n_157), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_160), .B(n_176), .Y(n_175) );
INVx5_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_160), .A2(n_174), .B1(n_521), .B2(n_523), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_SL g546 ( .A1(n_161), .A2(n_202), .B(n_547), .C(n_548), .Y(n_546) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_162), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_163), .A2(n_183), .B1(n_191), .B2(n_192), .Y(n_182) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_165), .A2(n_169), .B(n_177), .Y(n_168) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_166), .B(n_223), .Y(n_222) );
AO21x1_ASAP7_75t_L g558 ( .A1(n_166), .A2(n_559), .B(n_562), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_166), .B(n_514), .C(n_559), .Y(n_577) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_168), .B(n_274), .Y(n_288) );
INVx2_ASAP7_75t_L g298 ( .A(n_168), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_168), .B(n_277), .Y(n_311) );
OR2x2_ASAP7_75t_L g322 ( .A(n_168), .B(n_274), .Y(n_322) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_168), .B(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g380 ( .A(n_168), .Y(n_380) );
AND2x2_ASAP7_75t_L g426 ( .A(n_168), .B(n_180), .Y(n_426) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_173), .A2(n_490), .B(n_512), .C(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_173), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_174), .A2(n_494), .B1(n_537), .B2(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_174), .A2(n_494), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g207 ( .A(n_178), .Y(n_207) );
INVx2_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_178), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_178), .A2(n_526), .B(n_534), .Y(n_525) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_178), .A2(n_545), .B(n_552), .Y(n_544) );
INVx3_ASAP7_75t_SL g299 ( .A(n_179), .Y(n_299) );
OR2x2_ASAP7_75t_L g352 ( .A(n_179), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
INVx3_ASAP7_75t_L g274 ( .A(n_180), .Y(n_274) );
AND2x2_ASAP7_75t_L g341 ( .A(n_180), .B(n_196), .Y(n_341) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_180), .Y(n_409) );
AOI33xp33_ASAP7_75t_L g413 ( .A1(n_180), .A2(n_342), .A3(n_349), .B1(n_358), .B2(n_414), .B3(n_415), .Y(n_413) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_193), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_181), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_181), .A2(n_197), .B(n_205), .Y(n_196) );
INVx2_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
INVx2_ASAP7_75t_L g204 ( .A(n_184), .Y(n_204) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g186 ( .A1(n_187), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_186) );
INVx2_ASAP7_75t_L g189 ( .A(n_187), .Y(n_189) );
INVx4_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_195), .B(n_277), .Y(n_276) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_195), .B(n_337), .C(n_339), .Y(n_336) );
AND2x2_ASAP7_75t_L g362 ( .A(n_195), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_195), .B(n_369), .Y(n_372) );
AND2x2_ASAP7_75t_L g425 ( .A(n_195), .B(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g281 ( .A(n_196), .Y(n_281) );
OR2x2_ASAP7_75t_L g375 ( .A(n_196), .B(n_274), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_204), .Y(n_200) );
INVx2_ASAP7_75t_L g494 ( .A(n_202), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_202), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_202), .A2(n_509), .B(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_204), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_207), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_207), .B(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_234), .Y(n_208) );
AOI32xp33_ASAP7_75t_L g326 ( .A1(n_209), .A2(n_327), .A3(n_329), .B1(n_331), .B2(n_334), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_209), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g429 ( .A(n_209), .Y(n_429) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g361 ( .A(n_210), .B(n_345), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_210), .B(n_307), .Y(n_381) );
AND2x2_ASAP7_75t_L g449 ( .A(n_210), .B(n_367), .Y(n_449) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
INVx3_ASAP7_75t_L g270 ( .A(n_211), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_211), .B(n_268), .Y(n_284) );
OR2x2_ASAP7_75t_L g289 ( .A(n_211), .B(n_267), .Y(n_289) );
INVx1_ASAP7_75t_L g296 ( .A(n_211), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_211), .B(n_278), .Y(n_304) );
AND2x2_ASAP7_75t_L g306 ( .A(n_211), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_211), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g359 ( .A(n_211), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_211), .B(n_444), .Y(n_443) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_214), .B(n_221), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_218), .A2(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
INVx1_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_221), .A2(n_484), .B(n_495), .Y(n_483) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_221), .A2(n_507), .B(n_515), .Y(n_506) );
INVx2_ASAP7_75t_L g268 ( .A(n_224), .Y(n_268) );
AND2x2_ASAP7_75t_L g314 ( .A(n_224), .B(n_235), .Y(n_314) );
AND2x2_ASAP7_75t_L g324 ( .A(n_224), .B(n_249), .Y(n_324) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_231), .B(n_232), .Y(n_224) );
INVx2_ASAP7_75t_L g444 ( .A(n_234), .Y(n_444) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_248), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_235), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
AND2x2_ASAP7_75t_L g329 ( .A(n_235), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g345 ( .A(n_235), .B(n_308), .Y(n_345) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
AND2x2_ASAP7_75t_L g307 ( .A(n_236), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g358 ( .A(n_236), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_236), .B(n_268), .Y(n_390) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
AND2x2_ASAP7_75t_L g269 ( .A(n_248), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g330 ( .A(n_248), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_248), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g367 ( .A(n_248), .Y(n_367) );
INVx1_ASAP7_75t_L g400 ( .A(n_248), .Y(n_400) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g278 ( .A(n_249), .B(n_268), .Y(n_278) );
INVx1_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g488 ( .A(n_255), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_255), .A2(n_550), .B(n_551), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_265), .B1(n_271), .B2(n_278), .C(n_279), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_262), .B(n_282), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_262), .B(n_345), .Y(n_422) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_264), .B(n_312), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_264), .B(n_273), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_264), .B(n_287), .Y(n_416) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g338 ( .A(n_268), .Y(n_338) );
AND2x2_ASAP7_75t_L g313 ( .A(n_269), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g391 ( .A(n_269), .Y(n_391) );
AND2x2_ASAP7_75t_L g323 ( .A(n_270), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_270), .B(n_293), .Y(n_339) );
AND2x2_ASAP7_75t_L g403 ( .A(n_270), .B(n_329), .Y(n_403) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g312 ( .A(n_274), .B(n_281), .Y(n_312) );
AND2x2_ASAP7_75t_L g408 ( .A(n_275), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_277), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_278), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_278), .B(n_285), .Y(n_373) );
AND2x2_ASAP7_75t_L g393 ( .A(n_278), .B(n_293), .Y(n_393) );
AND2x2_ASAP7_75t_L g414 ( .A(n_278), .B(n_358), .Y(n_414) );
OAI32xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_283), .A3(n_285), .B1(n_286), .B2(n_289), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_SL g287 ( .A(n_281), .Y(n_287) );
NAND2x1_ASAP7_75t_L g328 ( .A(n_281), .B(n_311), .Y(n_328) );
OR2x2_ASAP7_75t_L g332 ( .A(n_281), .B(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_281), .B(n_380), .Y(n_433) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_283), .A2(n_374), .B1(n_420), .B2(n_423), .C(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g334 ( .A(n_284), .B(n_307), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_284), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g412 ( .A(n_284), .B(n_345), .Y(n_412) );
INVxp67_ASAP7_75t_L g348 ( .A(n_285), .Y(n_348) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g418 ( .A(n_287), .B(n_405), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_287), .B(n_368), .Y(n_441) );
INVx1_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_289), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g434 ( .A(n_289), .B(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_294), .B(n_297), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_292), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g387 ( .A(n_296), .B(n_307), .Y(n_387) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g405 ( .A(n_298), .B(n_363), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_298), .B(n_362), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_299), .B(n_311), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_305), .C(n_315), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_301), .A2(n_336), .B1(n_340), .B2(n_343), .C(n_346), .Y(n_335) );
AOI31xp33_ASAP7_75t_L g430 ( .A1(n_301), .A2(n_431), .A3(n_432), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B1(n_311), .B2(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g431 ( .A(n_311), .Y(n_431) );
INVx1_ASAP7_75t_L g394 ( .A(n_312), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_314), .A2(n_438), .B(n_440), .C(n_442), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_319), .B2(n_323), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_320), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_322), .A2(n_356), .B1(n_375), .B2(n_411), .C(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g406 ( .A(n_323), .Y(n_406) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_326), .B(n_335), .C(n_350), .Y(n_325) );
OAI21xp33_ASAP7_75t_L g376 ( .A1(n_327), .A2(n_377), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_329), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g436 ( .A(n_330), .Y(n_436) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g374 ( .A(n_337), .B(n_357), .Y(n_374) );
INVx1_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g347 ( .A(n_341), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_341), .B(n_379), .Y(n_378) );
NOR4xp25_ASAP7_75t_L g346 ( .A(n_342), .B(n_347), .C(n_348), .D(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_361), .B2(n_362), .C1(n_364), .C2(n_368), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g448 ( .A(n_352), .Y(n_448) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_364), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp5_ASAP7_75t_SL g424 ( .A1(n_369), .A2(n_425), .B(n_427), .Y(n_424) );
NOR4xp25_ASAP7_75t_L g370 ( .A(n_371), .B(n_382), .C(n_395), .D(n_410), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B1(n_374), .B2(n_375), .C(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g451 ( .A(n_372), .Y(n_451) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_379), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OAI222xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_388), .B2(n_389), .C1(n_392), .C2(n_394), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_387), .A2(n_418), .B(n_419), .C(n_430), .Y(n_417) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OAI222xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_401), .B1(n_402), .B2(n_404), .C1(n_406), .C2(n_407), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_412), .A2(n_415), .B1(n_448), .B2(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_445), .B(n_447), .C(n_450), .Y(n_442) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g462 ( .A(n_455), .Y(n_462) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g463 ( .A1(n_461), .A2(n_464), .B(n_777), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_469), .A2(n_474), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx6_ASAP7_75t_L g776 ( .A(n_472), .Y(n_776) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_475), .B(n_731), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_635), .C(n_719), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_578), .C(n_600), .D(n_616), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_516), .B1(n_539), .B2(n_557), .C(n_564), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_496), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_480), .B(n_557), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_480), .B(n_618), .C(n_631), .D(n_633), .Y(n_630) );
INVxp67_ASAP7_75t_L g747 ( .A(n_480), .Y(n_747) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g629 ( .A(n_481), .B(n_567), .Y(n_629) );
AND2x2_ASAP7_75t_L g653 ( .A(n_481), .B(n_496), .Y(n_653) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g620 ( .A(n_482), .B(n_556), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_482), .B(n_641), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_482), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_482), .B(n_497), .Y(n_701) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g555 ( .A(n_483), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g584 ( .A(n_483), .B(n_497), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_483), .B(n_506), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B(n_493), .C(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_494), .A2(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g587 ( .A(n_496), .B(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_496), .A2(n_637), .B1(n_640), .B2(n_642), .C(n_646), .Y(n_636) );
AND2x2_ASAP7_75t_L g695 ( .A(n_496), .B(n_660), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_496), .B(n_677), .Y(n_729) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx3_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
AND2x2_ASAP7_75t_L g604 ( .A(n_497), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g658 ( .A(n_497), .B(n_573), .Y(n_658) );
AND2x2_ASAP7_75t_L g716 ( .A(n_497), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g557 ( .A(n_506), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
INVx1_ASAP7_75t_L g628 ( .A(n_506), .Y(n_628) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_506), .Y(n_634) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_556), .Y(n_679) );
OR2x2_ASAP7_75t_L g718 ( .A(n_506), .B(n_558), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_516), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
AND2x2_ASAP7_75t_L g714 ( .A(n_517), .B(n_711), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_517), .B(n_696), .Y(n_746) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g645 ( .A(n_518), .B(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g694 ( .A(n_518), .B(n_542), .Y(n_694) );
INVx1_ASAP7_75t_L g740 ( .A(n_518), .Y(n_740) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
AND2x2_ASAP7_75t_L g595 ( .A(n_519), .B(n_569), .Y(n_595) );
INVx1_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_519), .B(n_535), .Y(n_618) );
AND2x2_ASAP7_75t_L g686 ( .A(n_524), .B(n_594), .Y(n_686) );
INVx2_ASAP7_75t_L g751 ( .A(n_524), .Y(n_751) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
AND2x2_ASAP7_75t_L g568 ( .A(n_525), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g581 ( .A(n_525), .B(n_543), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_525), .B(n_542), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_525), .Y(n_615) );
INVx1_ASAP7_75t_L g632 ( .A(n_525), .Y(n_632) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_525), .Y(n_644) );
INVx2_ASAP7_75t_L g712 ( .A(n_525), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .Y(n_527) );
INVx2_ASAP7_75t_L g569 ( .A(n_535), .Y(n_569) );
BUFx2_ASAP7_75t_L g666 ( .A(n_535), .Y(n_666) );
AND2x2_ASAP7_75t_L g711 ( .A(n_535), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_541), .B(n_648), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_541), .A2(n_710), .B(n_724), .Y(n_734) );
AND2x2_ASAP7_75t_L g759 ( .A(n_541), .B(n_645), .Y(n_759) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g681 ( .A(n_543), .Y(n_681) );
AND2x2_ASAP7_75t_L g710 ( .A(n_543), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_544), .Y(n_594) );
INVx2_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
OR2x2_ASAP7_75t_L g580 ( .A(n_554), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g648 ( .A(n_554), .B(n_644), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_554), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g749 ( .A(n_554), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_554), .B(n_686), .Y(n_761) );
AND2x2_ASAP7_75t_L g640 ( .A(n_555), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g663 ( .A(n_555), .B(n_557), .Y(n_663) );
INVx2_ASAP7_75t_L g575 ( .A(n_556), .Y(n_575) );
AND2x2_ASAP7_75t_L g603 ( .A(n_556), .B(n_576), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_556), .B(n_628), .Y(n_684) );
AND2x2_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g745 ( .A(n_557), .Y(n_745) );
AND2x2_ASAP7_75t_L g757 ( .A(n_557), .B(n_620), .Y(n_757) );
AND2x2_ASAP7_75t_L g583 ( .A(n_558), .B(n_573), .Y(n_583) );
INVx1_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g576 ( .A(n_563), .B(n_577), .Y(n_576) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_567), .B(n_614), .Y(n_623) );
OR2x2_ASAP7_75t_L g755 ( .A(n_567), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_613), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_568), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g739 ( .A(n_568), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g763 ( .A(n_568), .B(n_610), .Y(n_763) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_569), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g750 ( .A(n_569), .B(n_613), .Y(n_750) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g602 ( .A(n_572), .B(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g764 ( .A(n_572), .Y(n_764) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
AND2x2_ASAP7_75t_L g650 ( .A(n_575), .B(n_583), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_575), .B(n_718), .Y(n_744) );
INVx2_ASAP7_75t_L g589 ( .A(n_576), .Y(n_589) );
INVx3_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
OR2x2_ASAP7_75t_L g669 ( .A(n_576), .B(n_670), .Y(n_669) );
AOI311xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .A3(n_584), .B(n_585), .C(n_596), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_579), .A2(n_617), .B(n_619), .C(n_621), .Y(n_616) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g601 ( .A(n_581), .Y(n_601) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_583), .B(n_599), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_583), .B(n_584), .Y(n_752) );
AND2x2_ASAP7_75t_L g674 ( .A(n_584), .B(n_588), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_590), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g732 ( .A(n_588), .B(n_620), .Y(n_732) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_589), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g626 ( .A(n_589), .Y(n_626) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g617 ( .A(n_593), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g662 ( .A(n_595), .Y(n_662) );
AND2x4_ASAP7_75t_L g724 ( .A(n_595), .B(n_693), .Y(n_724) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_598), .A2(n_664), .B1(n_676), .B2(n_680), .C1(n_682), .C2(n_686), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_604), .C(n_607), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_601), .B(n_645), .Y(n_668) );
INVx1_ASAP7_75t_L g690 ( .A(n_603), .Y(n_690) );
INVx1_ASAP7_75t_L g624 ( .A(n_605), .Y(n_624) );
OR2x2_ASAP7_75t_L g689 ( .A(n_606), .B(n_690), .Y(n_689) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .B(n_614), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_608), .B(n_626), .C(n_627), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_608), .A2(n_645), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_612), .Y(n_665) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_613), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g722 ( .A(n_613), .Y(n_722) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_613), .Y(n_738) );
INVx2_ASAP7_75t_L g696 ( .A(n_614), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_618), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g670 ( .A(n_620), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_629), .C(n_630), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_624), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g758 ( .A(n_624), .Y(n_758) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g639 ( .A(n_631), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_631), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_645), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_631), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g730 ( .A(n_631), .B(n_665), .Y(n_730) );
BUFx3_ASAP7_75t_L g693 ( .A(n_632), .Y(n_693) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND5xp2_ASAP7_75t_L g635 ( .A(n_636), .B(n_654), .C(n_675), .D(n_687), .E(n_702), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI32xp33_ASAP7_75t_L g727 ( .A1(n_639), .A2(n_666), .A3(n_682), .B1(n_728), .B2(n_730), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_641), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g651 ( .A(n_645), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_651), .B2(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_661), .B1(n_663), .B2(n_664), .C(n_667), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g726 ( .A(n_658), .B(n_677), .Y(n_726) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_663), .A2(n_724), .B1(n_742), .B2(n_747), .C(n_748), .Y(n_741) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_L g707 ( .A(n_666), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g685 ( .A(n_677), .Y(n_685) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_698), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_696), .A2(n_743), .B1(n_745), .B2(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_708), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B(n_715), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g756 ( .A(n_711), .Y(n_756) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_725), .C(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_735), .C(n_760), .Y(n_731) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_732), .Y(n_736) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_741), .C(n_753), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B(n_752), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g770 ( .A(n_767), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
endmodule