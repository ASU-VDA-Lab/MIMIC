module real_jpeg_2797_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_32),
.B1(n_35),
.B2(n_77),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_1),
.A2(n_61),
.B1(n_62),
.B2(n_77),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_3),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_32),
.B1(n_35),
.B2(n_124),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_124),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_124),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_85),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_6),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_137)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_54),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_26),
.C(n_28),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_8),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_25),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_8),
.B(n_61),
.C(n_65),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_8),
.B(n_117),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_8),
.B(n_59),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_212),
.Y(n_277)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_11),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_146),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_11),
.A2(n_32),
.B1(n_35),
.B2(n_146),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_146),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_12),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_32),
.B1(n_35),
.B2(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_13),
.A2(n_45),
.B1(n_61),
.B2(n_62),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_15),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_177),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_177),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_177),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_78),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_39),
.B1(n_55),
.B2(n_56),
.Y(n_22)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_25),
.B(n_174),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_27),
.A2(n_28),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_28),
.B(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_32),
.B(n_202),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_32),
.B(n_49),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_35),
.A2(n_43),
.A3(n_48),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_47),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_51)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_43),
.A2(n_75),
.B(n_212),
.C(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_43),
.B(n_212),
.Y(n_213)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_46),
.A2(n_54),
.B1(n_145),
.B2(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_75),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_47),
.A2(n_84),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_47),
.B(n_123),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_47),
.A2(n_121),
.B(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.C(n_74),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_70),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_83),
.C(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_59),
.A2(n_66),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_59),
.A2(n_66),
.B1(n_140),
.B2(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_59),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_69),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_60),
.A2(n_100),
.B1(n_101),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_60),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_60),
.A2(n_219),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_60),
.A2(n_100),
.B1(n_195),
.B2(n_245),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_61),
.B(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_66),
.A2(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_66),
.B(n_198),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_73),
.B1(n_89),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_71),
.A2(n_73),
.B1(n_98),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_71),
.A2(n_73),
.B1(n_185),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_71),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_71),
.A2(n_216),
.B(n_278),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_73),
.A2(n_142),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_73),
.A2(n_173),
.B(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_75),
.A2(n_144),
.B(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_83),
.B1(n_103),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_86),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_153),
.B(n_326),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_149),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_125),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_95),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_95),
.B(n_125),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_95),
.B(n_150),
.Y(n_328)
);

FAx1_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.CI(n_106),
.CON(n_95),
.SN(n_95)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_100),
.A2(n_197),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_113),
.B(n_120),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_108),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_113),
.B1(n_120),
.B2(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_117),
.B(n_118),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_117),
.B1(n_137),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_114),
.A2(n_212),
.B(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_115),
.A2(n_116),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_115),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_115),
.A2(n_116),
.B1(n_192),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_115),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_115),
.A2(n_116),
.B1(n_237),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_116),
.A2(n_191),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_116),
.B(n_206),
.Y(n_239)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_117),
.A2(n_205),
.B(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.C(n_143),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_134),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_135),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_143),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_148),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_149),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_178),
.B(n_325),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_155),
.B(n_158),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_159),
.B(n_162),
.Y(n_323)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_164),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.C(n_175),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_165),
.A2(n_166),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_167),
.B(n_169),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_176),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_320),
.B(n_324),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_289),
.B(n_317),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_231),
.B(n_288),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_207),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_207),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.C(n_199),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_183),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_187),
.C(n_190),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_193),
.B(n_199),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_221),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_208),
.B(n_222),
.C(n_230),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_220),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_209),
.B(n_215),
.C(n_217),
.Y(n_302)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_283),
.B(n_287),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_272),
.B(n_282),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_254),
.B(n_271),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_248),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_248),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B1(n_246),
.B2(n_247),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_243),
.C(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_265),
.B(n_270),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_264),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_263),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_304),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_303),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_303),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_301),
.C(n_302),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_295),
.C(n_299),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_299),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_316),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_310),
.C(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);


endmodule