module fake_jpeg_9794_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_27),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_19),
.C(n_33),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_28),
.C(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_74),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_24),
.B1(n_35),
.B2(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_79),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_44),
.B1(n_48),
.B2(n_19),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_92),
.B1(n_101),
.B2(n_34),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_48),
.B1(n_22),
.B2(n_21),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_91),
.B1(n_34),
.B2(n_20),
.Y(n_138)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_84),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_93),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_0),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_28),
.B(n_22),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_18),
.B1(n_35),
.B2(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_23),
.B1(n_35),
.B2(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_74),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_23),
.B1(n_18),
.B2(n_33),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_21),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_31),
.Y(n_137)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_57),
.B(n_39),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_56),
.C(n_28),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_22),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_101),
.Y(n_144)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_128),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_105),
.C(n_110),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_80),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_54),
.B1(n_66),
.B2(n_69),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_127),
.B1(n_70),
.B2(n_94),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_47),
.A3(n_20),
.B1(n_17),
.B2(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_147),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_95),
.B1(n_97),
.B2(n_87),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_162),
.B1(n_142),
.B2(n_123),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_110),
.C(n_83),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_130),
.C(n_122),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_87),
.B1(n_93),
.B2(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_86),
.B1(n_98),
.B2(n_81),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_112),
.B1(n_84),
.B2(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_168),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_96),
.B(n_75),
.C(n_109),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_40),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_70),
.B1(n_77),
.B2(n_114),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_132),
.B(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_39),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_200),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_135),
.B(n_131),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_181),
.A2(n_185),
.B(n_208),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_117),
.C(n_130),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_177),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_145),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_129),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_190),
.C(n_198),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_129),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_120),
.B1(n_135),
.B2(n_131),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_199),
.B1(n_163),
.B2(n_150),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_132),
.B1(n_121),
.B2(n_141),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_134),
.B1(n_141),
.B2(n_76),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_134),
.C(n_103),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_0),
.C(n_1),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_15),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_17),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_198),
.C(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_212),
.A2(n_237),
.B(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_218),
.C(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_152),
.C(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_221),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_157),
.B(n_167),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_223),
.B(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_152),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_226),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_158),
.B(n_166),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_149),
.B(n_158),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_171),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_228),
.B1(n_191),
.B2(n_184),
.Y(n_239)
);

XNOR2x2_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_161),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_236),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_232),
.B1(n_227),
.B2(n_196),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_154),
.B1(n_76),
.B2(n_20),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_234),
.B1(n_194),
.B2(n_185),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_204),
.B1(n_206),
.B2(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_17),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_209),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_250),
.B1(n_236),
.B2(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_201),
.B1(n_210),
.B2(n_202),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_230),
.B1(n_228),
.B2(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_253),
.C(n_256),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_202),
.B1(n_205),
.B2(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_193),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_220),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_193),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_260),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_225),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_6),
.C(n_12),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_214),
.B(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_239),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_240),
.A2(n_214),
.B(n_218),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_270),
.B(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_265),
.A2(n_269),
.B1(n_15),
.B2(n_3),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_213),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_274),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_247),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_11),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_1),
.B(n_2),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_2),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_281),
.B1(n_269),
.B2(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_256),
.C(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_287),
.C(n_292),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_259),
.C(n_258),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_252),
.B1(n_253),
.B2(n_244),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_276),
.B1(n_271),
.B2(n_262),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_244),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_9),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

OAI221xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.C(n_4),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_263),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_268),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_279),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_282),
.B(n_266),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_266),
.C(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_297),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_280),
.B(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_296),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_287),
.C(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_3),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_302),
.B1(n_306),
.B2(n_307),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_309),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_308),
.B1(n_319),
.B2(n_315),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_318),
.B(n_300),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_326),
.B(n_322),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_303),
.B(n_299),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_327),
.B(n_321),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_323),
.B(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_3),
.C(n_4),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_4),
.Y(n_337)
);


endmodule