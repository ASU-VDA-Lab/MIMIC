module fake_jpeg_30167_n_501 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_501);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_501;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_19),
.A2(n_8),
.B(n_14),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_26),
.C(n_35),
.Y(n_144)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_59),
.B(n_63),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_24),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_8),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_21),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_7),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_9),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_26),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_99),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_57),
.B1(n_77),
.B2(n_61),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_100),
.A2(n_109),
.B1(n_120),
.B2(n_128),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_28),
.B1(n_46),
.B2(n_27),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_127),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_27),
.B1(n_48),
.B2(n_41),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_41),
.B1(n_48),
.B2(n_27),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_114),
.A2(n_124),
.B1(n_126),
.B2(n_132),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_70),
.B1(n_92),
.B2(n_76),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_41),
.B1(n_48),
.B2(n_36),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_51),
.A2(n_46),
.B1(n_47),
.B2(n_40),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_52),
.A2(n_23),
.B1(n_38),
.B2(n_44),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_55),
.A2(n_47),
.B1(n_40),
.B2(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_136),
.A2(n_155),
.B1(n_17),
.B2(n_50),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_53),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_44),
.C(n_43),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_73),
.C(n_96),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_54),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_64),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_82),
.B1(n_69),
.B2(n_87),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_59),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_162),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_159),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_64),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_190),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_168),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_186),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_56),
.B1(n_83),
.B2(n_94),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_167),
.A2(n_173),
.B1(n_195),
.B2(n_150),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_54),
.B(n_81),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_81),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_103),
.B(n_53),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_43),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_102),
.A2(n_97),
.B1(n_89),
.B2(n_93),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_23),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_177),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_125),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_74),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_23),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_183),
.Y(n_228)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_44),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_72),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_191),
.Y(n_245)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_134),
.A2(n_84),
.B1(n_65),
.B2(n_85),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_108),
.B(n_38),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_106),
.A2(n_44),
.B(n_43),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_193),
.A2(n_154),
.B(n_146),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_106),
.B(n_11),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_204),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_111),
.A2(n_43),
.B1(n_38),
.B2(n_91),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_206),
.B1(n_121),
.B2(n_131),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_132),
.A2(n_114),
.B1(n_141),
.B2(n_110),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_182),
.B(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_111),
.B(n_17),
.C(n_50),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_121),
.C(n_141),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_10),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_123),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_205),
.Y(n_242)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g271 ( 
.A1(n_212),
.A2(n_220),
.B(n_163),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_231),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_139),
.B1(n_122),
.B2(n_116),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_217),
.A2(n_226),
.B1(n_233),
.B2(n_234),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_158),
.A2(n_172),
.A3(n_170),
.B1(n_183),
.B2(n_162),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_190),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_191),
.C(n_157),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_227),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_155),
.B1(n_109),
.B2(n_126),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_148),
.C(n_145),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_157),
.A2(n_116),
.B1(n_139),
.B2(n_138),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_160),
.A2(n_138),
.B1(n_123),
.B2(n_133),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_201),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_241),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_160),
.A2(n_130),
.B1(n_150),
.B2(n_50),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_243),
.B1(n_203),
.B2(n_180),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_157),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_1),
.C(n_2),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_186),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_177),
.A2(n_9),
.B(n_13),
.C(n_12),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_176),
.B(n_197),
.C(n_198),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_253),
.A2(n_259),
.B1(n_267),
.B2(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_178),
.B(n_186),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_271),
.B(n_274),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_211),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_261),
.B(n_265),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_264),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_204),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_220),
.A2(n_161),
.B1(n_174),
.B2(n_185),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_211),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_268),
.B(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_214),
.B(n_209),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_273),
.B(n_13),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_159),
.B(n_165),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_240),
.A2(n_161),
.B1(n_174),
.B2(n_206),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_289),
.B1(n_290),
.B2(n_238),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_208),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_209),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_156),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_202),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_281),
.B(n_282),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_208),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_239),
.B(n_205),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_184),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_219),
.A2(n_225),
.B1(n_234),
.B2(n_208),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_287),
.B1(n_238),
.B2(n_232),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_219),
.A2(n_181),
.B1(n_196),
.B2(n_188),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_233),
.A2(n_175),
.B1(n_11),
.B2(n_9),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_226),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_293),
.C(n_305),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_216),
.C(n_227),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_215),
.B1(n_210),
.B2(n_224),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_307),
.B1(n_311),
.B2(n_253),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_259),
.A2(n_231),
.B1(n_218),
.B2(n_244),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_216),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_228),
.B1(n_221),
.B2(n_207),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_228),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_314),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_248),
.C(n_221),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_238),
.B(n_249),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_315),
.A2(n_327),
.B(n_261),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_242),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_320),
.A2(n_266),
.B1(n_283),
.B2(n_264),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_251),
.B(n_250),
.C(n_237),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_276),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_268),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_229),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_279),
.B(n_246),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_328),
.A2(n_335),
.B1(n_319),
.B2(n_322),
.Y(n_382)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_260),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_299),
.C(n_297),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_307),
.A2(n_251),
.B1(n_267),
.B2(n_304),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_336),
.A2(n_347),
.B(n_291),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_303),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_273),
.Y(n_342)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_285),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_322),
.C(n_313),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_353),
.B1(n_310),
.B2(n_308),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_294),
.A2(n_275),
.B1(n_281),
.B2(n_256),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_345),
.A2(n_351),
.B1(n_306),
.B2(n_312),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_287),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_350),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_281),
.B1(n_290),
.B2(n_262),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_354),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_308),
.A2(n_316),
.B1(n_298),
.B2(n_320),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_286),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_255),
.B(n_280),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_357),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_303),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_317),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_360),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_314),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_297),
.B(n_270),
.CI(n_269),
.CON(n_360),
.SN(n_360)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_361),
.A2(n_364),
.B1(n_374),
.B2(n_387),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_291),
.B1(n_299),
.B2(n_327),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_365),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_305),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_372),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_343),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_337),
.A2(n_323),
.B1(n_293),
.B2(n_325),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_380),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_379),
.B1(n_382),
.B2(n_332),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_306),
.B(n_321),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_357),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_345),
.A2(n_312),
.B1(n_309),
.B2(n_319),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_309),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_384),
.C(n_385),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_288),
.C(n_313),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_336),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_337),
.B1(n_338),
.B2(n_330),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_302),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_351),
.C(n_341),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_401),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_380),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_334),
.Y(n_397)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_358),
.Y(n_398)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_386),
.A2(n_330),
.B1(n_329),
.B2(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_360),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_408),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_389),
.B(n_360),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_301),
.C(n_272),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_332),
.C(n_329),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_407),
.C(n_383),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_406),
.A2(n_361),
.B1(n_364),
.B2(n_377),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_347),
.C(n_350),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_373),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_387),
.A2(n_355),
.B1(n_348),
.B2(n_340),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_409),
.A2(n_379),
.B1(n_376),
.B2(n_362),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_373),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_411),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_377),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_339),
.C(n_331),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_413),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_416),
.A2(n_393),
.B1(n_404),
.B2(n_403),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_417),
.A2(n_432),
.B1(n_406),
.B2(n_410),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_415),
.A2(n_378),
.B(n_363),
.Y(n_419)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_424),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_413),
.A2(n_384),
.B(n_374),
.Y(n_422)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_411),
.A2(n_390),
.B(n_385),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_395),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_407),
.B(n_375),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_394),
.C(n_396),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_397),
.A2(n_381),
.B(n_331),
.Y(n_430)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_409),
.A2(n_301),
.B(n_257),
.C(n_321),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_302),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_408),
.Y(n_448)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_446),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_439),
.A2(n_416),
.B1(n_393),
.B2(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_392),
.C(n_405),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_444),
.C(n_426),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_398),
.Y(n_441)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_394),
.C(n_396),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_451),
.Y(n_460)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_428),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_414),
.B1(n_432),
.B2(n_257),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_450),
.A2(n_417),
.B1(n_423),
.B2(n_433),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_427),
.B(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_434),
.B(n_399),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_453),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_464),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_419),
.B(n_425),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_456),
.Y(n_470)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_445),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_462),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_442),
.A2(n_430),
.B(n_418),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_458),
.B(n_461),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_450),
.A2(n_447),
.B1(n_445),
.B2(n_443),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_439),
.A2(n_432),
.B1(n_401),
.B2(n_402),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_466),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_429),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_432),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_437),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_472),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_438),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g473 ( 
.A(n_463),
.B(n_438),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_473),
.A2(n_453),
.B(n_446),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_460),
.A2(n_444),
.B(n_440),
.Y(n_474)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_477),
.A2(n_457),
.B1(n_458),
.B2(n_454),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_462),
.C(n_464),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_469),
.C(n_471),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_468),
.B(n_466),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_483),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_455),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_476),
.B(n_459),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_485),
.A2(n_486),
.B(n_487),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_424),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_258),
.C(n_246),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_486),
.A2(n_478),
.B(n_475),
.C(n_479),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_487),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_483),
.C(n_484),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_495),
.B(n_496),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_493),
.B(n_481),
.Y(n_495)
);

NAND4xp25_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_491),
.C(n_490),
.D(n_489),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_498),
.B(n_497),
.Y(n_499)
);

AOI31xp33_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_480),
.A3(n_229),
.B(n_237),
.Y(n_500)
);

OAI321xp33_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_237),
.A3(n_12),
.B1(n_5),
.B2(n_4),
.C(n_1),
.Y(n_501)
);


endmodule