module fake_jpeg_9567_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_14),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_53),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_17),
.B1(n_19),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_40),
.B1(n_32),
.B2(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_27),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_27),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_15),
.C(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_29),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_31),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_31),
.A2(n_24),
.B1(n_29),
.B2(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_43),
.B1(n_62),
.B2(n_27),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_16),
.B(n_30),
.C(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_51),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_37),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_58),
.Y(n_88)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_77),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_0),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_53),
.B(n_67),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_45),
.CI(n_54),
.CON(n_87),
.SN(n_87)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_56),
.B1(n_55),
.B2(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_100),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_74),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_70),
.B1(n_83),
.B2(n_72),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_48),
.A3(n_46),
.B1(n_44),
.B2(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_101),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_56),
.B1(n_43),
.B2(n_44),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_104),
.B1(n_77),
.B2(n_64),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_23),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_78),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_116),
.B(n_92),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_124),
.B1(n_89),
.B2(n_103),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_65),
.B1(n_72),
.B2(n_79),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_115),
.B(n_117),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_95),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_74),
.B1(n_59),
.B2(n_23),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_75),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_88),
.C(n_91),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_78),
.B1(n_59),
.B2(n_81),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_86),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_150),
.C(n_37),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_144),
.B(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_137),
.B1(n_38),
.B2(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_103),
.B1(n_93),
.B2(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_100),
.B1(n_97),
.B2(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_113),
.B1(n_112),
.B2(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_94),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_94),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_87),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_119),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_100),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_149),
.A3(n_129),
.B1(n_138),
.B2(n_135),
.C1(n_137),
.C2(n_145),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_87),
.C(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_169),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_88),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_163),
.C(n_164),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_41),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_116),
.B1(n_117),
.B2(n_115),
.C(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NOR4xp25_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_115),
.C(n_97),
.D(n_104),
.Y(n_157)
);

OA21x2_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_156),
.B(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_81),
.B1(n_73),
.B2(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_99),
.B1(n_28),
.B2(n_38),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_166),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_125),
.C(n_37),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_170),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_37),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_41),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_130),
.B1(n_133),
.B2(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_129),
.A3(n_148),
.B1(n_146),
.B2(n_150),
.C1(n_137),
.C2(n_135),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_178),
.B(n_99),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_129),
.A3(n_150),
.B1(n_139),
.B2(n_132),
.C1(n_131),
.C2(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_164),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_183),
.B(n_23),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_161),
.B1(n_158),
.B2(n_155),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_23),
.B1(n_99),
.B2(n_41),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_184),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_8),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_41),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_159),
.C(n_162),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_191),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_185),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_200),
.C(n_205),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

AOI321xp33_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_155),
.A3(n_162),
.B1(n_163),
.B2(n_154),
.C(n_171),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_206),
.B(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_160),
.B1(n_99),
.B2(n_2),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_180),
.B1(n_196),
.B2(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_41),
.C(n_23),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_183),
.C(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_198),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_174),
.B(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_178),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_214),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_186),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_190),
.C(n_1),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_12),
.C(n_11),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_227),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_221),
.B1(n_220),
.B2(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_207),
.B1(n_202),
.B2(n_208),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_230),
.B1(n_215),
.B2(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_13),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_232),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_242),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_210),
.C(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_0),
.C(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_237),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_212),
.A3(n_210),
.B1(n_12),
.B2(n_10),
.C(n_9),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_242),
.B1(n_4),
.B2(n_5),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_0),
.C(n_3),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_232),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_235),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_247),
.C(n_4),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_4),
.B(n_6),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_256),
.C(n_7),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_7),
.B1(n_237),
.B2(n_223),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_255),
.Y(n_258)
);


endmodule