module fake_jpeg_28291_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_3),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_22),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_16),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_32),
.B1(n_23),
.B2(n_19),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_60),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_20),
.B(n_23),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_61),
.C(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_15),
.B(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_44),
.B1(n_49),
.B2(n_41),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_74),
.B1(n_38),
.B2(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_41),
.C(n_43),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_52),
.C(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_41),
.B1(n_38),
.B2(n_21),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_83),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_74),
.B1(n_69),
.B2(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_69),
.B(n_41),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_90),
.B(n_81),
.C(n_75),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_87),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

AO221x1_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_68),
.B1(n_62),
.B2(n_80),
.C(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_89),
.C(n_84),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_84),
.A3(n_85),
.B1(n_21),
.B2(n_11),
.C(n_12),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_94),
.B1(n_91),
.B2(n_12),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);


endmodule