module real_aes_16874_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_0), .A2(n_50), .B1(n_566), .B2(n_570), .Y(n_565) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_0), .Y(n_629) );
INVx1_ASAP7_75t_L g594 ( .A(n_1), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_1), .B(n_551), .Y(n_602) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g508 ( .A(n_3), .Y(n_508) );
INVx1_ASAP7_75t_L g514 ( .A(n_4), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_4), .A2(n_14), .B1(n_613), .B2(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_5), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g499 ( .A(n_6), .Y(n_499) );
INVx1_ASAP7_75t_L g505 ( .A(n_6), .Y(n_505) );
INVx1_ASAP7_75t_L g704 ( .A(n_7), .Y(n_704) );
INVx2_ASAP7_75t_L g489 ( .A(n_8), .Y(n_489) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_9), .A2(n_29), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g538 ( .A(n_10), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_11), .B(n_201), .Y(n_200) );
XNOR2xp5_ASAP7_75t_L g477 ( .A(n_12), .B(n_478), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_13), .Y(n_225) );
INVx1_ASAP7_75t_L g525 ( .A(n_14), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_15), .B(n_91), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_16), .B(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_17), .Y(n_153) );
INVx1_ASAP7_75t_L g693 ( .A(n_18), .Y(n_693) );
INVx1_ASAP7_75t_L g500 ( .A(n_19), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_20), .Y(n_229) );
INVx1_ASAP7_75t_L g491 ( .A(n_21), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_21), .A2(n_59), .B1(n_611), .B2(n_613), .Y(n_610) );
INVx2_ASAP7_75t_L g488 ( .A(n_22), .Y(n_488) );
INVx1_ASAP7_75t_L g533 ( .A(n_22), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_23), .B(n_126), .Y(n_171) );
INVx2_ASAP7_75t_L g677 ( .A(n_24), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_25), .B(n_87), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_26), .B(n_143), .Y(n_203) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_27), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_27), .A2(n_50), .B1(n_634), .B2(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g541 ( .A(n_28), .Y(n_541) );
AND2x2_ASAP7_75t_L g231 ( .A(n_30), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_31), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_32), .B(n_91), .Y(n_257) );
INVx1_ASAP7_75t_L g699 ( .A(n_32), .Y(n_699) );
BUFx2_ASAP7_75t_L g705 ( .A(n_33), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_34), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g720 ( .A(n_34), .Y(n_720) );
BUFx3_ASAP7_75t_L g497 ( .A(n_35), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_36), .B(n_261), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_37), .A2(n_116), .B(n_124), .C(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g83 ( .A(n_38), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_38), .Y(n_663) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_40), .A2(n_42), .B1(n_175), .B2(n_185), .Y(n_184) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_41), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_43), .B(n_106), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_44), .B(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_45), .Y(n_230) );
INVx1_ASAP7_75t_L g522 ( .A(n_46), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_47), .B(n_175), .Y(n_174) );
BUFx3_ASAP7_75t_L g701 ( .A(n_48), .Y(n_701) );
INVx1_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_51), .Y(n_190) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_52), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_53), .B(n_106), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_54), .B(n_113), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_55), .B(n_87), .C(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g577 ( .A(n_56), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_57), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g535 ( .A(n_59), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_60), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_61), .B(n_126), .Y(n_158) );
INVx1_ASAP7_75t_L g713 ( .A(n_61), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_62), .B(n_120), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_63), .A2(n_71), .B1(n_91), .B2(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g689 ( .A(n_63), .Y(n_689) );
BUFx3_ASAP7_75t_L g551 ( .A(n_64), .Y(n_551) );
INVx1_ASAP7_75t_L g555 ( .A(n_64), .Y(n_555) );
INVx1_ASAP7_75t_L g583 ( .A(n_65), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_66), .B(n_126), .Y(n_156) );
NAND2xp33_ASAP7_75t_SL g141 ( .A(n_67), .B(n_115), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_68), .B(n_155), .Y(n_170) );
INVx1_ASAP7_75t_L g486 ( .A(n_69), .Y(n_486) );
INVx1_ASAP7_75t_L g532 ( .A(n_69), .Y(n_532) );
INVx2_ASAP7_75t_L g601 ( .A(n_69), .Y(n_601) );
INVx1_ASAP7_75t_L g552 ( .A(n_70), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g114 ( .A(n_72), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_73), .B(n_143), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g137 ( .A(n_74), .B(n_115), .C(n_136), .Y(n_137) );
INVx1_ASAP7_75t_SL g690 ( .A(n_75), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_76), .B(n_113), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_77), .B(n_91), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_94), .B(n_476), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
AND2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_85), .Y(n_81) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_82), .A2(n_180), .A3(n_188), .B(n_189), .Y(n_179) );
INVx2_ASAP7_75t_L g221 ( .A(n_82), .Y(n_221) );
BUFx10_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx10_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_84), .Y(n_665) );
INVxp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g723 ( .A1(n_86), .A2(n_664), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_89), .Y(n_86) );
O2A1O1Ixp5_ASAP7_75t_L g152 ( .A1(n_87), .A2(n_153), .B(n_154), .C(n_156), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_87), .A2(n_173), .B(n_174), .Y(n_172) );
INVx6_ASAP7_75t_L g183 ( .A(n_87), .Y(n_183) );
BUFx8_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g117 ( .A(n_88), .Y(n_117) );
INVx2_ASAP7_75t_L g122 ( .A(n_88), .Y(n_122) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx3_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
INVx1_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_93), .Y(n_175) );
INVx1_ASAP7_75t_L g185 ( .A(n_93), .Y(n_185) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_93), .Y(n_197) );
INVx2_ASAP7_75t_L g226 ( .A(n_93), .Y(n_226) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_96), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_408), .Y(n_96) );
NAND4xp25_ASAP7_75t_L g97 ( .A(n_98), .B(n_283), .C(n_323), .D(n_372), .Y(n_97) );
NOR2xp67_ASAP7_75t_L g98 ( .A(n_99), .B(n_232), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_146), .B1(n_204), .B2(n_213), .Y(n_99) );
INVx1_ASAP7_75t_L g404 ( .A(n_100), .Y(n_404) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_101), .B(n_251), .Y(n_320) );
AND2x2_ASAP7_75t_L g351 ( .A(n_101), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_129), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_102), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g275 ( .A(n_102), .Y(n_275) );
AND2x2_ASAP7_75t_L g450 ( .A(n_102), .B(n_318), .Y(n_450) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g215 ( .A(n_103), .Y(n_215) );
AND2x2_ASAP7_75t_L g303 ( .A(n_103), .B(n_265), .Y(n_303) );
AND2x2_ASAP7_75t_L g347 ( .A(n_103), .B(n_252), .Y(n_347) );
OR2x2_ASAP7_75t_L g365 ( .A(n_103), .B(n_366), .Y(n_365) );
INVx4_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g269 ( .A(n_104), .B(n_252), .Y(n_269) );
BUFx2_ASAP7_75t_L g326 ( .A(n_104), .Y(n_326) );
OR2x2_ASAP7_75t_L g334 ( .A(n_104), .B(n_292), .Y(n_334) );
INVx1_ASAP7_75t_L g389 ( .A(n_104), .Y(n_389) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_110), .Y(n_104) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_SL g127 ( .A(n_107), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g132 ( .A(n_107), .Y(n_132) );
INVx2_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_118), .B(n_127), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_114), .B(n_116), .Y(n_111) );
OAI22xp33_ASAP7_75t_L g228 ( .A1(n_113), .A2(n_175), .B1(n_229), .B2(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_116), .A2(n_139), .B(n_141), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_116), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_116), .A2(n_256), .B(n_257), .Y(n_255) );
BUFx4f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_121), .B1(n_123), .B2(n_125), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_120), .A2(n_158), .B(n_159), .Y(n_157) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g187 ( .A(n_122), .Y(n_187) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_126), .A2(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_128), .A2(n_134), .B(n_138), .Y(n_133) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_128), .A2(n_152), .B(n_157), .Y(n_151) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_128), .A2(n_169), .B(n_172), .Y(n_168) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_128), .A2(n_194), .B(n_198), .Y(n_193) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_128), .A2(n_255), .B(n_258), .Y(n_254) );
AND2x2_ASAP7_75t_L g216 ( .A(n_129), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g328 ( .A(n_129), .B(n_305), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_129), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g366 ( .A(n_130), .Y(n_366) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_130), .Y(n_371) );
AND2x2_ASAP7_75t_L g388 ( .A(n_130), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g278 ( .A(n_131), .B(n_218), .Y(n_278) );
INVx1_ASAP7_75t_L g292 ( .A(n_131), .Y(n_292) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_142), .Y(n_131) );
INVx1_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
NAND2x1_ASAP7_75t_L g146 ( .A(n_147), .B(n_162), .Y(n_146) );
AND2x4_ASAP7_75t_L g453 ( .A(n_147), .B(n_381), .Y(n_453) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
INVxp67_ASAP7_75t_SL g212 ( .A(n_148), .Y(n_212) );
BUFx3_ASAP7_75t_L g247 ( .A(n_148), .Y(n_247) );
INVx1_ASAP7_75t_L g313 ( .A(n_148), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_148), .B(n_165), .Y(n_316) );
AND2x2_ASAP7_75t_L g341 ( .A(n_148), .B(n_192), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_148), .Y(n_344) );
AND2x2_ASAP7_75t_L g376 ( .A(n_148), .B(n_241), .Y(n_376) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_161), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_150), .A2(n_151), .B(n_161), .Y(n_242) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_150), .A2(n_254), .B(n_263), .Y(n_253) );
OAI21xp33_ASAP7_75t_SL g281 ( .A1(n_150), .A2(n_254), .B(n_263), .Y(n_281) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_177), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g285 ( .A(n_164), .B(n_271), .Y(n_285) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g311 ( .A(n_166), .B(n_298), .Y(n_311) );
AND2x2_ASAP7_75t_L g340 ( .A(n_166), .B(n_179), .Y(n_340) );
OR2x2_ASAP7_75t_L g436 ( .A(n_166), .B(n_179), .Y(n_436) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_176), .Y(n_166) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_167), .A2(n_193), .B(n_203), .Y(n_192) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_167), .A2(n_168), .B(n_176), .Y(n_210) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_167), .A2(n_193), .B(n_203), .Y(n_241) );
INVx2_ASAP7_75t_L g182 ( .A(n_175), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_175), .A2(n_195), .B(n_196), .Y(n_194) );
AND2x2_ASAP7_75t_L g315 ( .A(n_177), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g464 ( .A(n_177), .Y(n_464) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
OR2x2_ASAP7_75t_L g398 ( .A(n_178), .B(n_208), .Y(n_398) );
INVx1_ASAP7_75t_L g420 ( .A(n_178), .Y(n_420) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_192), .Y(n_178) );
AND2x2_ASAP7_75t_L g236 ( .A(n_179), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g271 ( .A(n_179), .B(n_241), .Y(n_271) );
INVx1_ASAP7_75t_L g298 ( .A(n_179), .Y(n_298) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_179), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_179), .B(n_192), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B1(n_184), .B2(n_186), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_186), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
INVx2_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
AND2x2_ASAP7_75t_L g322 ( .A(n_192), .B(n_242), .Y(n_322) );
INVx2_ASAP7_75t_L g261 ( .A(n_197), .Y(n_261) );
AOI21x1_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR3x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .C(n_211), .Y(n_205) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_208), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g321 ( .A(n_208), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g361 ( .A(n_208), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_208), .B(n_384), .Y(n_416) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_209), .B(n_297), .Y(n_357) );
AND2x2_ASAP7_75t_L g381 ( .A(n_209), .B(n_241), .Y(n_381) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g392 ( .A(n_212), .B(n_271), .Y(n_392) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_215), .B(n_278), .Y(n_457) );
AND2x4_ASAP7_75t_L g449 ( .A(n_216), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_216), .B(n_269), .Y(n_463) );
INVx2_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
INVx1_ASAP7_75t_L g268 ( .A(n_217), .Y(n_268) );
INVx2_ASAP7_75t_L g353 ( .A(n_217), .Y(n_353) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g337 ( .A(n_218), .Y(n_337) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B(n_231), .Y(n_218) );
NOR2xp67_ASAP7_75t_SL g219 ( .A(n_220), .B(n_221), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_272), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_248), .B1(n_266), .B2(n_270), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_238), .B(n_243), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g300 ( .A(n_236), .B(n_247), .Y(n_300) );
AND2x2_ASAP7_75t_L g460 ( .A(n_236), .B(n_341), .Y(n_460) );
BUFx2_ASAP7_75t_L g331 ( .A(n_237), .Y(n_331) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g330 ( .A(n_240), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g245 ( .A(n_241), .Y(n_245) );
INVx1_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
INVx1_ASAP7_75t_L g422 ( .A(n_242), .Y(n_422) );
AOI31xp33_ASAP7_75t_L g440 ( .A1(n_243), .A2(n_441), .A3(n_442), .B(n_443), .Y(n_440) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_244), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_245), .B(n_340), .Y(n_439) );
INVx2_ASAP7_75t_L g467 ( .A(n_245), .Y(n_467) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_246), .Y(n_282) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g295 ( .A(n_247), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_247), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g425 ( .A(n_247), .B(n_385), .Y(n_425) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_264), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g336 ( .A(n_252), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g305 ( .A(n_253), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_262), .Y(n_258) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
INVx1_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
INVx1_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
AND2x2_ASAP7_75t_L g370 ( .A(n_269), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g426 ( .A(n_269), .B(n_353), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_270), .A2(n_343), .B(n_345), .Y(n_342) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_282), .Y(n_272) );
NAND3x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .C(n_279), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g444 ( .A(n_275), .B(n_364), .Y(n_444) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2x1_ASAP7_75t_SL g397 ( .A(n_277), .B(n_309), .Y(n_397) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g317 ( .A(n_278), .B(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_279), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_279), .B(n_388), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_279), .B(n_388), .Y(n_461) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g364 ( .A(n_281), .B(n_337), .Y(n_364) );
AND2x2_ASAP7_75t_L g284 ( .A(n_282), .B(n_285), .Y(n_284) );
AOI221x1_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_286), .B1(n_293), .B2(n_302), .C(n_306), .Y(n_283) );
AOI32xp33_ASAP7_75t_L g465 ( .A1(n_285), .A2(n_466), .A3(n_471), .B1(n_472), .B2(n_474), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_290), .B(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_292), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_292), .Y(n_308) );
OR2x2_ASAP7_75t_L g421 ( .A(n_292), .B(n_422), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .C(n_301), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g343 ( .A(n_296), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g360 ( .A(n_296), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_299), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_395) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g473 ( .A(n_303), .Y(n_473) );
INVx2_ASAP7_75t_L g318 ( .A(n_305), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B(n_314), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g442 ( .A(n_311), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_312), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_319), .B2(n_321), .Y(n_314) );
AND2x4_ASAP7_75t_L g411 ( .A(n_317), .B(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g470 ( .A(n_318), .Y(n_470) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g349 ( .A(n_322), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_322), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_322), .B(n_350), .Y(n_441) );
AOI211x1_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B(n_332), .C(n_358), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR3x2_ASAP7_75t_L g433 ( .A(n_326), .B(n_328), .C(n_329), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_327), .A2(n_349), .B1(n_351), .B2(n_354), .Y(n_348) );
NOR2x1p5_ASAP7_75t_SL g327 ( .A(n_328), .B(n_329), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_328), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g350 ( .A(n_331), .Y(n_350) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_338), .B(n_342), .C(n_348), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_340), .B(n_344), .Y(n_355) );
INVx1_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_340), .B(n_447), .Y(n_455) );
OAI32xp33_ASAP7_75t_L g430 ( .A1(n_341), .A2(n_386), .A3(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g447 ( .A(n_341), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_341), .B(n_361), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_344), .B(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g391 ( .A(n_350), .B(n_376), .Y(n_391) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g400 ( .A(n_353), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_356), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_367), .B2(n_369), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g387 ( .A(n_364), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_364), .B(n_371), .Y(n_475) );
INVx1_ASAP7_75t_SL g401 ( .A(n_365), .Y(n_401) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_395), .C(n_402), .Y(n_372) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_386), .B(n_390), .Y(n_373) );
NOR2xp33_ASAP7_75t_SL g374 ( .A(n_375), .B(n_379), .Y(n_374) );
INVxp67_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .C(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_388), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g403 ( .A(n_391), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_396), .A2(n_447), .B1(n_448), .B2(n_451), .C(n_452), .Y(n_446) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI32xp33_ASAP7_75t_L g402 ( .A1(n_399), .A2(n_403), .A3(n_404), .B1(n_405), .B2(n_407), .Y(n_402) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_405), .A2(n_415), .B1(n_416), .B2(n_417), .C(n_423), .Y(n_414) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_427), .C(n_445), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_414), .Y(n_409) );
AOI211x1_ASAP7_75t_L g427 ( .A1(n_410), .A2(n_428), .B(n_430), .C(n_437), .Y(n_427) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR2x1_ASAP7_75t_SL g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g429 ( .A(n_420), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AO21x1_ASAP7_75t_L g437 ( .A1(n_426), .A2(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g471 ( .A(n_442), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_458), .Y(n_445) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI21xp33_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_462), .Y(n_459) );
NOR2xp67_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g468 ( .A(n_467), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_661), .B2(n_666), .C(n_714), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_478), .A2(n_715), .B1(n_719), .B2(n_721), .Y(n_714) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_539), .C(n_597), .D(n_627), .Y(n_479) );
OAI33xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_490), .A3(n_507), .B1(n_519), .B2(n_526), .B3(n_534), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx4f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g620 ( .A(n_484), .Y(n_620) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_484), .Y(n_660) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g596 ( .A(n_485), .Y(n_596) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g682 ( .A(n_487), .Y(n_682) );
NAND2xp33_ASAP7_75t_SL g487 ( .A(n_488), .B(n_489), .Y(n_487) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_488), .Y(n_658) );
INVx1_ASAP7_75t_L g676 ( .A(n_488), .Y(n_676) );
INVx3_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
BUFx3_ASAP7_75t_L g637 ( .A(n_489), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B1(n_500), .B2(n_501), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_494), .A2(n_535), .B1(n_536), .B2(n_538), .Y(n_534) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x4_ASAP7_75t_L g645 ( .A(n_496), .B(n_530), .Y(n_645) );
OR2x4_ASAP7_75t_L g651 ( .A(n_496), .B(n_647), .Y(n_651) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_497), .Y(n_506) );
INVx2_ASAP7_75t_L g513 ( .A(n_497), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_497), .B(n_505), .Y(n_518) );
AND2x4_ASAP7_75t_L g631 ( .A(n_497), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g512 ( .A(n_499), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_500), .A2(n_538), .B1(n_607), .B2(n_622), .C(n_625), .Y(n_621) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g537 ( .A(n_503), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
BUFx2_ASAP7_75t_L g641 ( .A(n_504), .Y(n_641) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g632 ( .A(n_505), .Y(n_632) );
BUFx2_ASAP7_75t_L g638 ( .A(n_506), .Y(n_638) );
INVx2_ASAP7_75t_L g674 ( .A(n_506), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_514), .B2(n_515), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_508), .A2(n_522), .B1(n_604), .B2(n_607), .C(n_610), .Y(n_603) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx8_ASAP7_75t_L g521 ( .A(n_511), .Y(n_521) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_511), .Y(n_648) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g524 ( .A(n_517), .Y(n_524) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g654 ( .A(n_518), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_523), .B2(n_525), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND3x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .C(n_533), .Y(n_529) );
AND2x4_ASAP7_75t_L g642 ( .A(n_530), .B(n_631), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_530), .Y(n_647) );
OR2x6_ASAP7_75t_L g653 ( .A(n_530), .B(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_L g675 ( .A(n_530), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI31xp33_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_558), .A3(n_576), .B(n_591), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_552), .B2(n_553), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_541), .A2(n_552), .B1(n_644), .B2(n_646), .Y(n_643) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g556 ( .A(n_547), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g563 ( .A(n_547), .B(n_548), .Y(n_563) );
INVx1_ASAP7_75t_L g573 ( .A(n_547), .Y(n_573) );
INVx2_ASAP7_75t_L g581 ( .A(n_547), .Y(n_581) );
INVx2_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
NAND2x1_ASAP7_75t_L g609 ( .A(n_547), .B(n_548), .Y(n_609) );
INVx2_ASAP7_75t_L g557 ( .A(n_548), .Y(n_557) );
BUFx2_ASAP7_75t_L g569 ( .A(n_548), .Y(n_569) );
INVx1_ASAP7_75t_L g582 ( .A(n_548), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_548), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g606 ( .A(n_548), .B(n_581), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_548), .B(n_590), .Y(n_615) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g575 ( .A(n_550), .Y(n_575) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g568 ( .A(n_551), .Y(n_568) );
AND2x4_ASAP7_75t_L g571 ( .A(n_551), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g618 ( .A(n_551), .B(n_594), .Y(n_618) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B(n_565), .C(n_574), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g574 ( .A(n_562), .B(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g578 ( .A(n_568), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g587 ( .A(n_568), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_583), .B2(n_584), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_577), .A2(n_583), .B1(n_650), .B2(n_652), .Y(n_649) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_579), .Y(n_626) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g612 ( .A(n_580), .Y(n_612) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_603), .B1(n_616), .B2(n_621), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx3_ASAP7_75t_L g624 ( .A(n_606), .Y(n_624) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI31xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_643), .A3(n_649), .B(n_655), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_633), .C(n_642), .Y(n_628) );
BUFx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
AND2x4_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
CKINVDCx14_ASAP7_75t_R g655 ( .A(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g684 ( .A(n_663), .Y(n_684) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_665), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g724 ( .A(n_665), .B(n_684), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_685), .B1(n_708), .B2(n_712), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx12f_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g716 ( .A(n_669), .Y(n_716) );
BUFx8_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_677), .B(n_678), .C(n_683), .Y(n_670) );
AND2x2_ASAP7_75t_L g711 ( .A(n_671), .B(n_678), .Y(n_711) );
INVx4_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x6_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_673), .B(n_679), .C(n_682), .Y(n_678) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g681 ( .A(n_677), .Y(n_681) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g710 ( .A(n_683), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_685), .A2(n_712), .B1(n_716), .B2(n_717), .Y(n_715) );
XNOR2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_695), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_693), .B2(n_694), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_689), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_690), .Y(n_692) );
CKINVDCx14_ASAP7_75t_R g694 ( .A(n_693), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_702), .B2(n_703), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_704), .Y(n_707) );
INVx1_ASAP7_75t_L g706 ( .A(n_705), .Y(n_706) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g718 ( .A(n_709), .Y(n_718) );
OR2x6_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
endmodule