module real_jpeg_9998_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_26),
.B1(n_29),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_52),
.B1(n_61),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_8),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_101),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_26),
.B1(n_29),
.B2(n_101),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_101),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_9),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_54),
.B(n_58),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_9),
.A2(n_52),
.B1(n_61),
.B2(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_65),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_37),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_37),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_81),
.B1(n_82),
.B2(n_225),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_62),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_12),
.A2(n_34),
.B1(n_52),
.B2(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_52),
.B1(n_61),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_13),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_145),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_145),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_14),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_40),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_15),
.A2(n_28),
.B1(n_57),
.B2(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_15),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_15),
.A2(n_28),
.B1(n_52),
.B2(n_61),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_19),
.B(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.C(n_89),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_20),
.A2(n_21),
.B1(n_78),
.B2(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_49),
.C(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_24),
.A2(n_82),
.B(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_26),
.A2(n_29),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_26),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_29),
.B(n_45),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_29),
.B(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_30),
.A2(n_31),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_32),
.A2(n_81),
.B(n_209),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_36),
.A2(n_44),
.B(n_95),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_38),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_37),
.B(n_69),
.Y(n_253)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_38),
.A2(n_74),
.B1(n_248),
.B2(n_253),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_46),
.B(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_41),
.A2(n_44),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_41),
.A2(n_44),
.B1(n_215),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_41),
.A2(n_44),
.B1(n_238),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_41),
.A2(n_121),
.B(n_246),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_43),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_44),
.B(n_149),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_66),
.B2(n_77),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_60),
.B(n_63),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_56),
.B1(n_60),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_51),
.A2(n_56),
.B1(n_100),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_51),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_52),
.A2(n_53),
.B(n_149),
.C(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.C(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_69),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_58),
.B(n_149),
.CON(n_248),
.SN(n_248)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_65),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_72),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_67),
.A2(n_139),
.B1(n_140),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_67),
.A2(n_139),
.B1(n_170),
.B2(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_67),
.B(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_73),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_68),
.B(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_68),
.A2(n_73),
.B1(n_193),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_73),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_78),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_88),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_80),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_84),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_81),
.A2(n_82),
.B1(n_207),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_81),
.A2(n_83),
.B(n_93),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_82),
.B(n_149),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_86),
.A2(n_97),
.B(n_123),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_94),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_105),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_116),
.CI(n_125),
.CON(n_105),
.SN(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B(n_124),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_156),
.B(n_279),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_153),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_130),
.B(n_153),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_135),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_134),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_136),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.C(n_146),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_198),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_179),
.B(n_197),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_199),
.C(n_278),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_176),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_169),
.B1(n_175),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_180),
.B(n_182),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_276),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_186),
.Y(n_276)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_191),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_194),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_272),
.B(n_277),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_257),
.B(n_271),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_241),
.B(n_256),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_232),
.B(n_240),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_221),
.B(n_231),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_210),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_220),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_220),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_242),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.CI(n_239),
.CON(n_235),
.SN(n_235)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_255),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_250),
.C(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_251),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_254),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_266),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_268),
.C(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);


endmodule