module fake_jpeg_23787_n_35 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2x1_ASAP7_75t_SL g18 ( 
.A(n_4),
.B(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_10),
.B(n_13),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.C(n_18),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_17),
.B1(n_18),
.B2(n_15),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_31),
.Y(n_33)
);

AOI221xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_29),
.B1(n_1),
.B2(n_5),
.C(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);


endmodule