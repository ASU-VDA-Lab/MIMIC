module real_jpeg_18096_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_290;
wire n_239;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_0),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_0),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_0),
.A2(n_254),
.B1(n_291),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_0),
.A2(n_291),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_0),
.A2(n_291),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_1),
.A2(n_153),
.B1(n_223),
.B2(n_228),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_1),
.A2(n_153),
.B1(n_278),
.B2(n_282),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_2),
.A2(n_101),
.B1(n_254),
.B2(n_257),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_2),
.A2(n_101),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_2),
.A2(n_101),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_4),
.A2(n_93),
.B1(n_328),
.B2(n_332),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_4),
.A2(n_93),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_4),
.A2(n_93),
.B1(n_321),
.B2(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_5),
.Y(n_405)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_5),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_158),
.B1(n_162),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_6),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_6),
.A2(n_164),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_6),
.A2(n_164),
.B1(n_534),
.B2(n_539),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_7),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_7),
.A2(n_177),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_9),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_11),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_11),
.A2(n_212),
.B1(n_328),
.B2(n_338),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_67),
.B1(n_137),
.B2(n_142),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_13),
.A2(n_67),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_13),
.A2(n_67),
.B1(n_553),
.B2(n_555),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_14),
.B(n_272),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g299 ( 
.A1(n_14),
.A2(n_300),
.A3(n_301),
.B1(n_304),
.B2(n_306),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_14),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_14),
.A2(n_305),
.B1(n_348),
.B2(n_351),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_14),
.B(n_260),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_14),
.A2(n_165),
.B1(n_466),
.B2(n_472),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_14),
.A2(n_271),
.B(n_499),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_16),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_16),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_17),
.A2(n_31),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_17),
.A2(n_31),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_17),
.A2(n_31),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_523),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_292),
.B(n_520),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_246),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_22),
.B(n_246),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_181),
.Y(n_22)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_23),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_69),
.C(n_106),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_24),
.B(n_69),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_26),
.A2(n_38),
.B1(n_253),
.B2(n_260),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_29),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_30),
.Y(n_227)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_37),
.A2(n_62),
.B1(n_63),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_37),
.A2(n_62),
.B1(n_347),
.B2(n_356),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_37),
.A2(n_62),
.B1(n_356),
.B2(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_37),
.A2(n_62),
.B1(n_364),
.B2(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_38),
.A2(n_260),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_46),
.B(n_54),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_43),
.Y(n_350)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_45),
.Y(n_230)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_45),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_45),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_46),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_52),
.Y(n_269)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_53),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_53),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_60),
.Y(n_383)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_62),
.Y(n_260)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_66),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_89),
.B1(n_97),
.B2(n_105),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_70),
.A2(n_97),
.B1(n_105),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_70),
.A2(n_89),
.B1(n_105),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_70),
.A2(n_105),
.B1(n_288),
.B2(n_498),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_70),
.A2(n_105),
.B1(n_217),
.B2(n_552),
.Y(n_551)
);

AO21x2_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_77),
.B(n_84),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_73),
.Y(n_265)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_77),
.A2(n_263),
.B1(n_270),
.B2(n_274),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_79),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_92),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_92),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_92),
.Y(n_501)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_103),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_103),
.Y(n_290)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_104),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_105),
.B(n_305),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_107),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_156),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_108),
.A2(n_109),
.B1(n_156),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_136),
.B1(n_146),
.B2(n_149),
.Y(n_109)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_110),
.B(n_149),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_110),
.A2(n_327),
.B1(n_336),
.B2(n_344),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_110),
.A2(n_146),
.B1(n_423),
.B2(n_426),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_110),
.A2(n_146),
.B1(n_327),
.B2(n_426),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_110),
.A2(n_344),
.B1(n_543),
.B2(n_544),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_125),
.Y(n_110)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_119),
.B2(n_122),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_117),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_118),
.Y(n_323)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_119),
.Y(n_311)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_121),
.Y(n_471)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_132),
.B2(n_134),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_134),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_136),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_139),
.Y(n_337)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_141),
.Y(n_331)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_141),
.Y(n_335)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_142),
.Y(n_427)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_148),
.B(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_154),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_156),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_165),
.B1(n_172),
.B2(n_178),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_157),
.A2(n_165),
.B1(n_276),
.B2(n_284),
.Y(n_275)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_161),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_206),
.B(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_165),
.A2(n_431),
.B1(n_437),
.B2(n_438),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_165),
.A2(n_448),
.B1(n_463),
.B2(n_466),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_167),
.Y(n_316)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_171),
.Y(n_283)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_171),
.Y(n_320)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_171),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_214),
.B1(n_244),
.B2(n_245),
.Y(n_181)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_182),
.B(n_245),
.C(n_559),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_204),
.B1(n_205),
.B2(n_213),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_183),
.B(n_205),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_194),
.B2(n_203),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_184),
.A2(n_203),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_184),
.A2(n_203),
.B1(n_381),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_194),
.Y(n_543)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_198),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_203),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_203),
.B(n_305),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_204),
.A2(n_205),
.B1(n_550),
.B2(n_551),
.Y(n_549)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_231),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_216),
.B(n_231),
.C(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_221),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_222),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_226),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B(n_235),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_233),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_243),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_237),
.A2(n_308),
.B1(n_314),
.B2(n_317),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_237),
.A2(n_277),
.B1(n_317),
.B2(n_375),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_237),
.A2(n_447),
.B1(n_452),
.B2(n_456),
.Y(n_446)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g437 ( 
.A(n_240),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_240),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_242),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.C(n_251),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_247),
.B(n_249),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_251),
.B(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_261),
.C(n_286),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_252),
.A2(n_286),
.B1(n_287),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_252),
.Y(n_510)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_253),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_261),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_275),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_262),
.B(n_275),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_268),
.Y(n_366)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_281),
.Y(n_400)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_504),
.B(n_518),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_486),
.B(n_503),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_389),
.B(n_485),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_360),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_297),
.B(n_360),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_326),
.C(n_345),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_298),
.B(n_482),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_307),
.B1(n_324),
.B2(n_325),
.Y(n_298)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_299),
.B(n_325),
.Y(n_378)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_305),
.B(n_407),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_SL g423 ( 
.A1(n_305),
.A2(n_406),
.B(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_305),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_308),
.Y(n_438)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_309),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_320),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_326),
.A2(n_345),
.B1(n_346),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_326),
.Y(n_483)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_376),
.B2(n_377),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_361),
.B(n_379),
.C(n_387),
.Y(n_502)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_370),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_363),
.B(n_372),
.C(n_373),
.Y(n_490)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_387),
.B2(n_388),
.Y(n_377)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_479),
.B(n_484),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_444),
.B(n_478),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_429),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_392),
.B(n_429),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_421),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_421),
.B1(n_422),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_397),
.A3(n_401),
.B1(n_406),
.B2(n_409),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_398),
.B(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_415),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_439),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_441),
.C(n_443),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_439)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_459),
.B(n_477),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_457),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_457),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_473),
.B(n_476),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.Y(n_460)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_464),
.Y(n_472)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_474),
.B(n_475),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_SL g484 ( 
.A(n_480),
.B(n_481),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_502),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_502),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_491),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_489),
.B(n_490),
.C(n_491),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_497),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_495),
.C(n_497),
.Y(n_513)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_507),
.B(n_514),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_507),
.C(n_519),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_511),
.C(n_513),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_508),
.B(n_517),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_SL g517 ( 
.A(n_511),
.B(n_513),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_516),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_560),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_558),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_525),
.B(n_558),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_528),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_546),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_530),
.A2(n_542),
.B(n_545),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_542),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_547),
.A2(n_548),
.B1(n_549),
.B2(n_557),
.Y(n_546)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_547),
.Y(n_557)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx3_ASAP7_75t_SL g555 ( 
.A(n_556),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);


endmodule