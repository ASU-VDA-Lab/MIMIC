module fake_ibex_1411_n_4073 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_898, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4073);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4073;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3674;
wire n_3255;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3904;
wire n_3135;
wire n_3440;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_3711;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3668;
wire n_3699;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3874;
wire n_1281;
wire n_3094;
wire n_3217;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_1237;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3855;
wire n_3357;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_3578;
wire n_954;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_1395;
wire n_998;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_4047;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_3557;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3682;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3434;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_961;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3745;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3333;
wire n_3096;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_3604;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_1542;
wire n_1586;
wire n_1362;
wire n_946;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_2207;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_3143;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_1193;
wire n_980;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_4038;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2148;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_3247;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g899 ( 
.A(n_701),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_878),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_849),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_884),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_77),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_76),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_828),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_808),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_308),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_192),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_862),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_561),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_816),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_174),
.Y(n_912)
);

BUFx5_ASAP7_75t_L g913 ( 
.A(n_199),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_143),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_155),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_36),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_53),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_395),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_664),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_187),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_792),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_173),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_323),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_306),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_516),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_655),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_774),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_345),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_1),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_783),
.Y(n_930)
);

CKINVDCx16_ASAP7_75t_R g931 ( 
.A(n_826),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_240),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_162),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_192),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_178),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_564),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_417),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_209),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_622),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_475),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_807),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_795),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_433),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_722),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_235),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_879),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_847),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_726),
.Y(n_948)
);

CKINVDCx14_ASAP7_75t_R g949 ( 
.A(n_654),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_817),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_378),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_791),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_431),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_72),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_861),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_90),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_283),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_864),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_755),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_861),
.Y(n_960)
);

CKINVDCx16_ASAP7_75t_R g961 ( 
.A(n_7),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_831),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_615),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_803),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_889),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_860),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_829),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_364),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_586),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_837),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_220),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_473),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_594),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_142),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_431),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_309),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_877),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_57),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_113),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_799),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_801),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_78),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_697),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_789),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_537),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_830),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_887),
.Y(n_987)
);

BUFx10_ASAP7_75t_L g988 ( 
.A(n_808),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_513),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_479),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_592),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_175),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_19),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_369),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_73),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_553),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_480),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_330),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_608),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_527),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_309),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_139),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_331),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_78),
.Y(n_1004)
);

BUFx2_ASAP7_75t_SL g1005 ( 
.A(n_402),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_276),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_677),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_835),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_819),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_441),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_814),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_129),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_351),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_401),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_654),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_830),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_599),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_795),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_550),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_534),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_841),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_886),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_55),
.Y(n_1023)
);

CKINVDCx16_ASAP7_75t_R g1024 ( 
.A(n_765),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_416),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_840),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_809),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_239),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_809),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_875),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_890),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_194),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_161),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_621),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_832),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_4),
.Y(n_1036)
);

CKINVDCx14_ASAP7_75t_R g1037 ( 
.A(n_524),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_317),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_383),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_130),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_64),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_63),
.Y(n_1042)
);

CKINVDCx16_ASAP7_75t_R g1043 ( 
.A(n_291),
.Y(n_1043)
);

CKINVDCx14_ASAP7_75t_R g1044 ( 
.A(n_689),
.Y(n_1044)
);

BUFx10_ASAP7_75t_L g1045 ( 
.A(n_128),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_888),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_857),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_5),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_512),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_199),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_603),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_713),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_787),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_884),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_834),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_855),
.Y(n_1056)
);

BUFx8_ASAP7_75t_SL g1057 ( 
.A(n_842),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_687),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_827),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_847),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_851),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_896),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_614),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_401),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_785),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_346),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_38),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_676),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_476),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_286),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_558),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_496),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_112),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_372),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_866),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_307),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_15),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_793),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_70),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_303),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_639),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_695),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_826),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_481),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_299),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_855),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_794),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_100),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_812),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_638),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_349),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_850),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_150),
.Y(n_1093)
);

INVxp33_ASAP7_75t_R g1094 ( 
.A(n_66),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_290),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_225),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_56),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_805),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_871),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_82),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_215),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_432),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_816),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_345),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_246),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_292),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_160),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_844),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_104),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_806),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_557),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_880),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_883),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_606),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_430),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_16),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_820),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_257),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_839),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_634),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_641),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_20),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_143),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_800),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_413),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_898),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_77),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_48),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_498),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_819),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_140),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_887),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_718),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_169),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_768),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_736),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_311),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_625),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_386),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_318),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_559),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_790),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_112),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_876),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_120),
.Y(n_1145)
);

BUFx2_ASAP7_75t_SL g1146 ( 
.A(n_758),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_635),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_167),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_768),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_751),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_603),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_541),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_312),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_55),
.Y(n_1154)
);

BUFx10_ASAP7_75t_L g1155 ( 
.A(n_778),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_823),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_314),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_878),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_443),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_856),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_352),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_843),
.Y(n_1162)
);

CKINVDCx16_ASAP7_75t_R g1163 ( 
.A(n_359),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_281),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_414),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_849),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_859),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_222),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_270),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_252),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_865),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_244),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_39),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_153),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_818),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_602),
.Y(n_1176)
);

BUFx5_ASAP7_75t_L g1177 ( 
.A(n_692),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_852),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_657),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_383),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_822),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_893),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_470),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_5),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_597),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_482),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_546),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_395),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_390),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_811),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_707),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_712),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_297),
.Y(n_1193)
);

BUFx5_ASAP7_75t_L g1194 ( 
.A(n_845),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_859),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_838),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_639),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_186),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_885),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_881),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_778),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_700),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_109),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_853),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_134),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_606),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_518),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_862),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_725),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_869),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_306),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_412),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_118),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_18),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_570),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_467),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_824),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_400),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_868),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_821),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_698),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_355),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_892),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_488),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_767),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_152),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_895),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_198),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_561),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_873),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_439),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_409),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_846),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_577),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_786),
.Y(n_1235)
);

BUFx2_ASAP7_75t_SL g1236 ( 
.A(n_867),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_90),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_634),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_270),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_280),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_310),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_858),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_874),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_662),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_832),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_136),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_709),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_159),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_320),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_213),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_765),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_854),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_118),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_548),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_38),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_863),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_49),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_897),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_872),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_187),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_572),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_209),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_100),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_371),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_279),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_796),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_276),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_339),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_447),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_376),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_143),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_356),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_810),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_805),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_51),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_664),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_804),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_41),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_215),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_482),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_836),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_798),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_681),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_271),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_896),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_68),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_833),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_848),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_717),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_825),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_188),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_422),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_40),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_264),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_335),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_699),
.Y(n_1296)
);

CKINVDCx16_ASAP7_75t_R g1297 ( 
.A(n_579),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_792),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_411),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_894),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_815),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_720),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_26),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_524),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_298),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_263),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_756),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_191),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_39),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_802),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_628),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_258),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_286),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_453),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_870),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_784),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_619),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_85),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_715),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_788),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_797),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_882),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_756),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_690),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_782),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_891),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_319),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_83),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_813),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_452),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_116),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_959),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_959),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_922),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_939),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1066),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_941),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1001),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1177),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1129),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1231),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1010),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_949),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_949),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1037),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1260),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_900),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1263),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1051),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_976),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1293),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_907),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_900),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_903),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_910),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_989),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_914),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_920),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_923),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_967),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_924),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1075),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_915),
.Y(n_1363)
);

INVxp33_ASAP7_75t_SL g1364 ( 
.A(n_1199),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1075),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_938),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_967),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1044),
.Y(n_1368)
);

CKINVDCx14_ASAP7_75t_R g1369 ( 
.A(n_1044),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_956),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_957),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_989),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_971),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1087),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1087),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_985),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_968),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_938),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1057),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_995),
.Y(n_1380)
);

CKINVDCx16_ASAP7_75t_R g1381 ( 
.A(n_961),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1252),
.Y(n_1382)
);

CKINVDCx16_ASAP7_75t_R g1383 ( 
.A(n_1043),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_997),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_992),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1002),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1057),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1014),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1017),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1108),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1019),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1020),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1177),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1177),
.Y(n_1394)
);

INVxp33_ASAP7_75t_L g1395 ( 
.A(n_899),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1023),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1003),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1025),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1034),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1039),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1032),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1110),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1042),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1048),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1049),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1088),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1095),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1110),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1000),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1096),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1097),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1102),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1003),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1164),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1164),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1106),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1168),
.Y(n_1417)
);

INVxp33_ASAP7_75t_L g1418 ( 
.A(n_905),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1120),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1121),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_941),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1032),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1128),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1131),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1138),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1036),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1139),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1153),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1289),
.B(n_0),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1154),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1161),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1273),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1174),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1185),
.Y(n_1434)
);

BUFx8_ASAP7_75t_L g1435 ( 
.A(n_1390),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1362),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1372),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1352),
.B(n_1163),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1364),
.A2(n_1241),
.B1(n_1297),
.B2(n_1211),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1366),
.A2(n_1328),
.B1(n_908),
.B2(n_912),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1337),
.Y(n_1441)
);

AOI22x1_ASAP7_75t_SL g1442 ( 
.A1(n_1378),
.A2(n_902),
.B1(n_1182),
.B2(n_1149),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1365),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1377),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1351),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1374),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1375),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1377),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1372),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1339),
.A2(n_1006),
.B(n_945),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1413),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1338),
.B(n_1287),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1402),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1337),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1342),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1432),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1334),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1393),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1394),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1349),
.B(n_1107),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1382),
.B(n_1045),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1343),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1332),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1354),
.A2(n_1070),
.B(n_1063),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1333),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1335),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1336),
.Y(n_1468)
);

CKINVDCx16_ASAP7_75t_R g1469 ( 
.A(n_1381),
.Y(n_1469)
);

NOR2x1_ASAP7_75t_L g1470 ( 
.A(n_1350),
.B(n_1157),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1383),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1355),
.A2(n_1070),
.B(n_1063),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1340),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1385),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1421),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1341),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1397),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1356),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1344),
.A2(n_917),
.B1(n_918),
.B2(n_916),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1346),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1348),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1426),
.B(n_919),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1357),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1369),
.A2(n_926),
.B1(n_928),
.B2(n_925),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1358),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1359),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1361),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1347),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_L g1489 ( 
.A(n_1353),
.B(n_913),
.Y(n_1489)
);

AND2x2_ASAP7_75t_SL g1490 ( 
.A(n_1434),
.B(n_931),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1370),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1401),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1371),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1373),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1422),
.B(n_1137),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1376),
.Y(n_1496)
);

CKINVDCx6p67_ASAP7_75t_R g1497 ( 
.A(n_1409),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1360),
.A2(n_932),
.B1(n_933),
.B2(n_929),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1380),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1387),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1384),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1386),
.B(n_935),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1388),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1389),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1395),
.B(n_1137),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1391),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1392),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1396),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1414),
.A2(n_904),
.B1(n_951),
.B2(n_943),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1367),
.B(n_1165),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1398),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1399),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1400),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1403),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1404),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1405),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1415),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1406),
.A2(n_1079),
.B(n_1071),
.Y(n_1518)
);

CKINVDCx6p67_ASAP7_75t_R g1519 ( 
.A(n_1417),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1407),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1418),
.B(n_1410),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1411),
.A2(n_936),
.B1(n_940),
.B2(n_937),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1429),
.B(n_1248),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1412),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1416),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1419),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1420),
.B(n_1024),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1423),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1424),
.Y(n_1529)
);

AND2x6_ASAP7_75t_L g1530 ( 
.A(n_1425),
.B(n_1268),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1427),
.B(n_1158),
.Y(n_1531)
);

INVxp33_ASAP7_75t_SL g1532 ( 
.A(n_1428),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1430),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1431),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1433),
.B(n_953),
.Y(n_1535)
);

INVx5_ASAP7_75t_L g1536 ( 
.A(n_1372),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1345),
.B(n_954),
.Y(n_1537)
);

AND2x6_ASAP7_75t_L g1538 ( 
.A(n_1372),
.B(n_1269),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1337),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1351),
.B(n_1308),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1362),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1362),
.Y(n_1542)
);

CKINVDCx8_ASAP7_75t_R g1543 ( 
.A(n_1363),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1345),
.B(n_1285),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1368),
.B(n_901),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1363),
.Y(n_1546)
);

INVx6_ASAP7_75t_L g1547 ( 
.A(n_1363),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1337),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1379),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1364),
.A2(n_969),
.B1(n_972),
.B2(n_963),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1362),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1352),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1345),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1372),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1337),
.Y(n_1555)
);

CKINVDCx6p67_ASAP7_75t_R g1556 ( 
.A(n_1363),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1368),
.B(n_909),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1351),
.B(n_913),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1337),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1362),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1372),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1351),
.B(n_913),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1338),
.A2(n_973),
.B1(n_978),
.B2(n_974),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1352),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1379),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1368),
.B(n_909),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1345),
.B(n_979),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1368),
.B(n_1029),
.Y(n_1568)
);

INVx6_ASAP7_75t_L g1569 ( 
.A(n_1363),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1352),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1362),
.Y(n_1571)
);

OAI22x1_ASAP7_75t_L g1572 ( 
.A1(n_1379),
.A2(n_1094),
.B1(n_991),
.B2(n_994),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1352),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1345),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1352),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1337),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1372),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1345),
.B(n_990),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1362),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1337),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1362),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1362),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1364),
.A2(n_998),
.B1(n_999),
.B2(n_996),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1345),
.B(n_1004),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1362),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1362),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1337),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1337),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1368),
.B(n_1196),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1362),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1337),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1372),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1556),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1497),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1519),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1465),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1472),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1473),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1519),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1546),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1469),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1521),
.B(n_934),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1458),
.Y(n_1603)
);

BUFx10_ASAP7_75t_L g1604 ( 
.A(n_1547),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1467),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1445),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_SL g1607 ( 
.A(n_1490),
.Y(n_1607)
);

NOR2xp67_ASAP7_75t_L g1608 ( 
.A(n_1471),
.B(n_0),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1476),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1435),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1569),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1543),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1543),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1494),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_R g1615 ( 
.A(n_1500),
.B(n_1549),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1505),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1565),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1517),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1456),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1518),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1530),
.B(n_1071),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1511),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_R g1623 ( 
.A(n_1526),
.B(n_1012),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1514),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1528),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1442),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1533),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1450),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1440),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1509),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1532),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1483),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1480),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1508),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1481),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1574),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1488),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1563),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1492),
.Y(n_1639)
);

AND2x6_ASAP7_75t_L g1640 ( 
.A(n_1527),
.B(n_1558),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1439),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1484),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1479),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1550),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1464),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1583),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1462),
.B(n_975),
.Y(n_1647)
);

CKINVDCx20_ASAP7_75t_R g1648 ( 
.A(n_1553),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1522),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1466),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1572),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1485),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1538),
.Y(n_1653)
);

CKINVDCx16_ASAP7_75t_R g1654 ( 
.A(n_1495),
.Y(n_1654)
);

AND3x2_ASAP7_75t_L g1655 ( 
.A(n_1540),
.B(n_1080),
.C(n_1069),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1498),
.Y(n_1656)
);

BUFx10_ASAP7_75t_L g1657 ( 
.A(n_1544),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1561),
.B(n_1013),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1438),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1463),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1504),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1507),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1478),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1502),
.A2(n_1216),
.B(n_1193),
.Y(n_1664)
);

INVxp33_ASAP7_75t_L g1665 ( 
.A(n_1452),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1437),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1577),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1537),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1516),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1538),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1538),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1468),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1489),
.B(n_1084),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1510),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1457),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_SL g1676 ( 
.A(n_1530),
.B(n_1090),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1525),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1567),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1578),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1584),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_R g1681 ( 
.A(n_1449),
.B(n_1091),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1529),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1482),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1536),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1536),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1474),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1562),
.B(n_913),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1477),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1554),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1534),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1534),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1461),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1535),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1561),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1592),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1592),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1444),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1448),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1436),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1523),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_R g1701 ( 
.A(n_1451),
.B(n_1122),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1552),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1443),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1564),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1491),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1486),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1446),
.Y(n_1707)
);

CKINVDCx16_ASAP7_75t_R g1708 ( 
.A(n_1545),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1570),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1447),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1573),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1575),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1453),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1487),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1493),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1496),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1499),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1557),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1503),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1566),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1501),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1568),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_R g1723 ( 
.A(n_1531),
.B(n_1125),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1589),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_R g1725 ( 
.A(n_1512),
.B(n_1127),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1454),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1506),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1513),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1515),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1541),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1524),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1542),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1551),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1560),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1470),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1571),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_R g1737 ( 
.A(n_1520),
.B(n_1212),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1579),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1581),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1582),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1585),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1586),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1590),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1459),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1460),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1441),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1441),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1455),
.Y(n_1748)
);

XNOR2xp5_ASAP7_75t_L g1749 ( 
.A(n_1455),
.B(n_1228),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1475),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1475),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1539),
.Y(n_1752)
);

CKINVDCx20_ASAP7_75t_R g1753 ( 
.A(n_1548),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1555),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1559),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1559),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1576),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1580),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1587),
.Y(n_1759)
);

BUFx10_ASAP7_75t_L g1760 ( 
.A(n_1588),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1591),
.A2(n_1237),
.B(n_1232),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1473),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1473),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_R g1764 ( 
.A(n_1546),
.B(n_1028),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_R g1765 ( 
.A(n_1546),
.B(n_1250),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1556),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1497),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1480),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1445),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1445),
.Y(n_1770)
);

CKINVDCx16_ASAP7_75t_R g1771 ( 
.A(n_1469),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1473),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1547),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1556),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1556),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1556),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1659),
.A2(n_1305),
.B1(n_1317),
.B2(n_1303),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1596),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1728),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1611),
.B(n_965),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1679),
.B(n_1770),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1753),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1705),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1745),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1597),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1610),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1598),
.Y(n_1787)
);

XOR2xp5_ASAP7_75t_L g1788 ( 
.A(n_1648),
.B(n_1016),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1620),
.Y(n_1789)
);

AND2x2_ASAP7_75t_SL g1790 ( 
.A(n_1676),
.B(n_1018),
.Y(n_1790)
);

AO22x2_ASAP7_75t_L g1791 ( 
.A1(n_1725),
.A2(n_1005),
.B1(n_1236),
.B2(n_1146),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1737),
.Y(n_1792)
);

AND2x2_ASAP7_75t_SL g1793 ( 
.A(n_1771),
.B(n_1026),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1604),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1693),
.B(n_1038),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1769),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1616),
.B(n_1040),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1762),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1634),
.B(n_1050),
.Y(n_1799)
);

INVx6_ASAP7_75t_L g1800 ( 
.A(n_1604),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1773),
.B(n_1053),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1623),
.A2(n_1065),
.B1(n_1083),
.B2(n_1055),
.Y(n_1802)
);

BUFx8_ASAP7_75t_SL g1803 ( 
.A(n_1594),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1619),
.Y(n_1804)
);

INVx5_ASAP7_75t_L g1805 ( 
.A(n_1760),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1647),
.B(n_982),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1639),
.B(n_1221),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1675),
.B(n_1033),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1772),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1615),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_SL g1812 ( 
.A(n_1735),
.Y(n_1812)
);

INVx4_ASAP7_75t_SL g1813 ( 
.A(n_1607),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1703),
.Y(n_1814)
);

INVx4_ASAP7_75t_L g1815 ( 
.A(n_1660),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1672),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1721),
.Y(n_1817)
);

AND2x6_ASAP7_75t_L g1818 ( 
.A(n_1614),
.B(n_993),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1640),
.A2(n_1712),
.B1(n_1686),
.B2(n_1688),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1617),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1699),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1602),
.B(n_1744),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1758),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1640),
.B(n_1067),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1706),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1637),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1714),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1715),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1707),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1710),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1749),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1665),
.B(n_1072),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1701),
.B(n_1073),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_SL g1834 ( 
.A(n_1765),
.B(n_1076),
.C(n_1074),
.Y(n_1834)
);

NOR3xp33_ASAP7_75t_L g1835 ( 
.A(n_1708),
.B(n_1147),
.C(n_1143),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1723),
.B(n_1077),
.Y(n_1836)
);

BUFx4f_ASAP7_75t_L g1837 ( 
.A(n_1640),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1761),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1640),
.B(n_1081),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1713),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1681),
.Y(n_1841)
);

INVx4_ASAP7_75t_L g1842 ( 
.A(n_1593),
.Y(n_1842)
);

INVx6_ASAP7_75t_L g1843 ( 
.A(n_1760),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1664),
.B(n_1716),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1717),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1657),
.B(n_1085),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1719),
.Y(n_1847)
);

INVx4_ASAP7_75t_SL g1848 ( 
.A(n_1607),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1727),
.B(n_1100),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1635),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1683),
.B(n_1104),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1729),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1731),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1670),
.B(n_1109),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1657),
.B(n_1114),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1726),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1608),
.B(n_1196),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1645),
.B(n_1116),
.Y(n_1858)
);

AND2x6_ASAP7_75t_L g1859 ( 
.A(n_1622),
.B(n_993),
.Y(n_1859)
);

NAND2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1603),
.B(n_1148),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1650),
.B(n_1118),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1768),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1599),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1768),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1776),
.B(n_1124),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1766),
.B(n_1123),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1718),
.Y(n_1867)
);

BUFx8_ASAP7_75t_SL g1868 ( 
.A(n_1767),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1605),
.B(n_906),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1666),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1601),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1730),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1739),
.Y(n_1873)
);

INVx2_ASAP7_75t_SL g1874 ( 
.A(n_1667),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1668),
.B(n_1134),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1618),
.B(n_1151),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1624),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1678),
.B(n_1140),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1720),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1625),
.Y(n_1880)
);

AND2x6_ASAP7_75t_L g1881 ( 
.A(n_1627),
.B(n_993),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1702),
.B(n_1141),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1774),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1687),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1761),
.Y(n_1885)
);

INVxp33_ASAP7_75t_L g1886 ( 
.A(n_1673),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1658),
.B(n_1609),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1722),
.B(n_1152),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1628),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1775),
.B(n_1162),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1628),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1724),
.Y(n_1892)
);

AND2x2_ASAP7_75t_SL g1893 ( 
.A(n_1655),
.B(n_1093),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1680),
.B(n_1638),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1628),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1663),
.Y(n_1896)
);

OR2x6_ASAP7_75t_L g1897 ( 
.A(n_1621),
.B(n_1245),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1684),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1671),
.B(n_1159),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1649),
.A2(n_1172),
.B1(n_1173),
.B2(n_1170),
.Y(n_1900)
);

NAND2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1677),
.B(n_1330),
.Y(n_1901)
);

XOR2xp5_ASAP7_75t_L g1902 ( 
.A(n_1641),
.B(n_1176),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1709),
.B(n_1179),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1711),
.A2(n_1184),
.B1(n_1186),
.B2(n_1180),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1633),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1697),
.A2(n_1188),
.B1(n_1189),
.B2(n_1187),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1694),
.B(n_911),
.Y(n_1907)
);

INVx4_ASAP7_75t_L g1908 ( 
.A(n_1612),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1613),
.B(n_1171),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1644),
.B(n_1203),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1732),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1733),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1738),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1734),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1736),
.B(n_1205),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1740),
.B(n_1206),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1700),
.B(n_1692),
.Y(n_1917)
);

NAND2x1p5_ASAP7_75t_L g1918 ( 
.A(n_1690),
.B(n_1756),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1646),
.B(n_1213),
.Y(n_1919)
);

INVxp67_ASAP7_75t_SL g1920 ( 
.A(n_1764),
.Y(n_1920)
);

BUFx2_ASAP7_75t_L g1921 ( 
.A(n_1698),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1600),
.B(n_1215),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1751),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1741),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1642),
.A2(n_988),
.B1(n_1155),
.B2(n_947),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1643),
.B(n_1218),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1742),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1752),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1695),
.B(n_1222),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1632),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1743),
.B(n_1224),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1595),
.B(n_1202),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1652),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_SL g1934 ( 
.A(n_1626),
.Y(n_1934)
);

INVx2_ASAP7_75t_SL g1935 ( 
.A(n_1696),
.Y(n_1935)
);

BUFx10_ASAP7_75t_L g1936 ( 
.A(n_1674),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1661),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1704),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1689),
.B(n_1229),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1685),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1759),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1656),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1662),
.B(n_1234),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1630),
.B(n_1283),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1669),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1682),
.A2(n_1240),
.B1(n_1244),
.B2(n_1238),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1757),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1691),
.Y(n_1948)
);

INVx4_ASAP7_75t_L g1949 ( 
.A(n_1651),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1748),
.B(n_1246),
.Y(n_1950)
);

INVx4_ASAP7_75t_L g1951 ( 
.A(n_1629),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1754),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1746),
.Y(n_1953)
);

AO22x2_ASAP7_75t_L g1954 ( 
.A1(n_1755),
.A2(n_1296),
.B1(n_952),
.B2(n_958),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1747),
.B(n_1270),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1611),
.B(n_946),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1596),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1611),
.B(n_962),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1596),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1604),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1596),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_L g1962 ( 
.A(n_1653),
.B(n_1276),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1596),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1596),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1604),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1606),
.B(n_1327),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1636),
.B(n_1267),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1728),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1615),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1654),
.B(n_1272),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1604),
.Y(n_1971)
);

AND2x6_ASAP7_75t_L g1972 ( 
.A(n_1596),
.B(n_993),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1728),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1728),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1636),
.B(n_1275),
.Y(n_1975)
);

AND2x6_ASAP7_75t_L g1976 ( 
.A(n_1596),
.B(n_1015),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1728),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_SL g1978 ( 
.A(n_1631),
.B(n_1278),
.Y(n_1978)
);

AND2x6_ASAP7_75t_L g1979 ( 
.A(n_1596),
.B(n_1015),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1596),
.Y(n_1980)
);

INVxp33_ASAP7_75t_L g1981 ( 
.A(n_1725),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1659),
.B(n_1331),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1636),
.B(n_1280),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1728),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1606),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1728),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1606),
.B(n_1284),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1728),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1640),
.A2(n_1294),
.B1(n_1295),
.B2(n_1286),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1604),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1728),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1753),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1728),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1604),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1611),
.B(n_966),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1596),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1728),
.Y(n_1997)
);

OR2x6_ASAP7_75t_L g1998 ( 
.A(n_1610),
.B(n_1301),
.Y(n_1998)
);

INVx4_ASAP7_75t_L g1999 ( 
.A(n_1610),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1604),
.Y(n_2000)
);

INVx5_ASAP7_75t_L g2001 ( 
.A(n_1750),
.Y(n_2001)
);

BUFx12f_ASAP7_75t_L g2002 ( 
.A(n_1811),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1778),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1815),
.B(n_980),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_2001),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1779),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1796),
.Y(n_2007)
);

AO22x2_ASAP7_75t_L g2008 ( 
.A1(n_1777),
.A2(n_1254),
.B1(n_1255),
.B2(n_1253),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1785),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_2001),
.B(n_983),
.Y(n_2010)
);

NAND2x1p5_ASAP7_75t_L g2011 ( 
.A(n_1805),
.B(n_1015),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_R g2012 ( 
.A(n_1969),
.B(n_1299),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1960),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1968),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1973),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1974),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1960),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1807),
.B(n_1304),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1805),
.B(n_1816),
.Y(n_2019)
);

NAND2x1p5_ASAP7_75t_L g2020 ( 
.A(n_1965),
.B(n_1041),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1977),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1984),
.Y(n_2022)
);

AO22x2_ASAP7_75t_L g2023 ( 
.A1(n_1788),
.A2(n_1262),
.B1(n_1264),
.B2(n_1257),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1986),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1988),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1789),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1985),
.B(n_1265),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1990),
.B(n_1041),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1813),
.B(n_1007),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1990),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1991),
.Y(n_2031)
);

INVxp67_ASAP7_75t_L g2032 ( 
.A(n_1978),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1851),
.A2(n_927),
.B1(n_930),
.B2(n_921),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1822),
.B(n_1271),
.Y(n_2034)
);

NAND3xp33_ASAP7_75t_L g2035 ( 
.A(n_1882),
.B(n_1064),
.C(n_1041),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1993),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1813),
.B(n_1009),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1997),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1967),
.B(n_1279),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1784),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1873),
.Y(n_2041)
);

INVxp67_ASAP7_75t_SL g2042 ( 
.A(n_1938),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1975),
.B(n_1291),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1983),
.B(n_1292),
.Y(n_2044)
);

AO22x2_ASAP7_75t_L g2045 ( 
.A1(n_1792),
.A2(n_1312),
.B1(n_1313),
.B2(n_1311),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1848),
.B(n_1022),
.Y(n_2046)
);

AO22x2_ASAP7_75t_L g2047 ( 
.A1(n_1817),
.A2(n_1318),
.B1(n_1314),
.B2(n_1046),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1787),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1848),
.B(n_1031),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1926),
.B(n_988),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1957),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1888),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1935),
.B(n_1047),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_1835),
.A2(n_944),
.B1(n_950),
.B2(n_948),
.C(n_942),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1800),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1959),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1798),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1837),
.A2(n_1105),
.B1(n_1115),
.B2(n_1101),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1860),
.B(n_1323),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1961),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1877),
.B(n_1054),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1910),
.B(n_1155),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1806),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1963),
.Y(n_2064)
);

AO22x2_ASAP7_75t_L g2065 ( 
.A1(n_1902),
.A2(n_1068),
.B1(n_1078),
.B2(n_1060),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1810),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1880),
.B(n_1086),
.Y(n_2067)
);

OAI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_1925),
.A2(n_960),
.B1(n_977),
.B2(n_970),
.C(n_955),
.Y(n_2068)
);

NOR3xp33_ASAP7_75t_L g2069 ( 
.A(n_1834),
.B(n_1325),
.C(n_1324),
.Y(n_2069)
);

NAND2x1p5_ASAP7_75t_L g2070 ( 
.A(n_1786),
.B(n_1064),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1964),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1843),
.Y(n_2072)
);

AO22x2_ASAP7_75t_L g2073 ( 
.A1(n_1902),
.A2(n_1099),
.B1(n_1103),
.B2(n_1098),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_1900),
.A2(n_981),
.B1(n_987),
.B2(n_986),
.C(n_984),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1980),
.Y(n_2075)
);

NAND2x1p5_ASAP7_75t_L g2076 ( 
.A(n_1999),
.B(n_1064),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1825),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1844),
.A2(n_1115),
.B1(n_1145),
.B2(n_1105),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1782),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1827),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1874),
.B(n_1117),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1828),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1868),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1919),
.B(n_1191),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1819),
.B(n_1321),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1982),
.B(n_1795),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1843),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1845),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1847),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1928),
.B(n_1119),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1876),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_1921),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1970),
.B(n_1008),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1852),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1853),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1875),
.B(n_1225),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1901),
.B(n_1966),
.Y(n_2097)
);

AO22x2_ASAP7_75t_L g2098 ( 
.A1(n_1942),
.A2(n_1132),
.B1(n_1136),
.B2(n_1130),
.Y(n_2098)
);

AO22x2_ASAP7_75t_L g2099 ( 
.A1(n_1808),
.A2(n_1150),
.B1(n_1160),
.B2(n_1144),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1987),
.B(n_1011),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1996),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1869),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1821),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1829),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1830),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1911),
.B(n_1181),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_1884),
.A2(n_1183),
.B(n_1197),
.C(n_1169),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1912),
.B(n_1192),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1840),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1833),
.B(n_1021),
.Y(n_2110)
);

BUFx8_ASAP7_75t_L g2111 ( 
.A(n_1934),
.Y(n_2111)
);

AO22x2_ASAP7_75t_L g2112 ( 
.A1(n_1920),
.A2(n_1209),
.B1(n_1210),
.B2(n_1200),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1856),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1872),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_1797),
.A2(n_1258),
.B1(n_1251),
.B2(n_1030),
.Y(n_2115)
);

CKINVDCx14_ASAP7_75t_R g2116 ( 
.A(n_1871),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1849),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1867),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1858),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1836),
.B(n_1027),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1861),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1823),
.Y(n_2122)
);

AO22x2_ASAP7_75t_L g2123 ( 
.A1(n_1954),
.A2(n_1219),
.B1(n_1220),
.B2(n_1217),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1878),
.B(n_1035),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1954),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1905),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1943),
.Y(n_2127)
);

BUFx6f_ASAP7_75t_L g2128 ( 
.A(n_1923),
.Y(n_2128)
);

A2O1A1Ixp33_ASAP7_75t_L g2129 ( 
.A1(n_1887),
.A2(n_1169),
.B(n_1197),
.C(n_1183),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_1914),
.B(n_1223),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1933),
.Y(n_2131)
);

BUFx3_ASAP7_75t_L g2132 ( 
.A(n_1992),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1937),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1799),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1945),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1846),
.B(n_1052),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_SL g2137 ( 
.A1(n_1791),
.A2(n_1058),
.B1(n_1061),
.B2(n_1056),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1855),
.B(n_1062),
.Y(n_2138)
);

AO22x1_ASAP7_75t_L g2139 ( 
.A1(n_1981),
.A2(n_1089),
.B1(n_1092),
.B2(n_1082),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1948),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1950),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_1936),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1814),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1989),
.A2(n_1214),
.B1(n_1226),
.B2(n_1198),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1794),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_SL g2146 ( 
.A1(n_1802),
.A2(n_1326),
.B1(n_1112),
.B2(n_1113),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1994),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1952),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1838),
.A2(n_1214),
.B1(n_1226),
.B2(n_1198),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_1906),
.B(n_1126),
.Y(n_2150)
);

AO22x2_ASAP7_75t_L g2151 ( 
.A1(n_1894),
.A2(n_1243),
.B1(n_1259),
.B2(n_1247),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1947),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1904),
.B(n_1133),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1955),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1903),
.B(n_1135),
.Y(n_2155)
);

CKINVDCx11_ASAP7_75t_R g2156 ( 
.A(n_1863),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1947),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1913),
.Y(n_2158)
);

NAND2x1p5_ASAP7_75t_L g2159 ( 
.A(n_2000),
.B(n_1111),
.Y(n_2159)
);

BUFx2_ASAP7_75t_L g2160 ( 
.A(n_1879),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1924),
.B(n_1266),
.Y(n_2161)
);

OR2x2_ASAP7_75t_SL g2162 ( 
.A(n_1831),
.B(n_1870),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1930),
.Y(n_2163)
);

OAI22xp5_ASAP7_75t_SL g2164 ( 
.A1(n_1793),
.A2(n_1319),
.B1(n_1322),
.B2(n_1310),
.Y(n_2164)
);

AND2x2_ASAP7_75t_SL g2165 ( 
.A(n_1893),
.B(n_1239),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1907),
.B(n_1142),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1946),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1824),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1826),
.B(n_1156),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1839),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1971),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1927),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1857),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_SL g2174 ( 
.A1(n_1841),
.A2(n_1166),
.B1(n_1175),
.B2(n_1167),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_1886),
.B(n_1922),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_1892),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_1898),
.B(n_1940),
.Y(n_2177)
);

NAND2x1p5_ASAP7_75t_L g2178 ( 
.A(n_1941),
.B(n_1111),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_L g2179 ( 
.A1(n_1832),
.A2(n_1261),
.B(n_1309),
.C(n_1249),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_1915),
.A2(n_1195),
.B1(n_1201),
.B2(n_1190),
.C(n_1178),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1897),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_1908),
.B(n_1274),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1883),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1916),
.B(n_1204),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1953),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1918),
.Y(n_2186)
);

AND2x4_ASAP7_75t_L g2187 ( 
.A(n_1854),
.B(n_1899),
.Y(n_2187)
);

AO22x2_ASAP7_75t_L g2188 ( 
.A1(n_1896),
.A2(n_1300),
.B1(n_1307),
.B2(n_1290),
.Y(n_2188)
);

INVx2_ASAP7_75t_SL g2189 ( 
.A(n_1820),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1885),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_1780),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1850),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1862),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1864),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_1801),
.Y(n_2195)
);

OAI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_1931),
.A2(n_1227),
.B1(n_1233),
.B2(n_1230),
.C(n_1208),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1998),
.Y(n_2197)
);

CKINVDCx16_ASAP7_75t_R g2198 ( 
.A(n_1842),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_1917),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1812),
.Y(n_2200)
);

AO22x2_ASAP7_75t_L g2201 ( 
.A1(n_1944),
.A2(n_1315),
.B1(n_1301),
.B2(n_1309),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1818),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_1929),
.B(n_1235),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1956),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1958),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1939),
.B(n_1242),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1995),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1909),
.B(n_1256),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1818),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1866),
.Y(n_2210)
);

AND2x6_ASAP7_75t_L g2211 ( 
.A(n_1889),
.B(n_1207),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1865),
.A2(n_1890),
.B1(n_1932),
.B2(n_1951),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_1962),
.Y(n_2213)
);

AO22x2_ASAP7_75t_L g2214 ( 
.A1(n_1949),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1859),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1859),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1859),
.Y(n_2217)
);

OR2x2_ASAP7_75t_SL g2218 ( 
.A(n_1881),
.B(n_1207),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1881),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1881),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1976),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1976),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1979),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_1891),
.A2(n_1281),
.B1(n_1282),
.B2(n_1277),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1979),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_1895),
.B(n_2),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_2001),
.B(n_1207),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1960),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1783),
.B(n_1288),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1779),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1796),
.B(n_1298),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_1783),
.B(n_3),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_1783),
.B(n_3),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_1960),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1779),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1778),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1778),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1779),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1778),
.Y(n_2239)
);

AND2x4_ASAP7_75t_L g2240 ( 
.A(n_1783),
.B(n_4),
.Y(n_2240)
);

NAND2x1p5_ASAP7_75t_L g2241 ( 
.A(n_2001),
.B(n_1306),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_1783),
.B(n_5),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1779),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1779),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_1783),
.B(n_6),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_1783),
.B(n_6),
.Y(n_2246)
);

OR2x2_ASAP7_75t_SL g2247 ( 
.A(n_1834),
.B(n_941),
.Y(n_2247)
);

NOR3xp33_ASAP7_75t_L g2248 ( 
.A(n_1781),
.B(n_1194),
.C(n_8),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1779),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_SL g2250 ( 
.A(n_1863),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1783),
.B(n_7),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1960),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1796),
.B(n_964),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1783),
.B(n_8),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1778),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1779),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1783),
.B(n_8),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1779),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1807),
.B(n_9),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1960),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1779),
.Y(n_2261)
);

AO22x1_ASAP7_75t_L g2262 ( 
.A1(n_1981),
.A2(n_1302),
.B1(n_1316),
.B2(n_1059),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_1783),
.B(n_9),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_1783),
.B(n_9),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1783),
.B(n_10),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1779),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1779),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1779),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1783),
.B(n_10),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_1804),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1779),
.Y(n_2271)
);

INVxp67_ASAP7_75t_L g2272 ( 
.A(n_1804),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1779),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1779),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1779),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_1783),
.B(n_11),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1779),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_1807),
.B(n_11),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_1777),
.B(n_11),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1779),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1779),
.Y(n_2281)
);

A2O1A1Ixp33_ASAP7_75t_L g2282 ( 
.A1(n_1884),
.A2(n_1320),
.B(n_1329),
.C(n_1316),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1778),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1796),
.B(n_1316),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_2001),
.B(n_1320),
.Y(n_2285)
);

INVx8_ASAP7_75t_L g2286 ( 
.A(n_2001),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1779),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_1790),
.A2(n_1329),
.B1(n_1320),
.B2(n_14),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1796),
.B(n_1320),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1796),
.B(n_1329),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1779),
.Y(n_2291)
);

OR2x6_ASAP7_75t_L g2292 ( 
.A(n_1809),
.B(n_12),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1779),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1778),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1779),
.Y(n_2295)
);

OAI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_1777),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1778),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1779),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1779),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_1778),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_1781),
.B(n_16),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_1796),
.B(n_18),
.Y(n_2302)
);

BUFx8_ASAP7_75t_L g2303 ( 
.A(n_1934),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1779),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_1790),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1778),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_1796),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1779),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_1783),
.B(n_17),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1779),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1779),
.Y(n_2311)
);

NOR3xp33_ASAP7_75t_L g2312 ( 
.A(n_1781),
.B(n_24),
.C(n_23),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_2001),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1779),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1779),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1779),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1778),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_1804),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1779),
.Y(n_2319)
);

OAI221xp5_ASAP7_75t_L g2320 ( 
.A1(n_1822),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.C(n_25),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1778),
.Y(n_2321)
);

INVxp67_ASAP7_75t_L g2322 ( 
.A(n_1804),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1779),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1779),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1778),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1779),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1779),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_1804),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1779),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1779),
.Y(n_2330)
);

OR2x2_ASAP7_75t_SL g2331 ( 
.A(n_1834),
.B(n_27),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1779),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1783),
.B(n_28),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1779),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_1777),
.B(n_29),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_1807),
.B(n_29),
.Y(n_2336)
);

NAND2x1p5_ASAP7_75t_L g2337 ( 
.A(n_2001),
.B(n_30),
.Y(n_2337)
);

AO22x2_ASAP7_75t_L g2338 ( 
.A1(n_1777),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2338)
);

AO22x2_ASAP7_75t_L g2339 ( 
.A1(n_1777),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_1960),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1779),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_1790),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2342)
);

AO22x2_ASAP7_75t_L g2343 ( 
.A1(n_1777),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_1783),
.B(n_35),
.Y(n_2344)
);

OR2x2_ASAP7_75t_SL g2345 ( 
.A(n_1834),
.B(n_36),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_1807),
.B(n_37),
.Y(n_2346)
);

OAI221xp5_ASAP7_75t_L g2347 ( 
.A1(n_1822),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.C(n_41),
.Y(n_2347)
);

AO22x2_ASAP7_75t_L g2348 ( 
.A1(n_1777),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_1960),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_1783),
.B(n_43),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_1803),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2001),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1779),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1783),
.B(n_44),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1779),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1960),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1779),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_1960),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1779),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1779),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1778),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_1884),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1783),
.B(n_46),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1779),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_1796),
.B(n_48),
.Y(n_2365)
);

AO22x2_ASAP7_75t_L g2366 ( 
.A1(n_1777),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_1796),
.Y(n_2367)
);

BUFx3_ASAP7_75t_L g2368 ( 
.A(n_2001),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1778),
.Y(n_2369)
);

OR2x2_ASAP7_75t_SL g2370 ( 
.A(n_1834),
.B(n_50),
.Y(n_2370)
);

NAND2xp33_ASAP7_75t_L g2371 ( 
.A(n_1972),
.B(n_51),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1807),
.B(n_50),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1783),
.B(n_52),
.Y(n_2373)
);

AOI22xp33_ASAP7_75t_L g2374 ( 
.A1(n_1790),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1778),
.Y(n_2375)
);

AOI22xp33_ASAP7_75t_L g2376 ( 
.A1(n_1790),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_1804),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1783),
.B(n_54),
.Y(n_2378)
);

AO22x2_ASAP7_75t_L g2379 ( 
.A1(n_1777),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1779),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1779),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2191),
.B(n_58),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2019),
.B(n_59),
.Y(n_2383)
);

OAI22xp5_ASAP7_75t_L g2384 ( 
.A1(n_2165),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2167),
.B(n_59),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2003),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2117),
.B(n_62),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2091),
.B(n_62),
.Y(n_2388)
);

O2A1O1Ixp33_ASAP7_75t_L g2389 ( 
.A1(n_2086),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2009),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2008),
.B(n_65),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2006),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2119),
.B(n_69),
.Y(n_2393)
);

NAND2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2019),
.B(n_2340),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2371),
.A2(n_71),
.B(n_72),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2121),
.B(n_73),
.Y(n_2396)
);

O2A1O1Ixp33_ASAP7_75t_SL g2397 ( 
.A1(n_2107),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2007),
.Y(n_2398)
);

NAND2x1p5_ASAP7_75t_L g2399 ( 
.A(n_2013),
.B(n_74),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2052),
.B(n_75),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2137),
.B(n_675),
.Y(n_2401)
);

HB1xp67_ASAP7_75t_L g2402 ( 
.A(n_2307),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2134),
.B(n_75),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2160),
.B(n_2032),
.Y(n_2404)
);

A2O1A1Ixp33_ASAP7_75t_L g2405 ( 
.A1(n_2301),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2190),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2026),
.Y(n_2407)
);

AO21x1_ASAP7_75t_L g2408 ( 
.A1(n_2125),
.A2(n_678),
.B(n_677),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2008),
.B(n_84),
.Y(n_2409)
);

AOI21x1_ASAP7_75t_L g2410 ( 
.A1(n_2221),
.A2(n_86),
.B(n_87),
.Y(n_2410)
);

O2A1O1Ixp33_ASAP7_75t_L g2411 ( 
.A1(n_2248),
.A2(n_2302),
.B(n_2365),
.C(n_2179),
.Y(n_2411)
);

O2A1O1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2296),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_2286),
.Y(n_2413)
);

BUFx2_ASAP7_75t_L g2414 ( 
.A(n_2367),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_2017),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_L g2416 ( 
.A1(n_2222),
.A2(n_89),
.B(n_91),
.Y(n_2416)
);

AOI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2190),
.A2(n_91),
.B(n_92),
.Y(n_2417)
);

AOI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2034),
.A2(n_92),
.B(n_93),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2030),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2014),
.B(n_2015),
.Y(n_2420)
);

INVx5_ASAP7_75t_L g2421 ( 
.A(n_2292),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2016),
.B(n_93),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2021),
.B(n_93),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2022),
.B(n_94),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2123),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2092),
.B(n_96),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2024),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2023),
.B(n_97),
.Y(n_2428)
);

OAI21x1_ASAP7_75t_L g2429 ( 
.A1(n_2223),
.A2(n_97),
.B(n_98),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2025),
.B(n_98),
.Y(n_2430)
);

OAI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2141),
.A2(n_99),
.B(n_100),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2127),
.A2(n_99),
.B(n_101),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_SL g2433 ( 
.A(n_2083),
.B(n_101),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2031),
.B(n_2036),
.Y(n_2434)
);

AOI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2023),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2435)
);

O2A1O1Ixp33_ASAP7_75t_L g2436 ( 
.A1(n_2312),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2199),
.B(n_106),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2038),
.B(n_2040),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2123),
.A2(n_2045),
.B1(n_2233),
.B2(n_2232),
.Y(n_2439)
);

AO32x1_ASAP7_75t_L g2440 ( 
.A1(n_2078),
.A2(n_109),
.A3(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2041),
.B(n_107),
.Y(n_2441)
);

BUFx12f_ASAP7_75t_L g2442 ( 
.A(n_2156),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2129),
.A2(n_108),
.B(n_110),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2230),
.B(n_110),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2030),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2235),
.B(n_111),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2238),
.B(n_114),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2051),
.A2(n_115),
.B(n_117),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2056),
.A2(n_117),
.B(n_118),
.Y(n_2449)
);

AOI22x1_ASAP7_75t_L g2450 ( 
.A1(n_2178),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2174),
.B(n_679),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2060),
.A2(n_119),
.B(n_120),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2375),
.A2(n_2071),
.B(n_2064),
.Y(n_2453)
);

A2O1A1Ixp33_ASAP7_75t_L g2454 ( 
.A1(n_2168),
.A2(n_122),
.B(n_119),
.C(n_121),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2098),
.B(n_121),
.Y(n_2455)
);

AOI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2075),
.A2(n_121),
.B(n_122),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2170),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2243),
.B(n_123),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2244),
.B(n_123),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2149),
.A2(n_124),
.B(n_125),
.Y(n_2460)
);

OAI22xp5_ASAP7_75t_L g2461 ( 
.A1(n_2232),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2118),
.B(n_126),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2101),
.A2(n_127),
.B(n_128),
.Y(n_2463)
);

BUFx2_ASAP7_75t_L g2464 ( 
.A(n_2292),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2236),
.A2(n_131),
.B(n_132),
.Y(n_2465)
);

A2O1A1Ixp33_ASAP7_75t_L g2466 ( 
.A1(n_2362),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2249),
.B(n_134),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2237),
.A2(n_135),
.B(n_136),
.Y(n_2468)
);

BUFx6f_ASAP7_75t_L g2469 ( 
.A(n_2228),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2239),
.A2(n_135),
.B(n_137),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2256),
.B(n_137),
.Y(n_2471)
);

BUFx4f_ASAP7_75t_L g2472 ( 
.A(n_2002),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2258),
.B(n_138),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2261),
.B(n_139),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2255),
.A2(n_140),
.B(n_141),
.Y(n_2475)
);

OAI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2240),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2283),
.A2(n_2297),
.B(n_2294),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2234),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2234),
.B(n_144),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2240),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2480)
);

OAI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2251),
.A2(n_145),
.B(n_146),
.Y(n_2481)
);

OAI321xp33_ASAP7_75t_L g2482 ( 
.A1(n_2305),
.A2(n_149),
.A3(n_151),
.B1(n_147),
.B2(n_148),
.C(n_150),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2266),
.B(n_2267),
.Y(n_2483)
);

AOI21xp5_ASAP7_75t_L g2484 ( 
.A1(n_2300),
.A2(n_148),
.B(n_149),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2268),
.Y(n_2485)
);

AOI21xp5_ASAP7_75t_L g2486 ( 
.A1(n_2306),
.A2(n_149),
.B(n_150),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2271),
.B(n_151),
.Y(n_2487)
);

O2A1O1Ixp33_ASAP7_75t_L g2488 ( 
.A1(n_2097),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2273),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2274),
.B(n_152),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2275),
.B(n_2277),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2280),
.B(n_2281),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2242),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2317),
.A2(n_154),
.B(n_155),
.Y(n_2494)
);

OAI22xp5_ASAP7_75t_L g2495 ( 
.A1(n_2242),
.A2(n_2246),
.B1(n_2257),
.B2(n_2245),
.Y(n_2495)
);

AO32x1_ASAP7_75t_L g2496 ( 
.A1(n_2225),
.A2(n_158),
.A3(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2287),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2321),
.A2(n_156),
.B(n_157),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2291),
.Y(n_2499)
);

NAND2x1p5_ASAP7_75t_L g2500 ( 
.A(n_2252),
.B(n_160),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2047),
.B(n_160),
.Y(n_2501)
);

O2A1O1Ixp33_ASAP7_75t_L g2502 ( 
.A1(n_2054),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2325),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_L g2504 ( 
.A(n_2342),
.B(n_163),
.C(n_164),
.Y(n_2504)
);

NOR2x1_ASAP7_75t_L g2505 ( 
.A(n_2005),
.B(n_164),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2212),
.B(n_680),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2293),
.B(n_165),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2295),
.B(n_166),
.Y(n_2508)
);

NOR2x1_ASAP7_75t_R g2509 ( 
.A(n_2351),
.B(n_166),
.Y(n_2509)
);

AOI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2262),
.A2(n_167),
.B(n_168),
.Y(n_2510)
);

A2O1A1Ixp33_ASAP7_75t_L g2511 ( 
.A1(n_2320),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2511)
);

AOI21x1_ASAP7_75t_L g2512 ( 
.A1(n_2253),
.A2(n_168),
.B(n_169),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2176),
.B(n_170),
.Y(n_2513)
);

BUFx8_ASAP7_75t_L g2514 ( 
.A(n_2250),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_2361),
.A2(n_170),
.B(n_171),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2369),
.A2(n_171),
.B(n_172),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2298),
.B(n_171),
.Y(n_2517)
);

AOI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_2282),
.A2(n_172),
.B(n_173),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_L g2519 ( 
.A1(n_2065),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2519)
);

AOI21xp5_ASAP7_75t_L g2520 ( 
.A1(n_2105),
.A2(n_2265),
.B(n_2254),
.Y(n_2520)
);

AOI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2269),
.A2(n_175),
.B(n_176),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2299),
.B(n_177),
.Y(n_2522)
);

O2A1O1Ixp33_ASAP7_75t_L g2523 ( 
.A1(n_2120),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2304),
.B(n_179),
.Y(n_2524)
);

O2A1O1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2110),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2252),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2308),
.B(n_181),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2065),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2270),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2310),
.B(n_182),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2311),
.Y(n_2531)
);

O2A1O1Ixp33_ASAP7_75t_L g2532 ( 
.A1(n_2039),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2333),
.A2(n_188),
.B(n_189),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2314),
.B(n_188),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2315),
.B(n_189),
.Y(n_2535)
);

NAND3xp33_ASAP7_75t_L g2536 ( 
.A(n_2035),
.B(n_190),
.C(n_191),
.Y(n_2536)
);

OR2x4_ASAP7_75t_L g2537 ( 
.A(n_2279),
.B(n_190),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_2260),
.Y(n_2538)
);

NAND2x1_ASAP7_75t_L g2539 ( 
.A(n_2211),
.B(n_2202),
.Y(n_2539)
);

AOI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2354),
.A2(n_193),
.B(n_194),
.Y(n_2540)
);

OAI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2363),
.A2(n_2378),
.B(n_2373),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2103),
.A2(n_2109),
.B(n_2104),
.Y(n_2542)
);

AOI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2113),
.A2(n_2114),
.B(n_2044),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2048),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2159),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2316),
.B(n_193),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2043),
.A2(n_195),
.B(n_196),
.Y(n_2547)
);

A2O1A1Ixp33_ASAP7_75t_L g2548 ( 
.A1(n_2347),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2319),
.B(n_195),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2163),
.A2(n_196),
.B(n_197),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_SL g2551 ( 
.A(n_2288),
.B(n_200),
.C(n_201),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_L g2552 ( 
.A1(n_2073),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2245),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_2553)
);

O2A1O1Ixp33_ASAP7_75t_L g2554 ( 
.A1(n_2018),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2323),
.B(n_205),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2073),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2324),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2047),
.B(n_208),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2326),
.B(n_209),
.Y(n_2559)
);

AOI21x1_ASAP7_75t_L g2560 ( 
.A1(n_2284),
.A2(n_210),
.B(n_211),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2327),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_2011),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2289),
.A2(n_210),
.B(n_211),
.Y(n_2563)
);

O2A1O1Ixp33_ASAP7_75t_L g2564 ( 
.A1(n_2100),
.A2(n_2335),
.B(n_2196),
.C(n_2180),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2329),
.B(n_212),
.Y(n_2565)
);

AOI21x1_ASAP7_75t_L g2566 ( 
.A1(n_2290),
.A2(n_214),
.B(n_216),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2349),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2349),
.B(n_682),
.Y(n_2568)
);

AOI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2135),
.A2(n_217),
.B(n_218),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2356),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2330),
.B(n_218),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2188),
.B(n_218),
.Y(n_2572)
);

AND2x2_ASAP7_75t_SL g2573 ( 
.A(n_2198),
.B(n_219),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2166),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2332),
.B(n_222),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2155),
.A2(n_223),
.B(n_224),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2334),
.Y(n_2577)
);

OAI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2184),
.A2(n_225),
.B(n_226),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2341),
.B(n_226),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2353),
.B(n_226),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2355),
.Y(n_2581)
);

OAI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2027),
.A2(n_2229),
.B(n_2063),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2357),
.B(n_227),
.Y(n_2583)
);

O2A1O1Ixp5_ASAP7_75t_L g2584 ( 
.A1(n_2085),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2359),
.B(n_227),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2360),
.Y(n_2586)
);

AOI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2140),
.A2(n_228),
.B(n_229),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_2227),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2057),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2128),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2364),
.B(n_230),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2188),
.B(n_231),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2380),
.B(n_2381),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2185),
.A2(n_231),
.B(n_232),
.Y(n_2594)
);

INVx2_ASAP7_75t_SL g2595 ( 
.A(n_2128),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2197),
.B(n_2195),
.Y(n_2596)
);

AOI21x1_ASAP7_75t_L g2597 ( 
.A1(n_2215),
.A2(n_2217),
.B(n_2216),
.Y(n_2597)
);

OAI21x1_ASAP7_75t_L g2598 ( 
.A1(n_2285),
.A2(n_233),
.B(n_234),
.Y(n_2598)
);

AO22x1_ASAP7_75t_L g2599 ( 
.A1(n_2111),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2126),
.A2(n_236),
.B(n_237),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2259),
.B(n_237),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2066),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2278),
.B(n_2336),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2131),
.A2(n_238),
.B(n_239),
.Y(n_2604)
);

INVxp67_ASAP7_75t_L g2605 ( 
.A(n_2272),
.Y(n_2605)
);

AOI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2124),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2133),
.A2(n_241),
.B(n_242),
.Y(n_2607)
);

O2A1O1Ixp33_ASAP7_75t_SL g2608 ( 
.A1(n_2213),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_2608)
);

AND2x6_ASAP7_75t_L g2609 ( 
.A(n_2246),
.B(n_245),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2257),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2241),
.B(n_683),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2346),
.B(n_248),
.Y(n_2612)
);

O2A1O1Ixp33_ASAP7_75t_L g2613 ( 
.A1(n_2136),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_L g2614 ( 
.A(n_2318),
.B(n_252),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2077),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2053),
.B(n_684),
.Y(n_2616)
);

OAI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2080),
.A2(n_253),
.B(n_254),
.Y(n_2617)
);

OAI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2082),
.A2(n_254),
.B(n_255),
.Y(n_2618)
);

BUFx8_ASAP7_75t_L g2619 ( 
.A(n_2158),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2322),
.Y(n_2620)
);

INVx5_ASAP7_75t_L g2621 ( 
.A(n_2183),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2328),
.B(n_256),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2372),
.B(n_256),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2053),
.B(n_685),
.Y(n_2624)
);

BUFx4f_ASAP7_75t_L g2625 ( 
.A(n_2337),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2088),
.A2(n_258),
.B(n_259),
.Y(n_2626)
);

O2A1O1Ixp33_ASAP7_75t_SL g2627 ( 
.A1(n_2219),
.A2(n_2059),
.B(n_2220),
.C(n_2209),
.Y(n_2627)
);

INVx1_ASAP7_75t_SL g2628 ( 
.A(n_2313),
.Y(n_2628)
);

AND2x4_ASAP7_75t_L g2629 ( 
.A(n_2187),
.B(n_260),
.Y(n_2629)
);

AOI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2089),
.A2(n_260),
.B(n_261),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2094),
.A2(n_261),
.B(n_262),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2095),
.A2(n_262),
.B(n_263),
.Y(n_2632)
);

INVx6_ASAP7_75t_L g2633 ( 
.A(n_2183),
.Y(n_2633)
);

AOI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2138),
.A2(n_265),
.B(n_266),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2172),
.B(n_267),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2070),
.B(n_685),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2263),
.A2(n_271),
.B1(n_268),
.B2(n_269),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2264),
.Y(n_2638)
);

CKINVDCx16_ASAP7_75t_R g2639 ( 
.A(n_2012),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2146),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2226),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2377),
.B(n_272),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2264),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2152),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2276),
.Y(n_2645)
);

AO22x1_ASAP7_75t_L g2646 ( 
.A1(n_2303),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2076),
.B(n_686),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2276),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2309),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2102),
.B(n_280),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2050),
.B(n_282),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2309),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2148),
.B(n_2061),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2061),
.B(n_284),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2067),
.B(n_285),
.Y(n_2655)
);

AOI21x1_ASAP7_75t_L g2656 ( 
.A1(n_2144),
.A2(n_287),
.B(n_288),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2344),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2152),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2344),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2350),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2154),
.A2(n_287),
.B(n_288),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2067),
.B(n_287),
.Y(n_2662)
);

INVx3_ASAP7_75t_L g2663 ( 
.A(n_2157),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2151),
.B(n_288),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2062),
.B(n_289),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2350),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2218),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2157),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2084),
.B(n_292),
.Y(n_2669)
);

OAI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2374),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_2670)
);

AOI21x1_ASAP7_75t_L g2671 ( 
.A1(n_2058),
.A2(n_295),
.B(n_296),
.Y(n_2671)
);

OAI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2153),
.A2(n_295),
.B(n_296),
.Y(n_2672)
);

A2O1A1Ixp33_ASAP7_75t_L g2673 ( 
.A1(n_2376),
.A2(n_301),
.B(n_299),
.C(n_300),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2224),
.A2(n_299),
.B(n_300),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2143),
.A2(n_301),
.B(n_302),
.Y(n_2675)
);

O2A1O1Ixp33_ASAP7_75t_L g2676 ( 
.A1(n_2208),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2150),
.B(n_304),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2096),
.B(n_2106),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2175),
.B(n_307),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2106),
.B(n_309),
.Y(n_2680)
);

INVxp67_ASAP7_75t_L g2681 ( 
.A(n_2204),
.Y(n_2681)
);

OAI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2093),
.A2(n_312),
.B(n_313),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2108),
.B(n_2130),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2081),
.B(n_688),
.Y(n_2684)
);

OA21x2_ASAP7_75t_L g2685 ( 
.A1(n_2181),
.A2(n_313),
.B(n_314),
.Y(n_2685)
);

AOI21xp5_ASAP7_75t_L g2686 ( 
.A1(n_2192),
.A2(n_315),
.B(n_316),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2201),
.A2(n_2099),
.B1(n_2379),
.B2(n_2366),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2193),
.A2(n_315),
.B(n_316),
.Y(n_2688)
);

OAI22xp5_ASAP7_75t_SL g2689 ( 
.A1(n_2162),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2689)
);

INVx3_ASAP7_75t_L g2690 ( 
.A(n_2352),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2338),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_2691)
);

O2A1O1Ixp5_ASAP7_75t_L g2692 ( 
.A1(n_2173),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_2692)
);

O2A1O1Ixp33_ASAP7_75t_L g2693 ( 
.A1(n_2069),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2693)
);

AOI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2194),
.A2(n_326),
.B(n_328),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2132),
.Y(n_2695)
);

INVx5_ASAP7_75t_L g2696 ( 
.A(n_2202),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2161),
.B(n_328),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2161),
.B(n_329),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2211),
.Y(n_2699)
);

NOR3xp33_ASAP7_75t_L g2700 ( 
.A(n_2139),
.B(n_330),
.C(n_331),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2169),
.A2(n_331),
.B(n_332),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2171),
.B(n_688),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2339),
.A2(n_2379),
.B1(n_2348),
.B2(n_2366),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2420),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2495),
.A2(n_2247),
.B1(n_2112),
.B2(n_2343),
.Y(n_2705)
);

INVx5_ASAP7_75t_L g2706 ( 
.A(n_2413),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2501),
.B(n_2343),
.Y(n_2707)
);

INVxp67_ASAP7_75t_L g2708 ( 
.A(n_2620),
.Y(n_2708)
);

OAI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2439),
.A2(n_2112),
.B1(n_2348),
.B2(n_2214),
.Y(n_2709)
);

OAI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2537),
.A2(n_2214),
.B1(n_2345),
.B2(n_2331),
.Y(n_2710)
);

AO32x1_ASAP7_75t_L g2711 ( 
.A1(n_2703),
.A2(n_2189),
.A3(n_2142),
.B1(n_2370),
.B2(n_2200),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2464),
.B(n_2042),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_R g2713 ( 
.A(n_2639),
.B(n_2116),
.Y(n_2713)
);

XOR2x2_ASAP7_75t_L g2714 ( 
.A(n_2573),
.B(n_2164),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2392),
.B(n_2205),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2434),
.Y(n_2716)
);

OAI22x1_ASAP7_75t_L g2717 ( 
.A1(n_2421),
.A2(n_2210),
.B1(n_2122),
.B2(n_2079),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2678),
.B(n_2079),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2544),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2413),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2438),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2683),
.B(n_2090),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2558),
.B(n_2010),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2589),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2406),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2419),
.B(n_2186),
.Y(n_2726)
);

NOR3xp33_ASAP7_75t_L g2727 ( 
.A(n_2689),
.B(n_2068),
.C(n_2231),
.Y(n_2727)
);

OAI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2411),
.A2(n_2115),
.B(n_2033),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2427),
.B(n_2207),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2625),
.B(n_2667),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2483),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2398),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2541),
.A2(n_2028),
.B(n_2020),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2414),
.Y(n_2734)
);

O2A1O1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2687),
.A2(n_2074),
.B(n_2182),
.C(n_2203),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2491),
.Y(n_2736)
);

HB1xp67_ASAP7_75t_L g2737 ( 
.A(n_2402),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2485),
.B(n_2489),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2492),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2602),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2419),
.B(n_2368),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2406),
.Y(n_2742)
);

AOI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2453),
.A2(n_2211),
.B(n_2010),
.Y(n_2743)
);

AOI21xp5_ASAP7_75t_L g2744 ( 
.A1(n_2477),
.A2(n_2206),
.B(n_2004),
.Y(n_2744)
);

O2A1O1Ixp5_ASAP7_75t_L g2745 ( 
.A1(n_2506),
.A2(n_2037),
.B(n_2046),
.C(n_2029),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2593),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2419),
.B(n_2469),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2572),
.B(n_2592),
.Y(n_2748)
);

AOI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2627),
.A2(n_2049),
.B(n_2046),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2497),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2543),
.A2(n_2542),
.B(n_2582),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2499),
.B(n_2177),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2615),
.Y(n_2753)
);

AOI21x1_ASAP7_75t_L g2754 ( 
.A1(n_2597),
.A2(n_2087),
.B(n_2358),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2531),
.B(n_2145),
.Y(n_2755)
);

O2A1O1Ixp33_ASAP7_75t_L g2756 ( 
.A1(n_2564),
.A2(n_2147),
.B(n_2072),
.C(n_2055),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2557),
.Y(n_2757)
);

CKINVDCx20_ASAP7_75t_R g2758 ( 
.A(n_2619),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2394),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2406),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2653),
.B(n_333),
.Y(n_2761)
);

A2O1A1Ixp33_ASAP7_75t_L g2762 ( 
.A1(n_2674),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_2762)
);

A2O1A1Ixp33_ASAP7_75t_SL g2763 ( 
.A1(n_2700),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_2763)
);

OAI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2435),
.A2(n_340),
.B1(n_337),
.B2(n_338),
.Y(n_2764)
);

O2A1O1Ixp33_ASAP7_75t_L g2765 ( 
.A1(n_2511),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2561),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2428),
.B(n_342),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2469),
.B(n_343),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2455),
.B(n_344),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2577),
.B(n_2581),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2386),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2514),
.Y(n_2772)
);

A2O1A1Ixp33_ASAP7_75t_L g2773 ( 
.A1(n_2412),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2390),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2407),
.Y(n_2775)
);

AOI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2611),
.A2(n_347),
.B(n_348),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2586),
.B(n_349),
.Y(n_2777)
);

O2A1O1Ixp33_ASAP7_75t_L g2778 ( 
.A1(n_2548),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2478),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2397),
.A2(n_350),
.B(n_352),
.Y(n_2780)
);

BUFx24_ASAP7_75t_SL g2781 ( 
.A(n_2519),
.Y(n_2781)
);

AOI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2539),
.A2(n_353),
.B(n_354),
.Y(n_2782)
);

CKINVDCx6p67_ASAP7_75t_R g2783 ( 
.A(n_2442),
.Y(n_2783)
);

CKINVDCx14_ASAP7_75t_R g2784 ( 
.A(n_2472),
.Y(n_2784)
);

O2A1O1Ixp33_ASAP7_75t_SL g2785 ( 
.A1(n_2405),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_2785)
);

O2A1O1Ixp33_ASAP7_75t_L g2786 ( 
.A1(n_2451),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2529),
.B(n_358),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2605),
.B(n_359),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_SL g2789 ( 
.A(n_2526),
.B(n_360),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2503),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2621),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2677),
.B(n_2651),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2526),
.B(n_2570),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2526),
.Y(n_2794)
);

HB1xp67_ASAP7_75t_L g2795 ( 
.A(n_2383),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2603),
.B(n_361),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_2609),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2636),
.A2(n_362),
.B(n_363),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2422),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2423),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2596),
.B(n_362),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2424),
.Y(n_2802)
);

AOI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2504),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2657),
.B(n_364),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2664),
.B(n_365),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2647),
.A2(n_366),
.B(n_367),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2570),
.Y(n_2807)
);

INVx8_ASAP7_75t_L g2808 ( 
.A(n_2383),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2641),
.A2(n_2443),
.B(n_2699),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2450),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2385),
.A2(n_366),
.B(n_368),
.Y(n_2811)
);

BUFx5_ASAP7_75t_L g2812 ( 
.A(n_2445),
.Y(n_2812)
);

OAI21xp33_ASAP7_75t_L g2813 ( 
.A1(n_2679),
.A2(n_2552),
.B(n_2528),
.Y(n_2813)
);

AOI33xp33_ASAP7_75t_L g2814 ( 
.A1(n_2391),
.A2(n_370),
.A3(n_372),
.B1(n_368),
.B2(n_369),
.B3(n_371),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2388),
.B(n_369),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_2538),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2556),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2633),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2656),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2409),
.B(n_373),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2633),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2638),
.B(n_2645),
.Y(n_2822)
);

AO32x2_ASAP7_75t_L g2823 ( 
.A1(n_2691),
.A2(n_376),
.A3(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2680),
.B(n_374),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2416),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2648),
.B(n_374),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2652),
.B(n_375),
.Y(n_2827)
);

INVx4_ASAP7_75t_L g2828 ( 
.A(n_2696),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2429),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2659),
.B(n_378),
.Y(n_2830)
);

A2O1A1Ixp33_ASAP7_75t_L g2831 ( 
.A1(n_2395),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2629),
.B(n_2400),
.Y(n_2832)
);

BUFx6f_ASAP7_75t_L g2833 ( 
.A(n_2668),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2660),
.B(n_380),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2430),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2668),
.B(n_381),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2666),
.B(n_381),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2588),
.B(n_381),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2481),
.A2(n_382),
.B(n_384),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2668),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2437),
.B(n_384),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2472),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2588),
.B(n_385),
.Y(n_2843)
);

INVx1_ASAP7_75t_SL g2844 ( 
.A(n_2415),
.Y(n_2844)
);

CKINVDCx14_ASAP7_75t_R g2845 ( 
.A(n_2695),
.Y(n_2845)
);

AND2x2_ASAP7_75t_SL g2846 ( 
.A(n_2433),
.B(n_387),
.Y(n_2846)
);

BUFx3_ASAP7_75t_L g2847 ( 
.A(n_2590),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_2562),
.B(n_388),
.Y(n_2848)
);

A2O1A1Ixp33_ASAP7_75t_L g2849 ( 
.A1(n_2502),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_2849)
);

AOI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2608),
.A2(n_391),
.B(n_392),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2614),
.B(n_391),
.Y(n_2851)
);

O2A1O1Ixp33_ASAP7_75t_L g2852 ( 
.A1(n_2616),
.A2(n_2684),
.B(n_2624),
.C(n_2436),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2441),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2545),
.B(n_393),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2598),
.Y(n_2855)
);

AO32x2_ASAP7_75t_L g2856 ( 
.A1(n_2425),
.A2(n_397),
.A3(n_394),
.B1(n_396),
.B2(n_398),
.Y(n_2856)
);

INVx4_ASAP7_75t_L g2857 ( 
.A(n_2696),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2509),
.B(n_394),
.Y(n_2858)
);

OAI22x1_ASAP7_75t_L g2859 ( 
.A1(n_2505),
.A2(n_402),
.B1(n_399),
.B2(n_401),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2681),
.B(n_403),
.Y(n_2860)
);

A2O1A1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2431),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2444),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_L g2863 ( 
.A(n_2696),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2671),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2460),
.A2(n_407),
.B(n_408),
.Y(n_2865)
);

INVx3_ASAP7_75t_L g2866 ( 
.A(n_2690),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2622),
.B(n_409),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2446),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2403),
.B(n_2387),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2393),
.B(n_410),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2396),
.B(n_412),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2447),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2518),
.A2(n_414),
.B(n_415),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2644),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2595),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_2697),
.B(n_415),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_R g2877 ( 
.A(n_2567),
.B(n_415),
.Y(n_2877)
);

CKINVDCx8_ASAP7_75t_R g2878 ( 
.A(n_2479),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2665),
.B(n_416),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2698),
.B(n_417),
.Y(n_2880)
);

O2A1O1Ixp33_ASAP7_75t_L g2881 ( 
.A1(n_2401),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_2881)
);

NAND2x1_ASAP7_75t_L g2882 ( 
.A(n_2685),
.B(n_418),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2458),
.Y(n_2883)
);

NAND2x1p5_ASAP7_75t_L g2884 ( 
.A(n_2628),
.B(n_419),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2576),
.A2(n_420),
.B(n_421),
.Y(n_2885)
);

AOI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2578),
.A2(n_420),
.B(n_421),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2669),
.B(n_422),
.Y(n_2887)
);

A2O1A1Ixp33_ASAP7_75t_SL g2888 ( 
.A1(n_2672),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_2888)
);

INVx2_ASAP7_75t_SL g2889 ( 
.A(n_2644),
.Y(n_2889)
);

NAND2xp33_ASAP7_75t_L g2890 ( 
.A(n_2399),
.B(n_424),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2404),
.A2(n_425),
.B(n_426),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2462),
.B(n_426),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2459),
.Y(n_2893)
);

OR2x6_ASAP7_75t_L g2894 ( 
.A(n_2599),
.B(n_427),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2410),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2513),
.B(n_428),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2690),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2467),
.B(n_429),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2658),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2471),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2663),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2642),
.B(n_430),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_L g2903 ( 
.A(n_2654),
.B(n_2655),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2473),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2646),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2617),
.B(n_432),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2618),
.A2(n_433),
.B(n_434),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2384),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2662),
.B(n_435),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2474),
.B(n_436),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2487),
.B(n_437),
.Y(n_2911)
);

OAI22x1_ASAP7_75t_L g2912 ( 
.A1(n_2640),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2490),
.B(n_437),
.Y(n_2913)
);

CKINVDCx14_ASAP7_75t_R g2914 ( 
.A(n_2461),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2426),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2507),
.B(n_440),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2508),
.B(n_2517),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2522),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2524),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2584),
.A2(n_441),
.B(n_442),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2527),
.Y(n_2921)
);

OAI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2673),
.A2(n_442),
.B(n_443),
.Y(n_2922)
);

A2O1A1Ixp33_ASAP7_75t_L g2923 ( 
.A1(n_2389),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2574),
.B(n_444),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2500),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2530),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2534),
.B(n_447),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2512),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2535),
.B(n_448),
.Y(n_2929)
);

INVx3_ASAP7_75t_L g2930 ( 
.A(n_2560),
.Y(n_2930)
);

AOI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2466),
.A2(n_448),
.B(n_449),
.Y(n_2931)
);

A2O1A1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2613),
.A2(n_2554),
.B(n_2532),
.C(n_2523),
.Y(n_2932)
);

BUFx2_ASAP7_75t_L g2933 ( 
.A(n_2546),
.Y(n_2933)
);

AOI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2440),
.A2(n_450),
.B(n_451),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2566),
.Y(n_2935)
);

A2O1A1Ixp33_ASAP7_75t_L g2936 ( 
.A1(n_2525),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_2936)
);

BUFx2_ASAP7_75t_L g2937 ( 
.A(n_2549),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2555),
.B(n_2559),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2440),
.A2(n_454),
.B(n_455),
.Y(n_2939)
);

OAI21x1_ASAP7_75t_L g2940 ( 
.A1(n_2510),
.A2(n_457),
.B(n_456),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2565),
.B(n_455),
.Y(n_2941)
);

A2O1A1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2693),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2571),
.Y(n_2943)
);

NOR3xp33_ASAP7_75t_L g2944 ( 
.A(n_2702),
.B(n_458),
.C(n_459),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2575),
.B(n_460),
.Y(n_2945)
);

BUFx3_ASAP7_75t_L g2946 ( 
.A(n_2382),
.Y(n_2946)
);

A2O1A1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2676),
.A2(n_2418),
.B(n_2488),
.C(n_2634),
.Y(n_2947)
);

OAI21x1_ASAP7_75t_L g2948 ( 
.A1(n_2417),
.A2(n_462),
.B(n_461),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2601),
.B(n_461),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2579),
.Y(n_2950)
);

AOI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2551),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2580),
.B(n_465),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2583),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2585),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2606),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2591),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2496),
.A2(n_466),
.B(n_467),
.Y(n_2957)
);

O2A1O1Ixp33_ASAP7_75t_L g2958 ( 
.A1(n_2454),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_2958)
);

NOR3xp33_ASAP7_75t_L g2959 ( 
.A(n_2476),
.B(n_468),
.C(n_469),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2496),
.A2(n_469),
.B(n_470),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2521),
.A2(n_471),
.B(n_472),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2685),
.Y(n_2962)
);

HB1xp67_ASAP7_75t_L g2963 ( 
.A(n_2480),
.Y(n_2963)
);

A2O1A1Ixp33_ASAP7_75t_L g2964 ( 
.A1(n_2547),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2612),
.B(n_473),
.Y(n_2965)
);

AOI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2408),
.A2(n_693),
.B(n_691),
.Y(n_2966)
);

INVx3_ASAP7_75t_L g2967 ( 
.A(n_2635),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2623),
.B(n_2650),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2493),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_2969)
);

BUFx8_ASAP7_75t_L g2970 ( 
.A(n_2553),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2610),
.A2(n_483),
.B1(n_480),
.B2(n_481),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2692),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2432),
.B(n_484),
.Y(n_2973)
);

AND2x4_ASAP7_75t_L g2974 ( 
.A(n_2533),
.B(n_485),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2568),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2540),
.B(n_486),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2536),
.Y(n_2977)
);

BUFx2_ASAP7_75t_SL g2978 ( 
.A(n_2637),
.Y(n_2978)
);

AND2x2_ASAP7_75t_SL g2979 ( 
.A(n_2643),
.B(n_486),
.Y(n_2979)
);

O2A1O1Ixp33_ASAP7_75t_L g2980 ( 
.A1(n_2457),
.A2(n_489),
.B(n_487),
.C(n_488),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2649),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2701),
.B(n_490),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2482),
.B(n_490),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2670),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_2984)
);

INVxp67_ASAP7_75t_L g2985 ( 
.A(n_2563),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2600),
.Y(n_2986)
);

OAI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2569),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2587),
.B(n_494),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2626),
.B(n_495),
.Y(n_2989)
);

OAI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2630),
.A2(n_497),
.B1(n_495),
.B2(n_496),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2631),
.B(n_2632),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2604),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2607),
.Y(n_2993)
);

OAI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2675),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_2994)
);

A2O1A1Ixp33_ASAP7_75t_L g2995 ( 
.A1(n_2661),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2594),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2686),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2688),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_2998)
);

BUFx2_ASAP7_75t_L g2999 ( 
.A(n_2448),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2694),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_3000)
);

CKINVDCx20_ASAP7_75t_R g3001 ( 
.A(n_2449),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2452),
.B(n_505),
.Y(n_3002)
);

OAI22xp5_ASAP7_75t_SL g3003 ( 
.A1(n_2456),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2463),
.B(n_508),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2465),
.B(n_509),
.Y(n_3005)
);

AOI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_2468),
.A2(n_509),
.B(n_510),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2470),
.B(n_510),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2475),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2484),
.A2(n_511),
.B(n_512),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2486),
.B(n_511),
.Y(n_3010)
);

AOI22xp5_ASAP7_75t_L g3011 ( 
.A1(n_2494),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_3011)
);

CKINVDCx11_ASAP7_75t_R g3012 ( 
.A(n_2498),
.Y(n_3012)
);

BUFx12f_ASAP7_75t_L g3013 ( 
.A(n_2515),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2516),
.B(n_514),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_SL g3015 ( 
.A1(n_2550),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_3015)
);

A2O1A1Ixp33_ASAP7_75t_L g3016 ( 
.A1(n_2682),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_3016)
);

A2O1A1Ixp33_ASAP7_75t_L g3017 ( 
.A1(n_2682),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2520),
.A2(n_519),
.B(n_520),
.Y(n_3018)
);

AO21x1_ASAP7_75t_L g3019 ( 
.A1(n_2703),
.A2(n_520),
.B(n_521),
.Y(n_3019)
);

BUFx4f_ASAP7_75t_L g3020 ( 
.A(n_2442),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_2737),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2771),
.Y(n_3022)
);

BUFx2_ASAP7_75t_SL g3023 ( 
.A(n_2758),
.Y(n_3023)
);

INVx5_ASAP7_75t_SL g3024 ( 
.A(n_2783),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2750),
.Y(n_3025)
);

NAND2x1p5_ASAP7_75t_L g3026 ( 
.A(n_2706),
.B(n_520),
.Y(n_3026)
);

OAI22xp5_ASAP7_75t_SL g3027 ( 
.A1(n_2846),
.A2(n_2914),
.B1(n_2784),
.B2(n_2845),
.Y(n_3027)
);

BUFx2_ASAP7_75t_L g3028 ( 
.A(n_2808),
.Y(n_3028)
);

INVx4_ASAP7_75t_L g3029 ( 
.A(n_2842),
.Y(n_3029)
);

BUFx6f_ASAP7_75t_L g3030 ( 
.A(n_2863),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2704),
.B(n_521),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2716),
.B(n_521),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2721),
.B(n_522),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2757),
.Y(n_3034)
);

INVx3_ASAP7_75t_L g3035 ( 
.A(n_2791),
.Y(n_3035)
);

AOI22xp33_ASAP7_75t_L g3036 ( 
.A1(n_2978),
.A2(n_525),
.B1(n_522),
.B2(n_523),
.Y(n_3036)
);

BUFx6f_ASAP7_75t_L g3037 ( 
.A(n_2863),
.Y(n_3037)
);

CKINVDCx20_ASAP7_75t_R g3038 ( 
.A(n_2772),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2863),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2731),
.B(n_2736),
.Y(n_3040)
);

INVx6_ASAP7_75t_L g3041 ( 
.A(n_2791),
.Y(n_3041)
);

INVx5_ASAP7_75t_L g3042 ( 
.A(n_2720),
.Y(n_3042)
);

BUFx3_ASAP7_75t_L g3043 ( 
.A(n_2847),
.Y(n_3043)
);

INVx1_ASAP7_75t_SL g3044 ( 
.A(n_2844),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_2816),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2759),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2739),
.B(n_522),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2875),
.Y(n_3048)
);

BUFx5_ASAP7_75t_L g3049 ( 
.A(n_2741),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_3020),
.Y(n_3050)
);

BUFx6f_ASAP7_75t_L g3051 ( 
.A(n_2725),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2748),
.B(n_523),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2970),
.A2(n_526),
.B1(n_523),
.B2(n_525),
.Y(n_3053)
);

CKINVDCx8_ASAP7_75t_R g3054 ( 
.A(n_2894),
.Y(n_3054)
);

INVx1_ASAP7_75t_SL g3055 ( 
.A(n_2713),
.Y(n_3055)
);

INVx2_ASAP7_75t_SL g3056 ( 
.A(n_2741),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2818),
.Y(n_3057)
);

INVx1_ASAP7_75t_SL g3058 ( 
.A(n_2877),
.Y(n_3058)
);

AND2x2_ASAP7_75t_SL g3059 ( 
.A(n_2858),
.B(n_2979),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2821),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2767),
.B(n_526),
.Y(n_3061)
);

INVx5_ASAP7_75t_L g3062 ( 
.A(n_2828),
.Y(n_3062)
);

CKINVDCx8_ASAP7_75t_R g3063 ( 
.A(n_2894),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2774),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2775),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2766),
.Y(n_3066)
);

NAND2x1p5_ASAP7_75t_L g3067 ( 
.A(n_2857),
.B(n_527),
.Y(n_3067)
);

NAND2x1_ASAP7_75t_L g3068 ( 
.A(n_2836),
.B(n_528),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2805),
.B(n_2820),
.Y(n_3069)
);

AOI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_2792),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_3070)
);

INVx5_ASAP7_75t_L g3071 ( 
.A(n_2725),
.Y(n_3071)
);

BUFx2_ASAP7_75t_L g3072 ( 
.A(n_2779),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2738),
.Y(n_3073)
);

CKINVDCx20_ASAP7_75t_R g3074 ( 
.A(n_2714),
.Y(n_3074)
);

BUFx6f_ASAP7_75t_L g3075 ( 
.A(n_2725),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2770),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_L g3077 ( 
.A(n_2742),
.Y(n_3077)
);

BUFx6f_ASAP7_75t_L g3078 ( 
.A(n_2742),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2719),
.Y(n_3079)
);

INVx3_ASAP7_75t_L g3080 ( 
.A(n_2878),
.Y(n_3080)
);

BUFx2_ASAP7_75t_R g3081 ( 
.A(n_2905),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2732),
.Y(n_3082)
);

INVx1_ASAP7_75t_SL g3083 ( 
.A(n_2734),
.Y(n_3083)
);

BUFx3_ASAP7_75t_L g3084 ( 
.A(n_2726),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2742),
.Y(n_3085)
);

INVx3_ASAP7_75t_SL g3086 ( 
.A(n_2854),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2760),
.Y(n_3087)
);

INVx2_ASAP7_75t_SL g3088 ( 
.A(n_2717),
.Y(n_3088)
);

INVx3_ASAP7_75t_SL g3089 ( 
.A(n_2730),
.Y(n_3089)
);

BUFx6f_ASAP7_75t_L g3090 ( 
.A(n_2760),
.Y(n_3090)
);

INVx6_ASAP7_75t_L g3091 ( 
.A(n_2812),
.Y(n_3091)
);

BUFx6f_ASAP7_75t_L g3092 ( 
.A(n_2760),
.Y(n_3092)
);

INVx6_ASAP7_75t_L g3093 ( 
.A(n_2812),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2813),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2790),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_2866),
.Y(n_3096)
);

INVx6_ASAP7_75t_SL g3097 ( 
.A(n_2836),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2724),
.Y(n_3098)
);

INVxp67_ASAP7_75t_SL g3099 ( 
.A(n_2795),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2709),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2740),
.Y(n_3101)
);

INVx5_ASAP7_75t_L g3102 ( 
.A(n_2794),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2753),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2746),
.B(n_2707),
.Y(n_3104)
);

INVx8_ASAP7_75t_L g3105 ( 
.A(n_2897),
.Y(n_3105)
);

INVx8_ASAP7_75t_L g3106 ( 
.A(n_2874),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2715),
.Y(n_3107)
);

BUFx2_ASAP7_75t_L g3108 ( 
.A(n_2807),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_2925),
.Y(n_3109)
);

AOI22xp33_ASAP7_75t_L g3110 ( 
.A1(n_2710),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_3110)
);

BUFx2_ASAP7_75t_L g3111 ( 
.A(n_2807),
.Y(n_3111)
);

BUFx3_ASAP7_75t_L g3112 ( 
.A(n_2833),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2799),
.B(n_536),
.Y(n_3113)
);

INVx3_ASAP7_75t_SL g3114 ( 
.A(n_2915),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2769),
.B(n_536),
.Y(n_3115)
);

INVx3_ASAP7_75t_L g3116 ( 
.A(n_2925),
.Y(n_3116)
);

CKINVDCx11_ASAP7_75t_R g3117 ( 
.A(n_3012),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2874),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2833),
.Y(n_3119)
);

INVx5_ASAP7_75t_L g3120 ( 
.A(n_2840),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2962),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2729),
.Y(n_3122)
);

BUFx4_ASAP7_75t_SL g3123 ( 
.A(n_2946),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2840),
.Y(n_3124)
);

INVx4_ASAP7_75t_L g3125 ( 
.A(n_2874),
.Y(n_3125)
);

BUFx5_ASAP7_75t_L g3126 ( 
.A(n_3013),
.Y(n_3126)
);

AND2x6_ASAP7_75t_L g3127 ( 
.A(n_2855),
.B(n_538),
.Y(n_3127)
);

BUFx12f_ASAP7_75t_L g3128 ( 
.A(n_2884),
.Y(n_3128)
);

INVx4_ASAP7_75t_L g3129 ( 
.A(n_2899),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_2752),
.Y(n_3130)
);

INVx5_ASAP7_75t_L g3131 ( 
.A(n_2889),
.Y(n_3131)
);

INVx1_ASAP7_75t_SL g3132 ( 
.A(n_2712),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2940),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2901),
.Y(n_3134)
);

CKINVDCx5p33_ASAP7_75t_R g3135 ( 
.A(n_2708),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2755),
.Y(n_3136)
);

INVx5_ASAP7_75t_L g3137 ( 
.A(n_2954),
.Y(n_3137)
);

INVx1_ASAP7_75t_SL g3138 ( 
.A(n_2723),
.Y(n_3138)
);

INVx2_ASAP7_75t_SL g3139 ( 
.A(n_2815),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2800),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2802),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2835),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2747),
.Y(n_3143)
);

INVx6_ASAP7_75t_SL g3144 ( 
.A(n_2974),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2777),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2853),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_2705),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2862),
.Y(n_3148)
);

CKINVDCx16_ASAP7_75t_R g3149 ( 
.A(n_2832),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2822),
.Y(n_3150)
);

BUFx6f_ASAP7_75t_L g3151 ( 
.A(n_2793),
.Y(n_3151)
);

BUFx12f_ASAP7_75t_L g3152 ( 
.A(n_2722),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2851),
.B(n_540),
.Y(n_3153)
);

BUFx3_ASAP7_75t_L g3154 ( 
.A(n_2718),
.Y(n_3154)
);

INVx4_ASAP7_75t_L g3155 ( 
.A(n_2933),
.Y(n_3155)
);

NOR2xp67_ASAP7_75t_SL g3156 ( 
.A(n_2983),
.B(n_542),
.Y(n_3156)
);

BUFx6f_ASAP7_75t_L g3157 ( 
.A(n_2954),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_2761),
.Y(n_3158)
);

BUFx6f_ASAP7_75t_L g3159 ( 
.A(n_2975),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2868),
.Y(n_3160)
);

BUFx2_ASAP7_75t_R g3161 ( 
.A(n_2796),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2975),
.Y(n_3162)
);

CKINVDCx6p67_ASAP7_75t_R g3163 ( 
.A(n_2859),
.Y(n_3163)
);

INVx3_ASAP7_75t_L g3164 ( 
.A(n_2975),
.Y(n_3164)
);

BUFx4_ASAP7_75t_SL g3165 ( 
.A(n_3001),
.Y(n_3165)
);

BUFx10_ASAP7_75t_L g3166 ( 
.A(n_2787),
.Y(n_3166)
);

INVx6_ASAP7_75t_SL g3167 ( 
.A(n_2781),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2937),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2956),
.Y(n_3169)
);

BUFx10_ASAP7_75t_L g3170 ( 
.A(n_2788),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2801),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2996),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2872),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2883),
.Y(n_3174)
);

INVx3_ASAP7_75t_L g3175 ( 
.A(n_2967),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2893),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2900),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2904),
.Y(n_3178)
);

INVx2_ASAP7_75t_SL g3179 ( 
.A(n_2867),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2918),
.Y(n_3180)
);

INVxp67_ASAP7_75t_SL g3181 ( 
.A(n_2963),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2919),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2921),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2902),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2926),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2943),
.Y(n_3186)
);

INVx4_ASAP7_75t_L g3187 ( 
.A(n_2924),
.Y(n_3187)
);

INVx2_ASAP7_75t_SL g3188 ( 
.A(n_2824),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2950),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_2880),
.Y(n_3190)
);

INVx1_ASAP7_75t_SL g3191 ( 
.A(n_2890),
.Y(n_3191)
);

OR2x6_ASAP7_75t_L g3192 ( 
.A(n_2749),
.B(n_543),
.Y(n_3192)
);

INVx1_ASAP7_75t_SL g3193 ( 
.A(n_2838),
.Y(n_3193)
);

BUFx6f_ASAP7_75t_L g3194 ( 
.A(n_2996),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2953),
.B(n_543),
.Y(n_3195)
);

INVx2_ASAP7_75t_SL g3196 ( 
.A(n_2843),
.Y(n_3196)
);

INVx2_ASAP7_75t_SL g3197 ( 
.A(n_2848),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2826),
.Y(n_3198)
);

INVx2_ASAP7_75t_SL g3199 ( 
.A(n_2768),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2827),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_L g3201 ( 
.A(n_2996),
.Y(n_3201)
);

BUFx6f_ASAP7_75t_L g3202 ( 
.A(n_2948),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2860),
.Y(n_3203)
);

BUFx2_ASAP7_75t_L g3204 ( 
.A(n_2823),
.Y(n_3204)
);

BUFx2_ASAP7_75t_L g3205 ( 
.A(n_2823),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2981),
.B(n_544),
.Y(n_3206)
);

INVxp67_ASAP7_75t_SL g3207 ( 
.A(n_2751),
.Y(n_3207)
);

INVx5_ASAP7_75t_L g3208 ( 
.A(n_3010),
.Y(n_3208)
);

CKINVDCx6p67_ASAP7_75t_R g3209 ( 
.A(n_2912),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2830),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2834),
.Y(n_3211)
);

BUFx3_ASAP7_75t_L g3212 ( 
.A(n_2949),
.Y(n_3212)
);

INVx5_ASAP7_75t_L g3213 ( 
.A(n_2928),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_SL g3214 ( 
.A(n_2986),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_2965),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2903),
.B(n_544),
.Y(n_3216)
);

BUFx6f_ASAP7_75t_L g3217 ( 
.A(n_2754),
.Y(n_3217)
);

BUFx2_ASAP7_75t_R g3218 ( 
.A(n_2892),
.Y(n_3218)
);

INVx3_ASAP7_75t_L g3219 ( 
.A(n_2882),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2837),
.Y(n_3220)
);

OAI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_2797),
.A2(n_546),
.B1(n_544),
.B2(n_545),
.Y(n_3221)
);

BUFx6f_ASAP7_75t_L g3222 ( 
.A(n_2928),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2928),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2864),
.Y(n_3224)
);

INVx8_ASAP7_75t_L g3225 ( 
.A(n_2756),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_2959),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.Y(n_3226)
);

BUFx3_ASAP7_75t_L g3227 ( 
.A(n_2804),
.Y(n_3227)
);

BUFx6f_ASAP7_75t_L g3228 ( 
.A(n_2935),
.Y(n_3228)
);

BUFx12f_ASAP7_75t_L g3229 ( 
.A(n_2999),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2935),
.Y(n_3230)
);

OR2x6_ASAP7_75t_L g3231 ( 
.A(n_2735),
.B(n_2865),
.Y(n_3231)
);

BUFx2_ASAP7_75t_L g3232 ( 
.A(n_2856),
.Y(n_3232)
);

INVx1_ASAP7_75t_SL g3233 ( 
.A(n_2789),
.Y(n_3233)
);

INVxp67_ASAP7_75t_SL g3234 ( 
.A(n_2743),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2935),
.Y(n_3235)
);

INVx1_ASAP7_75t_SL g3236 ( 
.A(n_2896),
.Y(n_3236)
);

BUFx12f_ASAP7_75t_L g3237 ( 
.A(n_2814),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2841),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3019),
.Y(n_3239)
);

BUFx12f_ASAP7_75t_L g3240 ( 
.A(n_2711),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2819),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2966),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_2976),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2711),
.Y(n_3244)
);

BUFx8_ASAP7_75t_L g3245 ( 
.A(n_2972),
.Y(n_3245)
);

AOI22xp5_ASAP7_75t_L g3246 ( 
.A1(n_2727),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_3246)
);

INVx5_ASAP7_75t_L g3247 ( 
.A(n_2930),
.Y(n_3247)
);

INVxp67_ASAP7_75t_L g3248 ( 
.A(n_2876),
.Y(n_3248)
);

INVx5_ASAP7_75t_L g3249 ( 
.A(n_2977),
.Y(n_3249)
);

NAND2x1p5_ASAP7_75t_L g3250 ( 
.A(n_2803),
.B(n_549),
.Y(n_3250)
);

INVx4_ASAP7_75t_L g3251 ( 
.A(n_2810),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2968),
.B(n_551),
.Y(n_3252)
);

NAND2x1p5_ASAP7_75t_L g3253 ( 
.A(n_2906),
.B(n_551),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_2909),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_2879),
.Y(n_3255)
);

BUFx4f_ASAP7_75t_L g3256 ( 
.A(n_2895),
.Y(n_3256)
);

CKINVDCx11_ASAP7_75t_R g3257 ( 
.A(n_2993),
.Y(n_3257)
);

BUFx3_ASAP7_75t_L g3258 ( 
.A(n_2887),
.Y(n_3258)
);

INVxp67_ASAP7_75t_SL g3259 ( 
.A(n_2825),
.Y(n_3259)
);

INVx4_ASAP7_75t_L g3260 ( 
.A(n_2829),
.Y(n_3260)
);

INVx4_ASAP7_75t_L g3261 ( 
.A(n_2992),
.Y(n_3261)
);

INVx1_ASAP7_75t_SL g3262 ( 
.A(n_2733),
.Y(n_3262)
);

INVx8_ASAP7_75t_L g3263 ( 
.A(n_2745),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2898),
.Y(n_3264)
);

BUFx6f_ASAP7_75t_L g3265 ( 
.A(n_3002),
.Y(n_3265)
);

BUFx3_ASAP7_75t_L g3266 ( 
.A(n_3003),
.Y(n_3266)
);

INVx1_ASAP7_75t_SL g3267 ( 
.A(n_2870),
.Y(n_3267)
);

BUFx10_ASAP7_75t_L g3268 ( 
.A(n_2982),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2869),
.B(n_552),
.Y(n_3269)
);

BUFx6f_ASAP7_75t_L g3270 ( 
.A(n_3007),
.Y(n_3270)
);

BUFx2_ASAP7_75t_L g3271 ( 
.A(n_2985),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2917),
.B(n_553),
.Y(n_3272)
);

BUFx6f_ASAP7_75t_L g3273 ( 
.A(n_3014),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_2764),
.Y(n_3274)
);

NAND2x1p5_ASAP7_75t_L g3275 ( 
.A(n_2908),
.B(n_554),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_2871),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3008),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2938),
.B(n_554),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2910),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2911),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_2973),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_2913),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2916),
.Y(n_3283)
);

INVxp67_ASAP7_75t_SL g3284 ( 
.A(n_2809),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_2988),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_2989),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2927),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2929),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2941),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2945),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2952),
.Y(n_3291)
);

INVx4_ASAP7_75t_L g3292 ( 
.A(n_2944),
.Y(n_3292)
);

OAI21x1_ASAP7_75t_L g3293 ( 
.A1(n_3242),
.A2(n_3133),
.B(n_3219),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3025),
.Y(n_3294)
);

OAI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3059),
.A2(n_2762),
.B(n_3016),
.Y(n_3295)
);

INVx4_ASAP7_75t_SL g3296 ( 
.A(n_3086),
.Y(n_3296)
);

A2O1A1Ixp33_ASAP7_75t_L g3297 ( 
.A1(n_3191),
.A2(n_2786),
.B(n_2881),
.C(n_2839),
.Y(n_3297)
);

OAI21x1_ASAP7_75t_L g3298 ( 
.A1(n_3277),
.A2(n_3241),
.B(n_3224),
.Y(n_3298)
);

AOI221xp5_ASAP7_75t_SL g3299 ( 
.A1(n_3027),
.A2(n_2728),
.B1(n_2817),
.B2(n_2955),
.C(n_2744),
.Y(n_3299)
);

OAI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_3054),
.A2(n_3017),
.B1(n_2951),
.B2(n_2861),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3069),
.B(n_555),
.Y(n_3301)
);

INVx1_ASAP7_75t_SL g3302 ( 
.A(n_3123),
.Y(n_3302)
);

OAI21x1_ASAP7_75t_L g3303 ( 
.A1(n_3207),
.A2(n_2782),
.B(n_2920),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3034),
.Y(n_3304)
);

AO21x2_ASAP7_75t_L g3305 ( 
.A1(n_3244),
.A2(n_2960),
.B(n_2957),
.Y(n_3305)
);

OAI21x1_ASAP7_75t_L g3306 ( 
.A1(n_3035),
.A2(n_3018),
.B(n_2991),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3066),
.Y(n_3307)
);

O2A1O1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_3248),
.A2(n_2763),
.B(n_2888),
.C(n_2932),
.Y(n_3308)
);

OAI221xp5_ASAP7_75t_L g3309 ( 
.A1(n_3054),
.A2(n_2849),
.B1(n_2942),
.B2(n_2773),
.C(n_2922),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_3164),
.A2(n_3284),
.B(n_3124),
.Y(n_3310)
);

OA21x2_ASAP7_75t_L g3311 ( 
.A1(n_3234),
.A2(n_2850),
.B(n_2780),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3022),
.Y(n_3312)
);

OA21x2_ASAP7_75t_L g3313 ( 
.A1(n_3262),
.A2(n_2939),
.B(n_2934),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3256),
.A2(n_2947),
.B(n_2852),
.Y(n_3314)
);

BUFx2_ASAP7_75t_L g3315 ( 
.A(n_3229),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3064),
.Y(n_3316)
);

AND2x4_ASAP7_75t_L g3317 ( 
.A(n_3168),
.B(n_2891),
.Y(n_3317)
);

CKINVDCx20_ASAP7_75t_R g3318 ( 
.A(n_3038),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3160),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3063),
.A2(n_2984),
.B1(n_2831),
.B2(n_2907),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3263),
.A2(n_2886),
.B(n_2885),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3173),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3174),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3065),
.Y(n_3324)
);

OAI21x1_ASAP7_75t_L g3325 ( 
.A1(n_3118),
.A2(n_3005),
.B(n_3004),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3138),
.B(n_556),
.Y(n_3326)
);

OAI21x1_ASAP7_75t_L g3327 ( 
.A1(n_3259),
.A2(n_3068),
.B(n_3121),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3176),
.Y(n_3328)
);

OAI21x1_ASAP7_75t_L g3329 ( 
.A1(n_3239),
.A2(n_3009),
.B(n_3006),
.Y(n_3329)
);

OR2x2_ASAP7_75t_L g3330 ( 
.A(n_3021),
.B(n_557),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3177),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3182),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3095),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3183),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3185),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3186),
.Y(n_3336)
);

OAI21x1_ASAP7_75t_L g3337 ( 
.A1(n_3109),
.A2(n_2776),
.B(n_2931),
.Y(n_3337)
);

BUFx3_ASAP7_75t_L g3338 ( 
.A(n_3043),
.Y(n_3338)
);

OAI21x1_ASAP7_75t_L g3339 ( 
.A1(n_3116),
.A2(n_2806),
.B(n_2798),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_3058),
.B(n_558),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3189),
.Y(n_3341)
);

CKINVDCx6p67_ASAP7_75t_R g3342 ( 
.A(n_3050),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3140),
.Y(n_3343)
);

AND2x4_ASAP7_75t_L g3344 ( 
.A(n_3155),
.B(n_3169),
.Y(n_3344)
);

OAI21x1_ASAP7_75t_SL g3345 ( 
.A1(n_3088),
.A2(n_2980),
.B(n_2958),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3141),
.Y(n_3346)
);

BUFx3_ASAP7_75t_L g3347 ( 
.A(n_3048),
.Y(n_3347)
);

INVx1_ASAP7_75t_SL g3348 ( 
.A(n_3023),
.Y(n_3348)
);

OR2x2_ASAP7_75t_L g3349 ( 
.A(n_3104),
.B(n_559),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3208),
.A2(n_2923),
.B1(n_2936),
.B2(n_3015),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3073),
.B(n_2811),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3076),
.B(n_2969),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3142),
.B(n_2971),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3179),
.B(n_559),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3079),
.Y(n_3355)
);

AO31x2_ASAP7_75t_L g3356 ( 
.A1(n_3260),
.A2(n_2987),
.A3(n_2990),
.B(n_2994),
.Y(n_3356)
);

OAI21x1_ASAP7_75t_L g3357 ( 
.A1(n_3146),
.A2(n_2873),
.B(n_2778),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3184),
.B(n_560),
.Y(n_3358)
);

INVx1_ASAP7_75t_SL g3359 ( 
.A(n_3165),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3148),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3178),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_3149),
.B(n_560),
.Y(n_3362)
);

OAI21x1_ASAP7_75t_L g3363 ( 
.A1(n_3180),
.A2(n_2765),
.B(n_2961),
.Y(n_3363)
);

INVx6_ASAP7_75t_L g3364 ( 
.A(n_3062),
.Y(n_3364)
);

BUFx6f_ASAP7_75t_L g3365 ( 
.A(n_3030),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3098),
.Y(n_3366)
);

OA21x2_ASAP7_75t_L g3367 ( 
.A1(n_3271),
.A2(n_2964),
.B(n_2995),
.Y(n_3367)
);

NOR3xp33_ASAP7_75t_L g3368 ( 
.A(n_3292),
.B(n_3252),
.C(n_3216),
.Y(n_3368)
);

AOI22xp33_ASAP7_75t_L g3369 ( 
.A1(n_3266),
.A2(n_2997),
.B1(n_3000),
.B2(n_2998),
.Y(n_3369)
);

O2A1O1Ixp33_ASAP7_75t_SL g3370 ( 
.A1(n_3055),
.A2(n_3011),
.B(n_564),
.C(n_562),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3101),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3150),
.B(n_2785),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3103),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3040),
.Y(n_3374)
);

INVx4_ASAP7_75t_L g3375 ( 
.A(n_3105),
.Y(n_3375)
);

OAI21x1_ASAP7_75t_L g3376 ( 
.A1(n_3253),
.A2(n_695),
.B(n_694),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3136),
.Y(n_3377)
);

BUFx6f_ASAP7_75t_L g3378 ( 
.A(n_3030),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3130),
.B(n_563),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3107),
.Y(n_3380)
);

OAI21x1_ASAP7_75t_L g3381 ( 
.A1(n_3175),
.A2(n_697),
.B(n_696),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3122),
.B(n_565),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3157),
.Y(n_3383)
);

OAI21x1_ASAP7_75t_L g3384 ( 
.A1(n_3275),
.A2(n_3250),
.B(n_3067),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3157),
.Y(n_3385)
);

BUFx6f_ASAP7_75t_L g3386 ( 
.A(n_3037),
.Y(n_3386)
);

OR2x2_ASAP7_75t_L g3387 ( 
.A(n_3082),
.B(n_566),
.Y(n_3387)
);

OAI21x1_ASAP7_75t_L g3388 ( 
.A1(n_3287),
.A2(n_3288),
.B(n_3026),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3099),
.Y(n_3389)
);

BUFx10_ASAP7_75t_L g3390 ( 
.A(n_3041),
.Y(n_3390)
);

OA21x2_ASAP7_75t_L g3391 ( 
.A1(n_3204),
.A2(n_567),
.B(n_568),
.Y(n_3391)
);

BUFx6f_ASAP7_75t_L g3392 ( 
.A(n_3037),
.Y(n_3392)
);

AND2x4_ASAP7_75t_L g3393 ( 
.A(n_3084),
.B(n_569),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3237),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3394)
);

OAI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_3209),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3052),
.B(n_3154),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_3028),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3181),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3083),
.B(n_573),
.Y(n_3399)
);

AND2x4_ASAP7_75t_L g3400 ( 
.A(n_3045),
.B(n_574),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3134),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3145),
.B(n_574),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3206),
.Y(n_3403)
);

OAI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3246),
.A2(n_575),
.B(n_576),
.Y(n_3404)
);

INVx4_ASAP7_75t_L g3405 ( 
.A(n_3062),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3205),
.Y(n_3406)
);

AO31x2_ASAP7_75t_L g3407 ( 
.A1(n_3261),
.A2(n_578),
.A3(n_576),
.B(n_577),
.Y(n_3407)
);

INVxp67_ASAP7_75t_SL g3408 ( 
.A(n_3072),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_3131),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3232),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3139),
.B(n_578),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3108),
.Y(n_3412)
);

OAI21x1_ASAP7_75t_L g3413 ( 
.A1(n_3031),
.A2(n_702),
.B(n_701),
.Y(n_3413)
);

CKINVDCx6p67_ASAP7_75t_R g3414 ( 
.A(n_3117),
.Y(n_3414)
);

OAI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3094),
.A2(n_580),
.B(n_581),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3053),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_3416)
);

AOI22x1_ASAP7_75t_L g3417 ( 
.A1(n_3128),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3111),
.Y(n_3418)
);

OAI21x1_ASAP7_75t_L g3419 ( 
.A1(n_3032),
.A2(n_3047),
.B(n_3033),
.Y(n_3419)
);

AND2x2_ASAP7_75t_L g3420 ( 
.A(n_3061),
.B(n_583),
.Y(n_3420)
);

OR3x4_ASAP7_75t_SL g3421 ( 
.A(n_3024),
.B(n_584),
.C(n_585),
.Y(n_3421)
);

BUFx2_ASAP7_75t_SL g3422 ( 
.A(n_3029),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3264),
.B(n_587),
.Y(n_3423)
);

AOI21x1_ASAP7_75t_L g3424 ( 
.A1(n_3192),
.A2(n_587),
.B(n_588),
.Y(n_3424)
);

BUFx5_ASAP7_75t_L g3425 ( 
.A(n_3127),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3265),
.Y(n_3426)
);

NAND2x1p5_ASAP7_75t_L g3427 ( 
.A(n_3042),
.B(n_588),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_3161),
.B(n_589),
.Y(n_3428)
);

OAI21x1_ASAP7_75t_L g3429 ( 
.A1(n_3279),
.A2(n_704),
.B(n_703),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3280),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3270),
.Y(n_3431)
);

OR2x2_ASAP7_75t_L g3432 ( 
.A(n_3132),
.B(n_589),
.Y(n_3432)
);

OAI21x1_ASAP7_75t_L g3433 ( 
.A1(n_3283),
.A2(n_705),
.B(n_704),
.Y(n_3433)
);

OAI21x1_ASAP7_75t_L g3434 ( 
.A1(n_3289),
.A2(n_706),
.B(n_705),
.Y(n_3434)
);

BUFx2_ASAP7_75t_L g3435 ( 
.A(n_3144),
.Y(n_3435)
);

AOI21xp33_ASAP7_75t_L g3436 ( 
.A1(n_3225),
.A2(n_590),
.B(n_591),
.Y(n_3436)
);

OAI21x1_ASAP7_75t_L g3437 ( 
.A1(n_3290),
.A2(n_707),
.B(n_706),
.Y(n_3437)
);

AND2x4_ASAP7_75t_L g3438 ( 
.A(n_3056),
.B(n_590),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_3057),
.Y(n_3439)
);

CKINVDCx5p33_ASAP7_75t_R g3440 ( 
.A(n_3114),
.Y(n_3440)
);

BUFx6f_ASAP7_75t_L g3441 ( 
.A(n_3039),
.Y(n_3441)
);

OAI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3187),
.A2(n_596),
.B1(n_593),
.B2(n_595),
.Y(n_3442)
);

OAI21x1_ASAP7_75t_L g3443 ( 
.A1(n_3291),
.A2(n_710),
.B(n_708),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3115),
.B(n_595),
.Y(n_3444)
);

BUFx3_ASAP7_75t_L g3445 ( 
.A(n_3060),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3198),
.B(n_598),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3214),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3273),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_L g3449 ( 
.A1(n_3113),
.A2(n_710),
.B(n_708),
.Y(n_3449)
);

OAI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_3163),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_3450)
);

INVx2_ASAP7_75t_SL g3451 ( 
.A(n_3131),
.Y(n_3451)
);

AND2x4_ASAP7_75t_L g3452 ( 
.A(n_3044),
.B(n_603),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3137),
.Y(n_3453)
);

AO31x2_ASAP7_75t_L g3454 ( 
.A1(n_3251),
.A2(n_607),
.A3(n_604),
.B(n_605),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_3126),
.B(n_604),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3231),
.A2(n_605),
.B(n_607),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3243),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3153),
.B(n_605),
.Y(n_3458)
);

OAI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3070),
.A2(n_608),
.B(n_609),
.Y(n_3459)
);

AOI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3274),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3231),
.A2(n_609),
.B(n_610),
.Y(n_3461)
);

OAI21x1_ASAP7_75t_L g3462 ( 
.A1(n_3195),
.A2(n_714),
.B(n_711),
.Y(n_3462)
);

OA21x2_ASAP7_75t_L g3463 ( 
.A1(n_3147),
.A2(n_3036),
.B(n_3100),
.Y(n_3463)
);

AO21x2_ASAP7_75t_L g3464 ( 
.A1(n_3269),
.A2(n_611),
.B(n_612),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3312),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_L g3466 ( 
.A1(n_3293),
.A2(n_3080),
.B(n_3046),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3316),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3294),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3324),
.Y(n_3469)
);

BUFx4f_ASAP7_75t_SL g3470 ( 
.A(n_3302),
.Y(n_3470)
);

BUFx2_ASAP7_75t_L g3471 ( 
.A(n_3344),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3304),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3333),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3307),
.Y(n_3474)
);

CKINVDCx20_ASAP7_75t_R g3475 ( 
.A(n_3318),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3355),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_3408),
.Y(n_3477)
);

BUFx2_ASAP7_75t_L g3478 ( 
.A(n_3425),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3396),
.B(n_3257),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3343),
.Y(n_3480)
);

BUFx2_ASAP7_75t_SL g3481 ( 
.A(n_3375),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3346),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3319),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3322),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3360),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3403),
.B(n_3236),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3389),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3401),
.B(n_3238),
.Y(n_3488)
);

BUFx2_ASAP7_75t_L g3489 ( 
.A(n_3425),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3323),
.Y(n_3490)
);

INVxp67_ASAP7_75t_L g3491 ( 
.A(n_3338),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3328),
.Y(n_3492)
);

OAI33xp33_ASAP7_75t_L g3493 ( 
.A1(n_3450),
.A2(n_3278),
.A3(n_3272),
.B1(n_3221),
.B2(n_3203),
.B3(n_3135),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3331),
.Y(n_3494)
);

BUFx3_ASAP7_75t_L g3495 ( 
.A(n_3347),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3374),
.B(n_3267),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3332),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3334),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3361),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3335),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3336),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3341),
.Y(n_3502)
);

HB1xp67_ASAP7_75t_L g3503 ( 
.A(n_3398),
.Y(n_3503)
);

BUFx2_ASAP7_75t_L g3504 ( 
.A(n_3425),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3366),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3371),
.Y(n_3506)
);

BUFx2_ASAP7_75t_L g3507 ( 
.A(n_3425),
.Y(n_3507)
);

AND2x4_ASAP7_75t_L g3508 ( 
.A(n_3296),
.B(n_3406),
.Y(n_3508)
);

OA21x2_ASAP7_75t_L g3509 ( 
.A1(n_3310),
.A2(n_3210),
.B(n_3200),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3430),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_L g3511 ( 
.A1(n_3368),
.A2(n_3171),
.B1(n_3215),
.B2(n_3212),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3453),
.Y(n_3512)
);

AOI21x1_ASAP7_75t_L g3513 ( 
.A1(n_3314),
.A2(n_3156),
.B(n_3199),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3377),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3373),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3298),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3380),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3412),
.Y(n_3518)
);

OA21x2_ASAP7_75t_L g3519 ( 
.A1(n_3327),
.A2(n_3220),
.B(n_3211),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3418),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3426),
.B(n_3188),
.Y(n_3521)
);

BUFx2_ASAP7_75t_L g3522 ( 
.A(n_3315),
.Y(n_3522)
);

OAI21x1_ASAP7_75t_L g3523 ( 
.A1(n_3306),
.A2(n_3110),
.B(n_3226),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3431),
.B(n_3276),
.Y(n_3524)
);

INVx1_ASAP7_75t_SL g3525 ( 
.A(n_3359),
.Y(n_3525)
);

OR2x2_ASAP7_75t_L g3526 ( 
.A(n_3410),
.B(n_3158),
.Y(n_3526)
);

INVx6_ASAP7_75t_L g3527 ( 
.A(n_3390),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3448),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3457),
.Y(n_3529)
);

OAI21x1_ASAP7_75t_L g3530 ( 
.A1(n_3303),
.A2(n_3247),
.B(n_3213),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3330),
.Y(n_3531)
);

BUFx2_ASAP7_75t_L g3532 ( 
.A(n_3315),
.Y(n_3532)
);

HB1xp67_ASAP7_75t_L g3533 ( 
.A(n_3397),
.Y(n_3533)
);

OAI21xp33_ASAP7_75t_SL g3534 ( 
.A1(n_3409),
.A2(n_3190),
.B(n_3233),
.Y(n_3534)
);

CKINVDCx20_ASAP7_75t_R g3535 ( 
.A(n_3414),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3383),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3385),
.Y(n_3537)
);

INVx4_ASAP7_75t_SL g3538 ( 
.A(n_3364),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3391),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3391),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3387),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3351),
.Y(n_3542)
);

HB1xp67_ASAP7_75t_L g3543 ( 
.A(n_3439),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_3405),
.B(n_3249),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3379),
.Y(n_3545)
);

INVx4_ASAP7_75t_L g3546 ( 
.A(n_3342),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3399),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3301),
.B(n_3282),
.Y(n_3548)
);

AND2x4_ASAP7_75t_L g3549 ( 
.A(n_3447),
.B(n_3137),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3432),
.Y(n_3550)
);

HB1xp67_ASAP7_75t_L g3551 ( 
.A(n_3445),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3372),
.Y(n_3552)
);

HB1xp67_ASAP7_75t_L g3553 ( 
.A(n_3451),
.Y(n_3553)
);

HB1xp67_ASAP7_75t_L g3554 ( 
.A(n_3326),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3295),
.A2(n_3254),
.B1(n_3285),
.B2(n_3281),
.Y(n_3555)
);

AOI22xp33_ASAP7_75t_L g3556 ( 
.A1(n_3309),
.A2(n_3281),
.B1(n_3286),
.B2(n_3285),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3382),
.Y(n_3557)
);

HB1xp67_ASAP7_75t_L g3558 ( 
.A(n_3477),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3471),
.B(n_3348),
.Y(n_3559)
);

AO31x2_ASAP7_75t_L g3560 ( 
.A1(n_3522),
.A2(n_3428),
.A3(n_3435),
.B(n_3362),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_R g3561 ( 
.A(n_3535),
.B(n_3440),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3487),
.Y(n_3562)
);

AO31x2_ASAP7_75t_L g3563 ( 
.A1(n_3522),
.A2(n_3395),
.A3(n_3340),
.B(n_3321),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3471),
.B(n_3452),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3478),
.B(n_3317),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3503),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3468),
.Y(n_3567)
);

OR2x2_ASAP7_75t_L g3568 ( 
.A(n_3477),
.B(n_3400),
.Y(n_3568)
);

CKINVDCx16_ASAP7_75t_R g3569 ( 
.A(n_3481),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3512),
.Y(n_3570)
);

CKINVDCx16_ASAP7_75t_R g3571 ( 
.A(n_3546),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3532),
.Y(n_3572)
);

XOR2xp5_ASAP7_75t_L g3573 ( 
.A(n_3475),
.B(n_3074),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3542),
.B(n_3356),
.Y(n_3574)
);

BUFx3_ASAP7_75t_L g3575 ( 
.A(n_3495),
.Y(n_3575)
);

CKINVDCx5p33_ASAP7_75t_R g3576 ( 
.A(n_3470),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3472),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3465),
.Y(n_3578)
);

INVxp67_ASAP7_75t_L g3579 ( 
.A(n_3543),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3467),
.Y(n_3580)
);

BUFx2_ASAP7_75t_L g3581 ( 
.A(n_3534),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3474),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3526),
.B(n_3349),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3552),
.B(n_3411),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3493),
.A2(n_3345),
.B1(n_3300),
.B2(n_3350),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3469),
.Y(n_3586)
);

OAI21x1_ASAP7_75t_L g3587 ( 
.A1(n_3466),
.A2(n_3424),
.B(n_3384),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3473),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3554),
.B(n_3458),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3476),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3533),
.B(n_3420),
.Y(n_3591)
);

CKINVDCx5p33_ASAP7_75t_R g3592 ( 
.A(n_3525),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3488),
.B(n_3444),
.Y(n_3593)
);

CKINVDCx16_ASAP7_75t_R g3594 ( 
.A(n_3479),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3524),
.B(n_3172),
.Y(n_3595)
);

CKINVDCx20_ASAP7_75t_R g3596 ( 
.A(n_3551),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_3527),
.Y(n_3597)
);

BUFx6f_ASAP7_75t_L g3598 ( 
.A(n_3527),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3480),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3482),
.Y(n_3600)
);

AO31x2_ASAP7_75t_L g3601 ( 
.A1(n_3489),
.A2(n_3442),
.A3(n_3320),
.B(n_3402),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_3491),
.Y(n_3602)
);

BUFx3_ASAP7_75t_L g3603 ( 
.A(n_3553),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3485),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3483),
.Y(n_3605)
);

HB1xp67_ASAP7_75t_L g3606 ( 
.A(n_3499),
.Y(n_3606)
);

CKINVDCx16_ASAP7_75t_R g3607 ( 
.A(n_3548),
.Y(n_3607)
);

BUFx2_ASAP7_75t_L g3608 ( 
.A(n_3538),
.Y(n_3608)
);

HB1xp67_ASAP7_75t_L g3609 ( 
.A(n_3518),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3520),
.Y(n_3610)
);

OR2x6_ASAP7_75t_L g3611 ( 
.A(n_3544),
.B(n_3422),
.Y(n_3611)
);

INVx6_ASAP7_75t_SL g3612 ( 
.A(n_3508),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3484),
.Y(n_3613)
);

AND2x4_ASAP7_75t_SL g3614 ( 
.A(n_3549),
.B(n_3393),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_3521),
.B(n_3194),
.Y(n_3615)
);

INVx2_ASAP7_75t_SL g3616 ( 
.A(n_3538),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3490),
.Y(n_3617)
);

INVx1_ASAP7_75t_SL g3618 ( 
.A(n_3496),
.Y(n_3618)
);

NOR2xp33_ASAP7_75t_L g3619 ( 
.A(n_3550),
.B(n_3081),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3492),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3536),
.Y(n_3621)
);

HB1xp67_ASAP7_75t_L g3622 ( 
.A(n_3505),
.Y(n_3622)
);

BUFx4f_ASAP7_75t_SL g3623 ( 
.A(n_3541),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3547),
.B(n_3218),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3622),
.Y(n_3625)
);

NAND2x1p5_ASAP7_75t_L g3626 ( 
.A(n_3575),
.B(n_3071),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3559),
.B(n_3564),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3599),
.Y(n_3628)
);

INVxp67_ASAP7_75t_SL g3629 ( 
.A(n_3558),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3609),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3607),
.B(n_3504),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3572),
.B(n_3507),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3615),
.B(n_3507),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_3606),
.B(n_3486),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3600),
.Y(n_3635)
);

HB1xp67_ASAP7_75t_L g3636 ( 
.A(n_3596),
.Y(n_3636)
);

HB1xp67_ASAP7_75t_L g3637 ( 
.A(n_3603),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3618),
.B(n_3545),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3574),
.B(n_3531),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3562),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3566),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3610),
.Y(n_3642)
);

HB1xp67_ASAP7_75t_L g3643 ( 
.A(n_3579),
.Y(n_3643)
);

CKINVDCx20_ASAP7_75t_R g3644 ( 
.A(n_3569),
.Y(n_3644)
);

HB1xp67_ASAP7_75t_L g3645 ( 
.A(n_3611),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3571),
.B(n_3557),
.Y(n_3646)
);

BUFx3_ASAP7_75t_L g3647 ( 
.A(n_3576),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3578),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3580),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3604),
.Y(n_3650)
);

OR2x6_ASAP7_75t_L g3651 ( 
.A(n_3608),
.B(n_3427),
.Y(n_3651)
);

OR2x2_ASAP7_75t_L g3652 ( 
.A(n_3570),
.B(n_3502),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3567),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3577),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3582),
.Y(n_3655)
);

CKINVDCx20_ASAP7_75t_R g3656 ( 
.A(n_3561),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3586),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3590),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3595),
.B(n_3528),
.Y(n_3659)
);

HB1xp67_ASAP7_75t_L g3660 ( 
.A(n_3568),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3605),
.B(n_3539),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3588),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3621),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3613),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3617),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3620),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3583),
.Y(n_3667)
);

OAI221xp5_ASAP7_75t_L g3668 ( 
.A1(n_3585),
.A2(n_3555),
.B1(n_3511),
.B2(n_3556),
.C(n_3299),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_3584),
.B(n_3506),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3589),
.B(n_3540),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_3612),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3565),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3581),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3591),
.Y(n_3674)
);

CKINVDCx20_ASAP7_75t_R g3675 ( 
.A(n_3594),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3593),
.B(n_3510),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3614),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3623),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3560),
.B(n_3515),
.Y(n_3679)
);

HB1xp67_ASAP7_75t_L g3680 ( 
.A(n_3592),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3587),
.Y(n_3681)
);

INVx3_ASAP7_75t_L g3682 ( 
.A(n_3616),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3601),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3625),
.B(n_3667),
.Y(n_3684)
);

HB1xp67_ASAP7_75t_L g3685 ( 
.A(n_3629),
.Y(n_3685)
);

OR2x2_ASAP7_75t_L g3686 ( 
.A(n_3667),
.B(n_3514),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3630),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3625),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3658),
.Y(n_3689)
);

INVxp67_ASAP7_75t_L g3690 ( 
.A(n_3637),
.Y(n_3690)
);

BUFx2_ASAP7_75t_L g3691 ( 
.A(n_3675),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_SL g3692 ( 
.A(n_3644),
.B(n_3597),
.Y(n_3692)
);

OR2x2_ASAP7_75t_L g3693 ( 
.A(n_3639),
.B(n_3517),
.Y(n_3693)
);

OR2x2_ASAP7_75t_L g3694 ( 
.A(n_3669),
.B(n_3494),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3661),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3664),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3640),
.B(n_3601),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3658),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3665),
.Y(n_3699)
);

NAND4xp25_ASAP7_75t_L g3700 ( 
.A(n_3668),
.B(n_3624),
.C(n_3394),
.D(n_3460),
.Y(n_3700)
);

HB1xp67_ASAP7_75t_L g3701 ( 
.A(n_3643),
.Y(n_3701)
);

BUFx3_ASAP7_75t_L g3702 ( 
.A(n_3656),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3645),
.B(n_3619),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3631),
.B(n_3598),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3641),
.B(n_3563),
.Y(n_3705)
);

BUFx6f_ASAP7_75t_L g3706 ( 
.A(n_3647),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3666),
.Y(n_3707)
);

BUFx4f_ASAP7_75t_L g3708 ( 
.A(n_3651),
.Y(n_3708)
);

OAI22xp33_ASAP7_75t_L g3709 ( 
.A1(n_3673),
.A2(n_3602),
.B1(n_3519),
.B2(n_3509),
.Y(n_3709)
);

OAI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3651),
.A2(n_3519),
.B1(n_3509),
.B2(n_3240),
.Y(n_3710)
);

INVx4_ASAP7_75t_L g3711 ( 
.A(n_3626),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3653),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3662),
.Y(n_3713)
);

BUFx2_ASAP7_75t_L g3714 ( 
.A(n_3636),
.Y(n_3714)
);

AOI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3683),
.A2(n_3436),
.B1(n_3308),
.B2(n_3370),
.C(n_3497),
.Y(n_3715)
);

INVx5_ASAP7_75t_L g3716 ( 
.A(n_3671),
.Y(n_3716)
);

NAND3xp33_ASAP7_75t_L g3717 ( 
.A(n_3681),
.B(n_3679),
.C(n_3680),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3654),
.Y(n_3718)
);

HB1xp67_ASAP7_75t_L g3719 ( 
.A(n_3660),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3642),
.Y(n_3720)
);

BUFx2_ASAP7_75t_L g3721 ( 
.A(n_3682),
.Y(n_3721)
);

OA21x2_ASAP7_75t_L g3722 ( 
.A1(n_3681),
.A2(n_3530),
.B(n_3516),
.Y(n_3722)
);

A2O1A1Ixp33_ASAP7_75t_L g3723 ( 
.A1(n_3671),
.A2(n_3456),
.B(n_3461),
.C(n_3438),
.Y(n_3723)
);

BUFx3_ASAP7_75t_L g3724 ( 
.A(n_3678),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_3646),
.Y(n_3725)
);

AOI22xp33_ASAP7_75t_L g3726 ( 
.A1(n_3674),
.A2(n_3268),
.B1(n_3097),
.B2(n_3258),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3655),
.Y(n_3727)
);

INVx3_ASAP7_75t_L g3728 ( 
.A(n_3677),
.Y(n_3728)
);

AOI22xp33_ASAP7_75t_L g3729 ( 
.A1(n_3672),
.A2(n_3255),
.B1(n_3170),
.B2(n_3166),
.Y(n_3729)
);

A2O1A1Ixp33_ASAP7_75t_L g3730 ( 
.A1(n_3634),
.A2(n_3358),
.B(n_3354),
.C(n_3388),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3648),
.Y(n_3731)
);

INVxp67_ASAP7_75t_SL g3732 ( 
.A(n_3649),
.Y(n_3732)
);

A2O1A1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_3627),
.A2(n_3633),
.B(n_3632),
.C(n_3676),
.Y(n_3733)
);

AOI21xp5_ASAP7_75t_SL g3734 ( 
.A1(n_3711),
.A2(n_3573),
.B(n_3455),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3708),
.A2(n_3670),
.B(n_3638),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3714),
.Y(n_3736)
);

HB1xp67_ASAP7_75t_L g3737 ( 
.A(n_3719),
.Y(n_3737)
);

BUFx2_ASAP7_75t_L g3738 ( 
.A(n_3721),
.Y(n_3738)
);

INVx4_ASAP7_75t_L g3739 ( 
.A(n_3706),
.Y(n_3739)
);

NAND2x1p5_ASAP7_75t_L g3740 ( 
.A(n_3716),
.B(n_3071),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3701),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_SL g3742 ( 
.A(n_3692),
.B(n_3417),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3685),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3694),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3695),
.B(n_3563),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3720),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3684),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3731),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3703),
.B(n_3659),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3706),
.Y(n_3750)
);

CKINVDCx5p33_ASAP7_75t_R g3751 ( 
.A(n_3702),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3690),
.Y(n_3752)
);

OR2x2_ASAP7_75t_L g3753 ( 
.A(n_3693),
.B(n_3652),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3686),
.Y(n_3754)
);

INVx3_ASAP7_75t_L g3755 ( 
.A(n_3716),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3700),
.A2(n_3245),
.B1(n_3152),
.B2(n_3464),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3716),
.B(n_3628),
.Y(n_3757)
);

HB1xp67_ASAP7_75t_L g3758 ( 
.A(n_3687),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_SL g3759 ( 
.A1(n_3730),
.A2(n_3421),
.B(n_3297),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3704),
.B(n_3628),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3728),
.B(n_3635),
.Y(n_3761)
);

INVx2_ASAP7_75t_SL g3762 ( 
.A(n_3724),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3696),
.Y(n_3763)
);

AOI221xp5_ASAP7_75t_L g3764 ( 
.A1(n_3697),
.A2(n_3650),
.B1(n_3498),
.B2(n_3501),
.C(n_3500),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3712),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3691),
.B(n_3657),
.Y(n_3766)
);

AOI222xp33_ASAP7_75t_L g3767 ( 
.A1(n_3725),
.A2(n_3459),
.B1(n_3404),
.B2(n_3423),
.C1(n_3446),
.C2(n_3369),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3733),
.B(n_3663),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3689),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3698),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3718),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3699),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3688),
.B(n_3705),
.Y(n_3773)
);

OAI33xp33_ASAP7_75t_L g3774 ( 
.A1(n_3709),
.A2(n_3416),
.A3(n_3352),
.B1(n_3529),
.B2(n_3353),
.B3(n_3537),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3707),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3727),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3732),
.B(n_3441),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3713),
.B(n_3441),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3722),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3726),
.B(n_3365),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3722),
.Y(n_3781)
);

INVx5_ASAP7_75t_SL g3782 ( 
.A(n_3729),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3736),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3737),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3743),
.B(n_3741),
.Y(n_3785)
);

OR2x2_ASAP7_75t_L g3786 ( 
.A(n_3752),
.B(n_3717),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3747),
.B(n_3710),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3766),
.Y(n_3788)
);

AND2x4_ASAP7_75t_L g3789 ( 
.A(n_3762),
.B(n_3723),
.Y(n_3789)
);

OR2x2_ASAP7_75t_L g3790 ( 
.A(n_3754),
.B(n_3419),
.Y(n_3790)
);

OR2x2_ASAP7_75t_L g3791 ( 
.A(n_3744),
.B(n_3745),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3782),
.B(n_3715),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3764),
.B(n_3523),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3753),
.B(n_3454),
.Y(n_3794)
);

BUFx2_ASAP7_75t_L g3795 ( 
.A(n_3739),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3738),
.B(n_3513),
.Y(n_3796)
);

OR2x2_ASAP7_75t_L g3797 ( 
.A(n_3763),
.B(n_3454),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3768),
.B(n_3378),
.Y(n_3798)
);

AND2x4_ASAP7_75t_L g3799 ( 
.A(n_3739),
.B(n_3096),
.Y(n_3799)
);

AND2x4_ASAP7_75t_L g3800 ( 
.A(n_3750),
.B(n_3755),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3763),
.B(n_3772),
.Y(n_3801)
);

CKINVDCx16_ASAP7_75t_R g3802 ( 
.A(n_3742),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3749),
.B(n_3386),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3772),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_3751),
.B(n_3089),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3776),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3761),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3776),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3760),
.B(n_3392),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3765),
.B(n_3407),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3734),
.B(n_3735),
.Y(n_3811)
);

BUFx2_ASAP7_75t_L g3812 ( 
.A(n_3777),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3775),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3800),
.B(n_3757),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3800),
.B(n_3758),
.Y(n_3815)
);

OR2x2_ASAP7_75t_L g3816 ( 
.A(n_3784),
.B(n_3773),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3795),
.B(n_3756),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3785),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3792),
.A2(n_3774),
.B1(n_3767),
.B2(n_3780),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3812),
.B(n_3778),
.Y(n_3820)
);

OAI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3811),
.A2(n_3759),
.B(n_3781),
.Y(n_3821)
);

OR2x2_ASAP7_75t_L g3822 ( 
.A(n_3783),
.B(n_3775),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3793),
.B(n_3771),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3801),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3788),
.B(n_3746),
.Y(n_3825)
);

OAI31xp33_ASAP7_75t_L g3826 ( 
.A1(n_3789),
.A2(n_3781),
.A3(n_3779),
.B(n_3740),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3794),
.B(n_3748),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3802),
.B(n_3769),
.Y(n_3828)
);

AND2x4_ASAP7_75t_L g3829 ( 
.A(n_3799),
.B(n_3770),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3798),
.B(n_3789),
.Y(n_3830)
);

INVxp67_ASAP7_75t_L g3831 ( 
.A(n_3805),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3807),
.Y(n_3832)
);

NOR2x1_ASAP7_75t_L g3833 ( 
.A(n_3799),
.B(n_3415),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3804),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3813),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3813),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3786),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3818),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3817),
.B(n_3803),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3815),
.B(n_3809),
.Y(n_3840)
);

INVx1_ASAP7_75t_SL g3841 ( 
.A(n_3828),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3837),
.B(n_3791),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3816),
.Y(n_3843)
);

INVx1_ASAP7_75t_SL g3844 ( 
.A(n_3814),
.Y(n_3844)
);

AO21x2_ASAP7_75t_L g3845 ( 
.A1(n_3821),
.A2(n_3808),
.B(n_3806),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3830),
.B(n_3787),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3820),
.B(n_3796),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3825),
.Y(n_3848)
);

OAI211xp5_ASAP7_75t_SL g3849 ( 
.A1(n_3826),
.A2(n_3790),
.B(n_3810),
.C(n_3797),
.Y(n_3849)
);

AND2x4_ASAP7_75t_L g3850 ( 
.A(n_3831),
.B(n_3196),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3832),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3819),
.B(n_3193),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3822),
.Y(n_3853)
);

CKINVDCx16_ASAP7_75t_R g3854 ( 
.A(n_3833),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3827),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3824),
.Y(n_3856)
);

INVx4_ASAP7_75t_L g3857 ( 
.A(n_3829),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3834),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3823),
.B(n_3197),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3829),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3834),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3835),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3835),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3836),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_3857),
.B(n_613),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3854),
.B(n_614),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3846),
.B(n_3227),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3842),
.B(n_615),
.Y(n_3868)
);

NOR2xp67_ASAP7_75t_L g3869 ( 
.A(n_3857),
.B(n_615),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3841),
.B(n_616),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3851),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3860),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3839),
.B(n_3847),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3844),
.B(n_616),
.Y(n_3874)
);

OR2x2_ASAP7_75t_L g3875 ( 
.A(n_3843),
.B(n_616),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3840),
.B(n_3376),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3840),
.B(n_3463),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3855),
.B(n_617),
.Y(n_3878)
);

AOI22xp33_ASAP7_75t_L g3879 ( 
.A1(n_3848),
.A2(n_3167),
.B1(n_3367),
.B2(n_3159),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3838),
.Y(n_3880)
);

INVx3_ASAP7_75t_L g3881 ( 
.A(n_3850),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3853),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3850),
.B(n_3413),
.Y(n_3883)
);

BUFx2_ASAP7_75t_L g3884 ( 
.A(n_3856),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3863),
.B(n_3449),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3862),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3859),
.B(n_3852),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3845),
.B(n_3462),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3862),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3864),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3858),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3861),
.B(n_618),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3866),
.A2(n_3849),
.B(n_3381),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3870),
.Y(n_3894)
);

OAI321xp33_ASAP7_75t_L g3895 ( 
.A1(n_3880),
.A2(n_3162),
.A3(n_3078),
.B1(n_3075),
.B2(n_3085),
.C(n_3077),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3874),
.B(n_618),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3868),
.B(n_619),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3869),
.Y(n_3898)
);

INVx3_ASAP7_75t_L g3899 ( 
.A(n_3881),
.Y(n_3899)
);

INVx2_ASAP7_75t_SL g3900 ( 
.A(n_3881),
.Y(n_3900)
);

OAI221xp5_ASAP7_75t_L g3901 ( 
.A1(n_3871),
.A2(n_3102),
.B1(n_3120),
.B2(n_3093),
.C(n_3091),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3873),
.B(n_3877),
.Y(n_3902)
);

XOR2xp5_ASAP7_75t_L g3903 ( 
.A(n_3875),
.B(n_620),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3867),
.B(n_621),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3888),
.B(n_622),
.Y(n_3905)
);

HB1xp67_ASAP7_75t_L g3906 ( 
.A(n_3878),
.Y(n_3906)
);

OAI32xp33_ASAP7_75t_L g3907 ( 
.A1(n_3891),
.A2(n_3129),
.A3(n_3125),
.B1(n_3112),
.B2(n_3119),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3887),
.B(n_623),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3892),
.A2(n_3433),
.B(n_3429),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3883),
.B(n_624),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3876),
.Y(n_3911)
);

OAI221xp5_ASAP7_75t_L g3912 ( 
.A1(n_3879),
.A2(n_3884),
.B1(n_3890),
.B2(n_3886),
.C(n_3889),
.Y(n_3912)
);

OAI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3885),
.A2(n_3437),
.B(n_3434),
.Y(n_3913)
);

AOI21xp33_ASAP7_75t_L g3914 ( 
.A1(n_3880),
.A2(n_625),
.B(n_626),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3873),
.B(n_625),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3873),
.B(n_626),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3866),
.A2(n_3443),
.B(n_3325),
.Y(n_3917)
);

INVxp33_ASAP7_75t_L g3918 ( 
.A(n_3865),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3873),
.B(n_627),
.Y(n_3919)
);

AOI221xp5_ASAP7_75t_L g3920 ( 
.A1(n_3882),
.A2(n_3202),
.B1(n_3162),
.B2(n_3151),
.C(n_3143),
.Y(n_3920)
);

INVxp67_ASAP7_75t_L g3921 ( 
.A(n_3865),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3872),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3872),
.Y(n_3923)
);

AOI311xp33_ASAP7_75t_L g3924 ( 
.A1(n_3882),
.A2(n_629),
.A3(n_627),
.B(n_628),
.C(n_630),
.Y(n_3924)
);

OAI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3882),
.A2(n_3339),
.B(n_3329),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3923),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3922),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3900),
.B(n_629),
.Y(n_3928)
);

NAND2x1p5_ASAP7_75t_L g3929 ( 
.A(n_3899),
.B(n_3051),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3915),
.B(n_629),
.Y(n_3930)
);

NOR2xp67_ASAP7_75t_SL g3931 ( 
.A(n_3899),
.B(n_3896),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3908),
.B(n_3902),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3911),
.Y(n_3933)
);

NAND2xp33_ASAP7_75t_SL g3934 ( 
.A(n_3918),
.B(n_3051),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3904),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3910),
.B(n_630),
.Y(n_3936)
);

OR2x2_ASAP7_75t_L g3937 ( 
.A(n_3916),
.B(n_630),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3919),
.Y(n_3938)
);

NAND2x1p5_ASAP7_75t_L g3939 ( 
.A(n_3897),
.B(n_3085),
.Y(n_3939)
);

OR2x2_ASAP7_75t_L g3940 ( 
.A(n_3905),
.B(n_631),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3898),
.B(n_632),
.Y(n_3941)
);

NAND3xp33_ASAP7_75t_L g3942 ( 
.A(n_3914),
.B(n_632),
.C(n_633),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3903),
.B(n_633),
.Y(n_3943)
);

INVxp33_ASAP7_75t_L g3944 ( 
.A(n_3906),
.Y(n_3944)
);

NAND2x1_ASAP7_75t_L g3945 ( 
.A(n_3894),
.B(n_3087),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3917),
.B(n_634),
.Y(n_3946)
);

NOR2x1_ASAP7_75t_L g3947 ( 
.A(n_3912),
.B(n_636),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3893),
.B(n_636),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3921),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3924),
.B(n_3090),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3913),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3909),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3926),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3933),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3926),
.Y(n_3955)
);

NAND2xp33_ASAP7_75t_SL g3956 ( 
.A(n_3948),
.B(n_3931),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3930),
.B(n_3920),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3932),
.B(n_3936),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3928),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3943),
.B(n_3907),
.Y(n_3960)
);

OAI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_3947),
.A2(n_3895),
.B(n_3925),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3929),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3950),
.Y(n_3963)
);

INVx1_ASAP7_75t_SL g3964 ( 
.A(n_3934),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3941),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3927),
.B(n_3901),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3937),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3939),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3951),
.B(n_3952),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_SL g3970 ( 
.A(n_3946),
.B(n_3092),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3940),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_L g3972 ( 
.A(n_3942),
.B(n_637),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3949),
.Y(n_3973)
);

OAI21xp33_ASAP7_75t_L g3974 ( 
.A1(n_3944),
.A2(n_637),
.B(n_638),
.Y(n_3974)
);

INVxp67_ASAP7_75t_L g3975 ( 
.A(n_3938),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3945),
.Y(n_3976)
);

AOI221x1_ASAP7_75t_L g3977 ( 
.A1(n_3935),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.C(n_643),
.Y(n_3977)
);

INVx1_ASAP7_75t_SL g3978 ( 
.A(n_3926),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3926),
.B(n_642),
.Y(n_3979)
);

NAND4xp25_ASAP7_75t_L g3980 ( 
.A(n_3958),
.B(n_645),
.C(n_643),
.D(n_644),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3954),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3963),
.B(n_3092),
.Y(n_3982)
);

NOR4xp25_ASAP7_75t_L g3983 ( 
.A(n_3978),
.B(n_645),
.C(n_643),
.D(n_644),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3976),
.Y(n_3984)
);

INVx1_ASAP7_75t_SL g3985 ( 
.A(n_3964),
.Y(n_3985)
);

INVxp67_ASAP7_75t_L g3986 ( 
.A(n_3972),
.Y(n_3986)
);

A2O1A1Ixp33_ASAP7_75t_SL g3987 ( 
.A1(n_3973),
.A2(n_648),
.B(n_646),
.C(n_647),
.Y(n_3987)
);

NOR3xp33_ASAP7_75t_L g3988 ( 
.A(n_3974),
.B(n_646),
.C(n_647),
.Y(n_3988)
);

NAND3xp33_ASAP7_75t_L g3989 ( 
.A(n_3969),
.B(n_648),
.C(n_649),
.Y(n_3989)
);

NOR3xp33_ASAP7_75t_L g3990 ( 
.A(n_3953),
.B(n_648),
.C(n_649),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3965),
.B(n_650),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3979),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3955),
.B(n_650),
.Y(n_3993)
);

NAND4xp25_ASAP7_75t_L g3994 ( 
.A(n_3960),
.B(n_653),
.C(n_651),
.D(n_652),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3957),
.Y(n_3995)
);

OR2x2_ASAP7_75t_L g3996 ( 
.A(n_3966),
.B(n_656),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_L g3997 ( 
.A(n_3962),
.B(n_657),
.Y(n_3997)
);

NAND4xp75_ASAP7_75t_L g3998 ( 
.A(n_3977),
.B(n_660),
.C(n_658),
.D(n_659),
.Y(n_3998)
);

NAND4xp25_ASAP7_75t_L g3999 ( 
.A(n_3956),
.B(n_660),
.C(n_658),
.D(n_659),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3967),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_L g4001 ( 
.A(n_3968),
.B(n_660),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3971),
.Y(n_4002)
);

OAI221xp5_ASAP7_75t_SL g4003 ( 
.A1(n_3985),
.A2(n_3984),
.B1(n_3981),
.B2(n_3996),
.C(n_3983),
.Y(n_4003)
);

OAI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3989),
.A2(n_3961),
.B(n_3975),
.Y(n_4004)
);

OAI221xp5_ASAP7_75t_L g4005 ( 
.A1(n_3988),
.A2(n_3970),
.B1(n_3959),
.B2(n_663),
.C(n_661),
.Y(n_4005)
);

AOI211xp5_ASAP7_75t_SL g4006 ( 
.A1(n_4001),
.A2(n_663),
.B(n_661),
.C(n_662),
.Y(n_4006)
);

OAI221xp5_ASAP7_75t_L g4007 ( 
.A1(n_3999),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.C(n_665),
.Y(n_4007)
);

OAI211xp5_ASAP7_75t_SL g4008 ( 
.A1(n_3995),
.A2(n_667),
.B(n_665),
.C(n_666),
.Y(n_4008)
);

OAI321xp33_ASAP7_75t_L g4009 ( 
.A1(n_4000),
.A2(n_669),
.A3(n_671),
.B1(n_666),
.B2(n_668),
.C(n_670),
.Y(n_4009)
);

AOI222xp33_ASAP7_75t_L g4010 ( 
.A1(n_3982),
.A2(n_3106),
.B1(n_3217),
.B2(n_3337),
.C1(n_670),
.C2(n_672),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3991),
.Y(n_4011)
);

OAI21xp33_ASAP7_75t_L g4012 ( 
.A1(n_3994),
.A2(n_3363),
.B(n_3357),
.Y(n_4012)
);

AND2x4_ASAP7_75t_L g4013 ( 
.A(n_4002),
.B(n_668),
.Y(n_4013)
);

AOI221xp5_ASAP7_75t_L g4014 ( 
.A1(n_3980),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.C(n_674),
.Y(n_4014)
);

O2A1O1Ixp33_ASAP7_75t_L g4015 ( 
.A1(n_3990),
.A2(n_673),
.B(n_674),
.C(n_714),
.Y(n_4015)
);

OAI211xp5_ASAP7_75t_L g4016 ( 
.A1(n_3997),
.A2(n_717),
.B(n_715),
.C(n_716),
.Y(n_4016)
);

AOI21xp33_ASAP7_75t_L g4017 ( 
.A1(n_3993),
.A2(n_719),
.B(n_721),
.Y(n_4017)
);

AOI221xp5_ASAP7_75t_L g4018 ( 
.A1(n_3986),
.A2(n_3201),
.B1(n_3223),
.B2(n_3228),
.C(n_3222),
.Y(n_4018)
);

AOI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3998),
.A2(n_3049),
.B1(n_3305),
.B2(n_3311),
.Y(n_4019)
);

AOI221xp5_ASAP7_75t_L g4020 ( 
.A1(n_3992),
.A2(n_3201),
.B1(n_3223),
.B2(n_3228),
.C(n_3222),
.Y(n_4020)
);

AOI21xp33_ASAP7_75t_L g4021 ( 
.A1(n_3987),
.A2(n_723),
.B(n_724),
.Y(n_4021)
);

OAI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3984),
.A2(n_3230),
.B1(n_3235),
.B2(n_3313),
.Y(n_4022)
);

OAI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_4003),
.A2(n_3313),
.B1(n_3230),
.B2(n_3235),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_4013),
.B(n_3049),
.Y(n_4024)
);

OAI211xp5_ASAP7_75t_L g4025 ( 
.A1(n_4014),
.A2(n_729),
.B(n_727),
.C(n_728),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_4013),
.B(n_728),
.Y(n_4026)
);

AOI21xp33_ASAP7_75t_L g4027 ( 
.A1(n_4015),
.A2(n_4007),
.B(n_4016),
.Y(n_4027)
);

AOI211xp5_ASAP7_75t_L g4028 ( 
.A1(n_4021),
.A2(n_4017),
.B(n_4005),
.C(n_4008),
.Y(n_4028)
);

OAI22xp33_ASAP7_75t_L g4029 ( 
.A1(n_4006),
.A2(n_732),
.B1(n_730),
.B2(n_731),
.Y(n_4029)
);

A2O1A1Ixp33_ASAP7_75t_SL g4030 ( 
.A1(n_4004),
.A2(n_733),
.B(n_731),
.C(n_732),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_4011),
.Y(n_4031)
);

AOI221xp5_ASAP7_75t_L g4032 ( 
.A1(n_4009),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.C(n_736),
.Y(n_4032)
);

OAI31xp33_ASAP7_75t_L g4033 ( 
.A1(n_4025),
.A2(n_4012),
.A3(n_4010),
.B(n_4022),
.Y(n_4033)
);

AOI321xp33_ASAP7_75t_L g4034 ( 
.A1(n_4028),
.A2(n_4019),
.A3(n_4020),
.B1(n_4018),
.B2(n_739),
.C(n_741),
.Y(n_4034)
);

AND2x4_ASAP7_75t_L g4035 ( 
.A(n_4031),
.B(n_737),
.Y(n_4035)
);

AOI21xp33_ASAP7_75t_L g4036 ( 
.A1(n_4030),
.A2(n_738),
.B(n_739),
.Y(n_4036)
);

AOI311xp33_ASAP7_75t_L g4037 ( 
.A1(n_4027),
.A2(n_742),
.A3(n_740),
.B(n_741),
.C(n_743),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_4026),
.B(n_742),
.Y(n_4038)
);

AOI21xp33_ASAP7_75t_L g4039 ( 
.A1(n_4029),
.A2(n_743),
.B(n_744),
.Y(n_4039)
);

OAI22xp5_ASAP7_75t_L g4040 ( 
.A1(n_4023),
.A2(n_747),
.B1(n_745),
.B2(n_746),
.Y(n_4040)
);

NOR3xp33_ASAP7_75t_L g4041 ( 
.A(n_4032),
.B(n_747),
.C(n_748),
.Y(n_4041)
);

OAI22xp33_ASAP7_75t_SL g4042 ( 
.A1(n_4024),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.Y(n_4042)
);

NAND4xp25_ASAP7_75t_L g4043 ( 
.A(n_4034),
.B(n_754),
.C(n_752),
.D(n_753),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_4035),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_4035),
.Y(n_4045)
);

OAI211xp5_ASAP7_75t_L g4046 ( 
.A1(n_4039),
.A2(n_760),
.B(n_757),
.C(n_759),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_4038),
.B(n_4037),
.Y(n_4047)
);

AOI221xp5_ASAP7_75t_L g4048 ( 
.A1(n_4036),
.A2(n_763),
.B1(n_761),
.B2(n_762),
.C(n_764),
.Y(n_4048)
);

NAND4xp25_ASAP7_75t_L g4049 ( 
.A(n_4033),
.B(n_763),
.C(n_761),
.D(n_762),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_4040),
.Y(n_4050)
);

CKINVDCx5p33_ASAP7_75t_R g4051 ( 
.A(n_4042),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_4041),
.B(n_764),
.Y(n_4052)
);

CKINVDCx5p33_ASAP7_75t_R g4053 ( 
.A(n_4051),
.Y(n_4053)
);

HB1xp67_ASAP7_75t_L g4054 ( 
.A(n_4047),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_4044),
.Y(n_4055)
);

CKINVDCx5p33_ASAP7_75t_R g4056 ( 
.A(n_4045),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_4054),
.Y(n_4057)
);

XNOR2xp5_ASAP7_75t_L g4058 ( 
.A(n_4056),
.B(n_4043),
.Y(n_4058)
);

OA22x2_ASAP7_75t_L g4059 ( 
.A1(n_4055),
.A2(n_4050),
.B1(n_4052),
.B2(n_4046),
.Y(n_4059)
);

AND3x4_ASAP7_75t_L g4060 ( 
.A(n_4053),
.B(n_4049),
.C(n_4048),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_4054),
.Y(n_4061)
);

XNOR2x1_ASAP7_75t_L g4062 ( 
.A(n_4060),
.B(n_766),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_4057),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_4061),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4062),
.Y(n_4065)
);

OAI21xp5_ASAP7_75t_L g4066 ( 
.A1(n_4065),
.A2(n_4064),
.B(n_4063),
.Y(n_4066)
);

OAI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_4066),
.A2(n_4058),
.B(n_4059),
.Y(n_4067)
);

INVxp33_ASAP7_75t_L g4068 ( 
.A(n_4067),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_4068),
.Y(n_4069)
);

AOI222xp33_ASAP7_75t_L g4070 ( 
.A1(n_4069),
.A2(n_771),
.B1(n_773),
.B2(n_769),
.C1(n_770),
.C2(n_772),
.Y(n_4070)
);

INVxp67_ASAP7_75t_L g4071 ( 
.A(n_4070),
.Y(n_4071)
);

AOI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_4071),
.A2(n_777),
.B1(n_775),
.B2(n_776),
.Y(n_4072)
);

AOI211xp5_ASAP7_75t_L g4073 ( 
.A1(n_4072),
.A2(n_781),
.B(n_779),
.C(n_780),
.Y(n_4073)
);


endmodule