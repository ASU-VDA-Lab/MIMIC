module fake_jpeg_3169_n_173 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_34),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_7),
.B(n_1),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_0),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_80),
.B1(n_60),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_58),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_57),
.B1(n_56),
.B2(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_57),
.B1(n_45),
.B2(n_53),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_66),
.B(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_97),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_71),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_27),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_52),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_88),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_12),
.C(n_13),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_47),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_20),
.C(n_21),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_47),
.B1(n_3),
.B2(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_117),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_84),
.B(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.C(n_112),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_111),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_6),
.CI(n_9),
.CON(n_121),
.SN(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_9),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_10),
.CI(n_11),
.CON(n_125),
.SN(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_126),
.Y(n_143)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_12),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_13),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_135),
.B1(n_117),
.B2(n_115),
.Y(n_138)
);

CKINVDCx10_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_14),
.Y(n_135)
);

NOR2x1_ASAP7_75t_R g142 ( 
.A(n_136),
.B(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_138),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_22),
.B(n_24),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_124),
.B(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_35),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_153),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_122),
.B1(n_125),
.B2(n_121),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_157),
.B1(n_149),
.B2(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_153),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_150),
.B1(n_144),
.B2(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_141),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_152),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_166),
.A3(n_162),
.B1(n_161),
.B2(n_163),
.C1(n_164),
.C2(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_145),
.B(n_147),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_148),
.C(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_44),
.Y(n_173)
);


endmodule