module fake_netlist_5_1207_n_1778 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1778);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1778;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g161 ( 
.A(n_43),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_47),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_71),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_52),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_30),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_50),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_17),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_48),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_56),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_81),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_98),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_84),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_128),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_29),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_82),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_67),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_34),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_45),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_122),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_32),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_97),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_83),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_99),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_124),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_26),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_20),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_100),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_101),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_92),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_88),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_55),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_144),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_80),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_44),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_113),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_70),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_90),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_142),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_53),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_6),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_15),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_58),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_36),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_55),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_22),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_69),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_52),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_73),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_148),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_42),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_126),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_48),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_64),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_32),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_57),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_141),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_28),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_39),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_91),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_8),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_109),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_61),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_149),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_86),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_76),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_39),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_13),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_159),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_119),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_75),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_79),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_59),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_85),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_15),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_62),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_34),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_49),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_25),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_154),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_49),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_4),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_44),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_22),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_77),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_53),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_27),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_190),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_173),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_255),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_298),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_224),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_168),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_194),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_179),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_181),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_173),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_173),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_0),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_200),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_173),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_215),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_215),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_215),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_215),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_186),
.B(n_0),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_215),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_284),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_180),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_185),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_250),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_166),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_186),
.B(n_2),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_224),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_191),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_196),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_192),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_282),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_207),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_253),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_214),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_162),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_161),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_161),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_178),
.B(n_2),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_164),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_219),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_164),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_170),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_261),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_220),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_163),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_170),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_227),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_222),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_178),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_181),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_175),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_175),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_228),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_232),
.B(n_112),
.Y(n_387)
);

BUFx6f_ASAP7_75t_SL g388 ( 
.A(n_174),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_172),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_182),
.B(n_3),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_176),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_176),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_177),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_177),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_199),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_358),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_330),
.B(n_289),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_289),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_206),
.B(n_199),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_340),
.B(n_322),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_333),
.B(n_174),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_247),
.B(n_206),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_353),
.B(n_226),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_371),
.B(n_174),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_336),
.A2(n_226),
.B(n_184),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_337),
.B(n_233),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_338),
.B(n_221),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_368),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_323),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_325),
.A2(n_169),
.B1(n_318),
.B2(n_302),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_239),
.B1(n_193),
.B2(n_268),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_341),
.A2(n_252),
.B(n_247),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_324),
.B(n_174),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_352),
.B(n_221),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_343),
.B(n_236),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_346),
.B(n_182),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_345),
.A2(n_171),
.B1(n_249),
.B2(n_314),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_348),
.B(n_261),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_184),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_378),
.B(n_212),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_359),
.B(n_189),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_356),
.B(n_189),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_354),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_364),
.A2(n_217),
.B1(n_304),
.B2(n_285),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_183),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_369),
.B(n_370),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_370),
.B(n_195),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_321),
.A2(n_271),
.B1(n_317),
.B2(n_252),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_372),
.B(n_374),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

CKINVDCx8_ASAP7_75t_R g464 ( 
.A(n_326),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_375),
.A2(n_262),
.B(n_254),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_261),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_327),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_426),
.B(n_329),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_380),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_398),
.B(n_344),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_400),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_417),
.A2(n_260),
.B1(n_313),
.B2(n_211),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_398),
.B(n_347),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_417),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_417),
.A2(n_357),
.B1(n_366),
.B2(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_419),
.B(n_350),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_399),
.B(n_379),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_416),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_417),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_419),
.B(n_355),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_426),
.B(n_360),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_399),
.B(n_363),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_427),
.B(n_230),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_365),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_399),
.B(n_261),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_409),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_444),
.B(n_373),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_421),
.B(n_381),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_464),
.B(n_386),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_436),
.B(n_384),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_405),
.B(n_377),
.Y(n_512)
);

AND2x4_ASAP7_75t_SL g513 ( 
.A(n_451),
.B(n_328),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_397),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_434),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_465),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_436),
.B(n_384),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_429),
.A2(n_428),
.B1(n_459),
.B2(n_440),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_421),
.B(n_240),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_465),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_464),
.B(n_435),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_397),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_436),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_241),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_431),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_450),
.A2(n_313),
.B1(n_211),
.B2(n_260),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_437),
.B(n_244),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_464),
.B(n_351),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_422),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_467),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_405),
.B(n_248),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_435),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_411),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_423),
.B(n_265),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_431),
.Y(n_547)
);

INVxp33_ASAP7_75t_SL g548 ( 
.A(n_428),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_423),
.B(n_269),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_457),
.B(n_385),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_459),
.A2(n_388),
.B1(n_342),
.B2(n_334),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_423),
.B(n_275),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_423),
.B(n_281),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_431),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_450),
.A2(n_271),
.B1(n_272),
.B2(n_317),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_411),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_411),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_427),
.B(n_406),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_427),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_406),
.B(n_387),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

INVxp33_ASAP7_75t_SL g564 ( 
.A(n_429),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_455),
.B(n_388),
.Y(n_566)
);

CKINVDCx11_ASAP7_75t_R g567 ( 
.A(n_427),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_441),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_454),
.A2(n_225),
.B1(n_319),
.B2(n_216),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_455),
.B(n_234),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_411),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_423),
.B(n_287),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_454),
.A2(n_273),
.B1(n_231),
.B2(n_238),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_422),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_463),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_463),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_450),
.B(n_234),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_430),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_460),
.B(n_230),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_450),
.B(n_188),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_401),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_450),
.B(n_288),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_401),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_450),
.B(n_234),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_439),
.B(n_292),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_401),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_441),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_430),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_411),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_441),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_430),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_432),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_460),
.B(n_203),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_403),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_432),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_403),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_403),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_457),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_458),
.B(n_299),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_441),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_432),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_439),
.B(n_294),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_458),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_404),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_458),
.B(n_299),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_412),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_458),
.A2(n_272),
.B1(n_254),
.B2(n_262),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_439),
.B(n_296),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_460),
.B(n_204),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_404),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_460),
.B(n_205),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_480),
.B(n_460),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_483),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_613),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_458),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_490),
.B(n_599),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_490),
.B(n_439),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_208),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_468),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_613),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_497),
.B(n_276),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_550),
.B(n_457),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_439),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_486),
.A2(n_305),
.B(n_279),
.C(n_283),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_468),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_609),
.B(n_261),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_491),
.B(n_213),
.C(n_209),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_497),
.B(n_276),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_618),
.B(n_439),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_569),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_519),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_483),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_469),
.B(n_237),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_609),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_472),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_542),
.B(n_442),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_569),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_604),
.B(n_461),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_520),
.A2(n_279),
.B1(n_283),
.B2(n_277),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_530),
.B(n_442),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_570),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_530),
.B(n_442),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_473),
.B(n_243),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_564),
.A2(n_524),
.B1(n_548),
.B2(n_523),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_478),
.A2(n_446),
.B1(n_442),
.B2(n_297),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_488),
.B(n_442),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_495),
.B(n_442),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_471),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_540),
.B(n_251),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_446),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_575),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_511),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_578),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_507),
.B(n_446),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_520),
.A2(n_277),
.B1(n_305),
.B2(n_446),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_526),
.B(n_446),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_476),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_502),
.B(n_584),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_476),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_531),
.B(n_446),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_472),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_585),
.A2(n_246),
.B1(n_195),
.B2(n_198),
.Y(n_674)
);

OAI221xp5_ASAP7_75t_L g675 ( 
.A1(n_475),
.A2(n_310),
.B1(n_264),
.B2(n_316),
.C(n_300),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_532),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_579),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_525),
.A2(n_420),
.B(n_229),
.C(n_218),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_519),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_479),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_535),
.B(n_452),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_563),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_579),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_511),
.B(n_461),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_544),
.A2(n_198),
.B1(n_316),
.B2(n_310),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_525),
.B(n_448),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

AO221x1_ASAP7_75t_L g688 ( 
.A1(n_524),
.A2(n_246),
.B1(n_218),
.B2(n_229),
.C(n_235),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_505),
.B(n_256),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_581),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_502),
.B(n_235),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_581),
.B(n_452),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_471),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_523),
.B(n_461),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_527),
.A2(n_300),
.B1(n_245),
.B2(n_264),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_586),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_529),
.B(n_257),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_532),
.B(n_452),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_547),
.B(n_452),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_605),
.A2(n_245),
.B1(n_242),
.B2(n_456),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_522),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_479),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_527),
.A2(n_242),
.B1(n_420),
.B2(n_456),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_586),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_474),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_588),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_474),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_477),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_547),
.B(n_452),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_534),
.B(n_456),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_534),
.B(n_456),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_588),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_481),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_536),
.B(n_404),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_410),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_497),
.B(n_385),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_538),
.A2(n_420),
.B1(n_453),
.B2(n_394),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_477),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_591),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_410),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_482),
.B(n_391),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_587),
.A2(n_608),
.B1(n_615),
.B2(n_590),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_470),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_484),
.B(n_391),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_506),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_482),
.B(n_410),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_485),
.B(n_415),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_481),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_485),
.B(n_415),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_496),
.B(n_415),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_497),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_560),
.B(n_453),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_591),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_506),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_493),
.B(n_227),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_528),
.B(n_392),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_496),
.B(n_424),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_499),
.B(n_424),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_499),
.B(n_424),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_489),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_497),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_559),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_559),
.B(n_392),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_503),
.A2(n_453),
.B1(n_395),
.B2(n_394),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_R g745 ( 
.A(n_529),
.B(n_258),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_494),
.B(n_259),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_503),
.B(n_425),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_600),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_600),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_602),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_572),
.B(n_393),
.C(n_293),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_508),
.B(n_425),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_498),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_602),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_508),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_SL g756 ( 
.A(n_592),
.B(n_266),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_514),
.Y(n_757)
);

O2A1O1Ixp5_ASAP7_75t_L g758 ( 
.A1(n_541),
.A2(n_418),
.B(n_425),
.C(n_447),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_513),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_514),
.A2(n_393),
.B(n_449),
.C(n_290),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_517),
.B(n_443),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_517),
.B(n_443),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_518),
.B(n_541),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_513),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_518),
.B(n_443),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_506),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_506),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_553),
.B(n_445),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_493),
.B(n_267),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_493),
.B(n_270),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_559),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_489),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_533),
.B(n_311),
.C(n_291),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_516),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_553),
.B(n_445),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_555),
.A2(n_227),
.B1(n_223),
.B2(n_201),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_603),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_555),
.A2(n_449),
.B(n_286),
.C(n_309),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_562),
.B(n_448),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_562),
.B(n_445),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_487),
.B(n_448),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_487),
.B(n_448),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_506),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_611),
.A2(n_466),
.B1(n_447),
.B2(n_201),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_545),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_603),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_610),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_623),
.A2(n_549),
.B(n_546),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_670),
.A2(n_554),
.B(n_552),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_758),
.A2(n_574),
.B(n_610),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_640),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_764),
.A2(n_595),
.B(n_487),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_762),
.B(n_561),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_760),
.A2(n_617),
.B(n_582),
.C(n_589),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_663),
.B(n_559),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_775),
.B(n_560),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_622),
.A2(n_617),
.B(n_502),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_641),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_644),
.B(n_493),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_619),
.A2(n_624),
.B(n_698),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_695),
.A2(n_614),
.B1(n_556),
.B2(n_502),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_666),
.A2(n_595),
.B(n_568),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_640),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_762),
.B(n_502),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_625),
.B(n_502),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_631),
.A2(n_595),
.B(n_568),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_625),
.B(n_566),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_637),
.A2(n_487),
.B(n_568),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_658),
.A2(n_595),
.B(n_568),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_682),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_684),
.B(n_509),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_643),
.B(n_492),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_663),
.B(n_559),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_651),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_644),
.B(n_606),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_675),
.A2(n_571),
.B(n_576),
.C(n_537),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_SL g818 ( 
.A1(n_760),
.A2(n_580),
.B(n_607),
.C(n_601),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_645),
.B(n_551),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_787),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_643),
.B(n_492),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_654),
.B(n_492),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_620),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_SL g825 ( 
.A(n_689),
.B(n_274),
.C(n_308),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_654),
.B(n_492),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_658),
.A2(n_606),
.B(n_545),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_682),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_647),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_695),
.A2(n_278),
.B(n_280),
.C(n_301),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_649),
.A2(n_312),
.B(n_307),
.C(n_306),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_668),
.A2(n_606),
.B(n_545),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_722),
.A2(n_606),
.B1(n_500),
.B2(n_557),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_644),
.B(n_592),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_687),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_672),
.A2(n_545),
.B(n_596),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_646),
.A2(n_545),
.B(n_596),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_788),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_699),
.A2(n_500),
.B(n_521),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_734),
.A2(n_592),
.B(n_596),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_673),
.B(n_303),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_687),
.A2(n_504),
.B(n_607),
.C(n_601),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_652),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_701),
.B(n_567),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_694),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_759),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_765),
.B(n_639),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_734),
.A2(n_767),
.B(n_676),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_767),
.A2(n_592),
.B(n_596),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_676),
.A2(n_592),
.B(n_596),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_676),
.A2(n_711),
.B(n_710),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_620),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_630),
.B(n_521),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_592),
.B(n_596),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_662),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_644),
.B(n_521),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_689),
.A2(n_521),
.B1(n_557),
.B2(n_594),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_725),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_657),
.B(n_557),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_621),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_664),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_736),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_681),
.A2(n_661),
.B(n_709),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_665),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_693),
.B(n_557),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_782),
.A2(n_558),
.B(n_573),
.Y(n_866)
);

OAI321xp33_ASAP7_75t_L g867 ( 
.A1(n_777),
.A2(n_447),
.A3(n_449),
.B1(n_295),
.B2(n_263),
.C(n_223),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_677),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_782),
.A2(n_558),
.B(n_573),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_783),
.A2(n_558),
.B(n_573),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_783),
.A2(n_558),
.B(n_573),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_693),
.B(n_594),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_649),
.A2(n_449),
.B(n_598),
.C(n_597),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_627),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_736),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_705),
.B(n_707),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_705),
.B(n_594),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_628),
.B(n_594),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_686),
.A2(n_612),
.B(n_598),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_746),
.A2(n_612),
.B(n_597),
.C(n_593),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_721),
.B(n_612),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_686),
.A2(n_612),
.B(n_593),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_735),
.B(n_299),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_780),
.A2(n_779),
.B(n_727),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_683),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_780),
.A2(n_583),
.B(n_580),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_501),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_650),
.A2(n_583),
.B(n_577),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_724),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_632),
.A2(n_577),
.B(n_565),
.C(n_543),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_708),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_638),
.B(n_642),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_708),
.B(n_501),
.Y(n_893)
);

AO21x1_ASAP7_75t_L g894 ( 
.A1(n_634),
.A2(n_565),
.B(n_543),
.Y(n_894)
);

CKINVDCx8_ASAP7_75t_R g895 ( 
.A(n_731),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_718),
.B(n_504),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_718),
.B(n_510),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_690),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_732),
.B(n_65),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_729),
.B(n_726),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_656),
.A2(n_539),
.B1(n_510),
.B2(n_466),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_653),
.A2(n_539),
.B(n_396),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_755),
.B(n_418),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_730),
.A2(n_396),
.B(n_402),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_737),
.A2(n_396),
.B(n_402),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_738),
.A2(n_408),
.B(n_396),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_755),
.B(n_659),
.Y(n_907)
);

NOR2x1_ASAP7_75t_L g908 ( 
.A(n_635),
.B(n_743),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_659),
.B(n_448),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_739),
.A2(n_402),
.B(n_407),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_746),
.A2(n_418),
.B(n_438),
.C(n_433),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_747),
.A2(n_402),
.B(n_407),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_667),
.A2(n_418),
.B1(n_448),
.B2(n_438),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_752),
.A2(n_407),
.B(n_408),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_678),
.A2(n_408),
.B(n_407),
.C(n_418),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_753),
.A2(n_466),
.B1(n_441),
.B2(n_448),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_716),
.B(n_66),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_634),
.A2(n_433),
.B(n_432),
.C(n_438),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_761),
.A2(n_408),
.B(n_433),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_697),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_L g921 ( 
.A1(n_660),
.A2(n_438),
.B(n_433),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_763),
.A2(n_441),
.B(n_466),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_766),
.A2(n_414),
.B(n_412),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_770),
.A2(n_3),
.B(n_5),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_660),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_725),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_770),
.B(n_771),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_696),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_771),
.B(n_201),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_757),
.B(n_448),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_757),
.B(n_448),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_655),
.B(n_412),
.C(n_414),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_731),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_725),
.A2(n_414),
.B(n_412),
.Y(n_934)
);

AO21x2_ASAP7_75t_L g935 ( 
.A1(n_678),
.A2(n_295),
.B(n_263),
.Y(n_935)
);

AOI21xp33_ASAP7_75t_L g936 ( 
.A1(n_777),
.A2(n_9),
.B(n_11),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_697),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_704),
.B(n_414),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_706),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_712),
.B(n_414),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_719),
.B(n_414),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_725),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_768),
.A2(n_414),
.B(n_412),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_768),
.B(n_201),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_733),
.B(n_748),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_768),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_667),
.A2(n_749),
.B1(n_750),
.B2(n_754),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_632),
.A2(n_223),
.B(n_263),
.C(n_295),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_768),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_778),
.B(n_744),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_744),
.B(n_414),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_731),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_786),
.A2(n_414),
.B(n_412),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_786),
.A2(n_412),
.B(n_441),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_674),
.A2(n_223),
.B(n_263),
.C(n_295),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_786),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_685),
.A2(n_745),
.B(n_774),
.Y(n_957)
);

BUFx8_ASAP7_75t_L g958 ( 
.A(n_721),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_786),
.A2(n_412),
.B(n_441),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_714),
.A2(n_412),
.B(n_441),
.Y(n_960)
);

CKINVDCx10_ASAP7_75t_R g961 ( 
.A(n_629),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_784),
.B(n_116),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_721),
.B(n_466),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_721),
.B(n_466),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_716),
.B(n_160),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_745),
.A2(n_9),
.B(n_11),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_715),
.A2(n_466),
.B(n_157),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_720),
.A2(n_12),
.B(n_16),
.C(n_21),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_626),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_769),
.A2(n_466),
.B(n_155),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_721),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_743),
.B(n_23),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_633),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_751),
.A2(n_466),
.B1(n_153),
.B2(n_151),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_703),
.A2(n_106),
.B1(n_147),
.B2(n_146),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_832),
.A2(n_703),
.B(n_781),
.Y(n_976)
);

OAI22x1_ASAP7_75t_L g977 ( 
.A1(n_820),
.A2(n_700),
.B1(n_785),
.B2(n_743),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_808),
.A2(n_925),
.B1(n_950),
.B2(n_927),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_937),
.B(n_772),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_797),
.B(n_772),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_925),
.A2(n_772),
.B1(n_742),
.B2(n_776),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_887),
.B(n_751),
.Y(n_982)
);

BUFx6f_ASAP7_75t_SL g983 ( 
.A(n_828),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_887),
.B(n_688),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_812),
.B(n_741),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_813),
.A2(n_692),
.B(n_756),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_817),
.A2(n_957),
.B(n_929),
.C(n_795),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_844),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_L g989 ( 
.A1(n_795),
.A2(n_773),
.B(n_669),
.C(n_671),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_936),
.A2(n_629),
.B(n_636),
.C(n_716),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_862),
.B(n_741),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_924),
.A2(n_629),
.B(n_636),
.C(n_691),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_825),
.A2(n_636),
.B1(n_742),
.B2(n_741),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_920),
.B(n_742),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_933),
.B(n_740),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_811),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_825),
.A2(n_717),
.B1(n_728),
.B2(n_713),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_862),
.A2(n_702),
.B1(n_680),
.B2(n_466),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_792),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_799),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_895),
.B(n_102),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_917),
.B(n_133),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_889),
.B(n_875),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_845),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_875),
.B(n_129),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_794),
.B(n_25),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_835),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_SL g1009 ( 
.A(n_796),
.B(n_814),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_819),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_858),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_807),
.A2(n_809),
.B(n_863),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_900),
.A2(n_117),
.B(n_115),
.C(n_107),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_802),
.A2(n_103),
.B1(n_96),
.B2(n_95),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_829),
.B(n_26),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_796),
.B(n_93),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_816),
.A2(n_87),
.B(n_68),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_952),
.B(n_814),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_822),
.A2(n_27),
.B(n_30),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_961),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_888),
.A2(n_33),
.B(n_35),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_835),
.B(n_33),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_816),
.A2(n_35),
.B(n_36),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_955),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_847),
.B(n_820),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_858),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_SL g1027 ( 
.A1(n_972),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_883),
.B(n_917),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_841),
.A2(n_45),
.B(n_46),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_965),
.B(n_47),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_858),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_843),
.B(n_51),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_841),
.B(n_51),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_860),
.B(n_54),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_855),
.B(n_54),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_861),
.B(n_57),
.Y(n_1036)
);

CKINVDCx6p67_ASAP7_75t_R g1037 ( 
.A(n_846),
.Y(n_1037)
);

AOI33xp33_ASAP7_75t_L g1038 ( 
.A1(n_968),
.A2(n_58),
.A3(n_61),
.B1(n_63),
.B2(n_64),
.B3(n_864),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_965),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_810),
.A2(n_63),
.B(n_851),
.Y(n_1040)
);

AO32x2_ASAP7_75t_L g1041 ( 
.A1(n_947),
.A2(n_975),
.A3(n_913),
.B1(n_818),
.B2(n_946),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_860),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_802),
.A2(n_932),
.B1(n_806),
.B2(n_945),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_926),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_955),
.A2(n_966),
.B(n_830),
.C(n_831),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_874),
.B(n_838),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_815),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_SL g1048 ( 
.A(n_958),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_SL g1049 ( 
.A(n_948),
.B(n_972),
.C(n_974),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_926),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_830),
.A2(n_831),
.B(n_867),
.C(n_944),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_944),
.B(n_800),
.C(n_805),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_881),
.A2(n_793),
.B(n_823),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_868),
.B(n_885),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_908),
.B(n_800),
.C(n_789),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_898),
.B(n_928),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_958),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_926),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_971),
.A2(n_852),
.B1(n_824),
.B2(n_907),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_884),
.A2(n_791),
.B(n_839),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_801),
.A2(n_798),
.B(n_859),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_939),
.B(n_899),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_821),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_926),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_826),
.A2(n_790),
.B(n_827),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_876),
.A2(n_891),
.B(n_848),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_878),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_824),
.B(n_852),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_880),
.A2(n_915),
.B(n_911),
.C(n_853),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_969),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_962),
.Y(n_1071)
);

AO21x1_ASAP7_75t_L g1072 ( 
.A1(n_859),
.A2(n_842),
.B(n_890),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_971),
.B(n_973),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_915),
.A2(n_818),
.B(n_873),
.C(n_921),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_836),
.A2(n_837),
.B(n_856),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_865),
.A2(n_877),
.B(n_872),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_942),
.B(n_949),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_893),
.B(n_897),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_896),
.B(n_892),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_930),
.A2(n_931),
.B(n_909),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_942),
.B(n_949),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_909),
.A2(n_869),
.B(n_871),
.Y(n_1082)
);

BUFx8_ASAP7_75t_SL g1083 ( 
.A(n_942),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_894),
.A2(n_906),
.B(n_918),
.C(n_967),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_942),
.B(n_949),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_833),
.A2(n_857),
.B1(n_892),
.B2(n_951),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_903),
.B(n_949),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_956),
.A2(n_946),
.B1(n_834),
.B2(n_962),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_866),
.A2(n_870),
.B(n_850),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_854),
.A2(n_840),
.B(n_849),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_901),
.A2(n_902),
.B(n_879),
.C(n_882),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_956),
.B(n_873),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_938),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_956),
.B(n_940),
.Y(n_1094)
);

AND2x4_ASAP7_75t_SL g1095 ( 
.A(n_956),
.B(n_916),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_941),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_904),
.A2(n_914),
.B(n_905),
.C(n_910),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_834),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_886),
.A2(n_912),
.B(n_919),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_963),
.A2(n_964),
.B1(n_935),
.B2(n_922),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_935),
.B(n_960),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_923),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_934),
.B(n_943),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_953),
.A2(n_954),
.B(n_959),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_970),
.A2(n_888),
.B(n_882),
.Y(n_1105)
);

BUFx12f_ASAP7_75t_L g1106 ( 
.A(n_828),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_936),
.A2(n_625),
.B(n_924),
.C(n_825),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_835),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_925),
.B(n_564),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_817),
.A2(n_625),
.B(n_808),
.C(n_486),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_917),
.B(n_731),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_811),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_804),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_813),
.A2(n_823),
.B(n_822),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_799),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_820),
.A2(n_524),
.B1(n_564),
.B2(n_523),
.C(n_548),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_832),
.A2(n_676),
.B(n_803),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_927),
.B(n_648),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_828),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1118),
.B(n_978),
.Y(n_1120)
);

NAND3x1_ASAP7_75t_L g1121 ( 
.A(n_1116),
.B(n_1109),
.C(n_1033),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1054),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_987),
.A2(n_1072),
.A3(n_1110),
.B(n_1086),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1012),
.A2(n_1065),
.B(n_1053),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1109),
.A2(n_1027),
.B1(n_1039),
.B2(n_1057),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1020),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1117),
.A2(n_1089),
.B(n_1082),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1043),
.A2(n_1091),
.A3(n_1040),
.B(n_1097),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1106),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_1061),
.A2(n_1084),
.B(n_1021),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1025),
.A2(n_982),
.B1(n_1111),
.B2(n_1039),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_976),
.A2(n_1066),
.B(n_1075),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1107),
.A2(n_1028),
.B(n_1007),
.C(n_1029),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_SL g1134 ( 
.A(n_1010),
.B(n_1115),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1083),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1069),
.A2(n_989),
.B(n_1076),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_997),
.B(n_1112),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_988),
.B(n_1004),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_983),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1060),
.A2(n_1078),
.B(n_1090),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_990),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1105),
.A2(n_1104),
.B(n_989),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1103),
.A2(n_977),
.A3(n_1092),
.B(n_1094),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1007),
.B(n_984),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1099),
.A2(n_1080),
.B(n_1074),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1070),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1060),
.A2(n_1102),
.B(n_1062),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1055),
.B(n_1094),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_1014),
.A2(n_1006),
.B(n_1016),
.C(n_1051),
.Y(n_1150)
);

AND2x6_ASAP7_75t_SL g1151 ( 
.A(n_1034),
.B(n_1022),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1084),
.A2(n_1114),
.B(n_1013),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_SL g1153 ( 
.A1(n_1003),
.A2(n_980),
.B1(n_1034),
.B2(n_1004),
.Y(n_1153)
);

BUFx4f_ASAP7_75t_SL g1154 ( 
.A(n_1037),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1059),
.A2(n_1079),
.A3(n_1088),
.B(n_1023),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_1030),
.A2(n_994),
.B1(n_1022),
.B2(n_1108),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1100),
.A2(n_1013),
.B(n_1102),
.Y(n_1157)
);

OA21x2_ASAP7_75t_L g1158 ( 
.A1(n_1052),
.A2(n_1055),
.B(n_986),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1046),
.B(n_1073),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1119),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1049),
.A2(n_1024),
.B(n_1045),
.C(n_1036),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_990),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1087),
.A2(n_985),
.B(n_992),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1042),
.B(n_1008),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1005),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1015),
.A2(n_1032),
.B(n_1035),
.C(n_991),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_1052),
.A2(n_998),
.B(n_1019),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1017),
.A2(n_1081),
.B1(n_1009),
.B2(n_1046),
.C(n_979),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_998),
.A2(n_999),
.B(n_993),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1073),
.B(n_1113),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1111),
.A2(n_1095),
.B(n_1077),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1085),
.A2(n_1056),
.B(n_1063),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1027),
.B(n_1038),
.C(n_1108),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1111),
.A2(n_1071),
.B1(n_1047),
.B2(n_1008),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1098),
.A2(n_1068),
.B(n_996),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1003),
.A2(n_995),
.B1(n_1001),
.B2(n_1018),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1018),
.B(n_996),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1067),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_983),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1098),
.A2(n_1003),
.B(n_1041),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1003),
.A2(n_1041),
.B(n_1050),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1003),
.A2(n_1041),
.B(n_1050),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1101),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1026),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1026),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1068),
.A2(n_1101),
.B(n_1064),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1026),
.A2(n_1058),
.B(n_1064),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1041),
.A2(n_1044),
.B(n_1026),
.Y(n_1188)
);

CKINVDCx9p33_ASAP7_75t_R g1189 ( 
.A(n_1048),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_980),
.A2(n_1058),
.B(n_1064),
.C(n_1002),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1058),
.A2(n_1064),
.B(n_1002),
.C(n_1048),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1044),
.A2(n_800),
.B(n_986),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_625),
.B1(n_1116),
.B2(n_1109),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_997),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1025),
.B(n_927),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1012),
.A2(n_1065),
.B(n_1053),
.Y(n_1197)
);

AOI211x1_ASAP7_75t_L g1198 ( 
.A1(n_1029),
.A2(n_936),
.B(n_924),
.C(n_966),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1025),
.B(n_936),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1101),
.A2(n_1055),
.B(n_987),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1110),
.A2(n_987),
.B(n_1107),
.Y(n_1201)
);

AND2x6_ASAP7_75t_L g1202 ( 
.A(n_1071),
.B(n_917),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1107),
.A2(n_1110),
.B(n_817),
.C(n_625),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1049),
.A2(n_927),
.B1(n_978),
.B2(n_825),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1110),
.A2(n_987),
.B(n_808),
.C(n_936),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1118),
.B(n_978),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1118),
.B(n_978),
.Y(n_1210)
);

AO32x2_ASAP7_75t_L g1211 ( 
.A1(n_978),
.A2(n_1043),
.A3(n_1086),
.B1(n_981),
.B2(n_524),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1118),
.B(n_978),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1214)
);

AOI221xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1029),
.A2(n_1107),
.B1(n_817),
.B2(n_1110),
.C(n_1045),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_987),
.A2(n_1072),
.A3(n_1110),
.B(n_1086),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1110),
.A2(n_625),
.B(n_1107),
.C(n_925),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1110),
.A2(n_695),
.B1(n_802),
.B2(n_649),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_1110),
.B(n_817),
.C(n_625),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1109),
.B(n_925),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1010),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_987),
.A2(n_1072),
.A3(n_1110),
.B(n_1086),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1025),
.A2(n_625),
.B1(n_1116),
.B2(n_1109),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1025),
.B(n_927),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_987),
.A2(n_1072),
.A3(n_1110),
.B(n_1086),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1010),
.Y(n_1233)
);

CKINVDCx11_ASAP7_75t_R g1234 ( 
.A(n_1106),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1000),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1118),
.B(n_978),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_775),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1106),
.B(n_775),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_990),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_987),
.A2(n_1072),
.A3(n_1110),
.B(n_1086),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1018),
.B(n_933),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1054),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1110),
.A2(n_695),
.B1(n_802),
.B2(n_649),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1107),
.A2(n_1110),
.B(n_817),
.C(n_625),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1083),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1109),
.B(n_925),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_990),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1110),
.A2(n_695),
.B1(n_802),
.B2(n_649),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_990),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1101),
.A2(n_1055),
.B(n_987),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1110),
.A2(n_987),
.B(n_1107),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1110),
.A2(n_987),
.B(n_1107),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1118),
.B(n_1109),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1025),
.A2(n_625),
.B(n_564),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1083),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1110),
.A2(n_695),
.B1(n_802),
.B2(n_649),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1109),
.B(n_925),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1012),
.A2(n_1117),
.B(n_1053),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1117),
.A2(n_1012),
.B(n_1089),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1110),
.A2(n_987),
.B(n_1107),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1256),
.A2(n_1193),
.B1(n_1228),
.B2(n_1199),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1199),
.A2(n_1125),
.B1(n_1218),
.B2(n_1258),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1218),
.A2(n_1244),
.B1(n_1258),
.B2(n_1249),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1145),
.A2(n_1262),
.B1(n_1253),
.B2(n_1252),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1244),
.A2(n_1249),
.B1(n_1259),
.B2(n_1247),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1250),
.Y(n_1268)
);

INVx5_ASAP7_75t_L g1269 ( 
.A(n_1202),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1250),
.B(n_1186),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1121),
.A2(n_1153),
.B1(n_1221),
.B2(n_1145),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1196),
.A2(n_1230),
.B1(n_1159),
.B2(n_1176),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1139),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1173),
.A2(n_1262),
.B1(n_1201),
.B2(n_1253),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1201),
.A2(n_1252),
.B1(n_1173),
.B2(n_1206),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1131),
.A2(n_1254),
.B1(n_1156),
.B2(n_1215),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1234),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1194),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1141),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1177),
.B(n_1242),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1159),
.A2(n_1120),
.B1(n_1210),
.B2(n_1213),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1160),
.Y(n_1282)
);

CKINVDCx6p67_ASAP7_75t_R g1283 ( 
.A(n_1135),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1235),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1203),
.A2(n_1220),
.B(n_1245),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1122),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1165),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1126),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1120),
.A2(n_1213),
.B1(n_1236),
.B2(n_1208),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1212),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1208),
.A2(n_1210),
.B1(n_1236),
.B2(n_1149),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1206),
.A2(n_1169),
.B1(n_1251),
.B2(n_1200),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1139),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1202),
.A2(n_1174),
.B1(n_1177),
.B2(n_1151),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1135),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1169),
.A2(n_1251),
.B1(n_1200),
.B2(n_1149),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1243),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1179),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1202),
.A2(n_1157),
.B1(n_1167),
.B2(n_1178),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1202),
.A2(n_1157),
.B1(n_1167),
.B2(n_1144),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1170),
.A2(n_1174),
.B1(n_1136),
.B2(n_1198),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1170),
.A2(n_1136),
.B1(n_1215),
.B2(n_1180),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1179),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_1237),
.Y(n_1304)
);

INVx11_ASAP7_75t_L g1305 ( 
.A(n_1154),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1137),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1168),
.A2(n_1138),
.B1(n_1135),
.B2(n_1246),
.Y(n_1307)
);

CKINVDCx9p33_ASAP7_75t_R g1308 ( 
.A(n_1226),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1180),
.A2(n_1246),
.B1(n_1257),
.B2(n_1181),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1172),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1133),
.B(n_1217),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1246),
.A2(n_1171),
.B1(n_1175),
.B2(n_1181),
.Y(n_1312)
);

INVx4_ASAP7_75t_SL g1313 ( 
.A(n_1143),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1242),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1129),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1224),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1191),
.A2(n_1186),
.B1(n_1166),
.B2(n_1161),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1233),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1143),
.B(n_1134),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1188),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1141),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1148),
.A2(n_1182),
.B1(n_1158),
.B2(n_1163),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1182),
.A2(n_1158),
.B1(n_1130),
.B2(n_1211),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1150),
.A2(n_1211),
.B1(n_1207),
.B2(n_1152),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1130),
.A2(n_1211),
.B1(n_1152),
.B2(n_1140),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1141),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1146),
.A2(n_1132),
.B1(n_1124),
.B2(n_1197),
.Y(n_1327)
);

INVx8_ASAP7_75t_L g1328 ( 
.A(n_1184),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1184),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1238),
.A2(n_1239),
.B1(n_1248),
.B2(n_1162),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1124),
.A2(n_1197),
.B1(n_1205),
.B2(n_1260),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1192),
.B(n_1214),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1248),
.A2(n_1185),
.B1(n_1216),
.B2(n_1227),
.Y(n_1333)
);

BUFx2_ASAP7_75t_SL g1334 ( 
.A(n_1187),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1183),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1190),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1204),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1232),
.B(n_1255),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1155),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1155),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1123),
.A2(n_1240),
.B1(n_1231),
.B2(n_1227),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1123),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1216),
.A2(n_1240),
.B1(n_1231),
.B2(n_1227),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1231),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1240),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1127),
.A2(n_1142),
.B1(n_1222),
.B2(n_1195),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1128),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1128),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1209),
.A2(n_1219),
.B1(n_1223),
.B2(n_1225),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1229),
.A2(n_1025),
.B1(n_1199),
.B2(n_1125),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1241),
.Y(n_1351)
);

INVx4_ASAP7_75t_SL g1352 ( 
.A(n_1261),
.Y(n_1352)
);

BUFx4f_ASAP7_75t_L g1353 ( 
.A(n_1135),
.Y(n_1353)
);

CKINVDCx6p67_ASAP7_75t_R g1354 ( 
.A(n_1189),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1126),
.Y(n_1355)
);

INVx8_ASAP7_75t_L g1356 ( 
.A(n_1250),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1164),
.Y(n_1357)
);

CKINVDCx16_ASAP7_75t_R g1358 ( 
.A(n_1135),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1126),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1160),
.Y(n_1360)
);

OAI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1193),
.A2(n_625),
.B(n_1228),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1234),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1147),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1193),
.B(n_1228),
.Y(n_1364)
);

BUFx4_ASAP7_75t_SL g1365 ( 
.A(n_1126),
.Y(n_1365)
);

CKINVDCx6p67_ASAP7_75t_R g1366 ( 
.A(n_1189),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1256),
.A2(n_1193),
.B1(n_1228),
.B2(n_1199),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1234),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1256),
.A2(n_1193),
.B1(n_1228),
.B2(n_1199),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1256),
.A2(n_1193),
.B1(n_1228),
.B2(n_1199),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1139),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1199),
.A2(n_1025),
.B1(n_1125),
.B2(n_564),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1147),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1147),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1256),
.A2(n_1193),
.B1(n_1228),
.B2(n_1199),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1147),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1234),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1342),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1277),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1273),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1269),
.B(n_1335),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1344),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1347),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1269),
.B(n_1313),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1296),
.B(n_1265),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1348),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1332),
.A2(n_1346),
.B(n_1327),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1320),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1320),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1365),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1310),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1296),
.B(n_1275),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1339),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1340),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1306),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1292),
.B(n_1319),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1292),
.B(n_1275),
.Y(n_1397)
);

CKINVDCx12_ASAP7_75t_R g1398 ( 
.A(n_1294),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1364),
.A2(n_1361),
.B1(n_1367),
.B2(n_1369),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1267),
.B(n_1266),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1270),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1357),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1343),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1343),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1352),
.Y(n_1405)
);

CKINVDCx12_ASAP7_75t_R g1406 ( 
.A(n_1365),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1332),
.A2(n_1338),
.B(n_1285),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1266),
.B(n_1274),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1270),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1346),
.A2(n_1327),
.B(n_1349),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1284),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1363),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1338),
.A2(n_1333),
.B(n_1311),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1373),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1337),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1374),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1317),
.B(n_1351),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1273),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1376),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1372),
.A2(n_1370),
.B1(n_1367),
.B2(n_1369),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1364),
.A2(n_1263),
.B(n_1375),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1333),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1351),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1312),
.A2(n_1289),
.B(n_1291),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1370),
.A2(n_1375),
.B1(n_1264),
.B2(n_1271),
.Y(n_1425)
);

AO21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1299),
.A2(n_1300),
.B(n_1323),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1349),
.A2(n_1331),
.B(n_1325),
.Y(n_1427)
);

INVxp33_ASAP7_75t_L g1428 ( 
.A(n_1360),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1278),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1287),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1341),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1345),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1341),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1281),
.Y(n_1434)
);

AO21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1299),
.A2(n_1300),
.B(n_1323),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1356),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1302),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1302),
.B(n_1322),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1324),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1356),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1273),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1350),
.A2(n_1272),
.B1(n_1276),
.B2(n_1309),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1312),
.A2(n_1301),
.B1(n_1307),
.B2(n_1282),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1301),
.B(n_1297),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1331),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1325),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1286),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1290),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1334),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1307),
.A2(n_1282),
.B1(n_1314),
.B2(n_1280),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1330),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1330),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1336),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1421),
.A2(n_1356),
.B(n_1353),
.C(n_1326),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1420),
.A2(n_1353),
.B(n_1321),
.C(n_1279),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1393),
.B(n_1358),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1425),
.A2(n_1326),
.B(n_1280),
.C(n_1371),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1399),
.A2(n_1316),
.B1(n_1293),
.B2(n_1304),
.C(n_1318),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1442),
.A2(n_1318),
.B(n_1329),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1394),
.B(n_1402),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1394),
.B(n_1329),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1424),
.A2(n_1326),
.B(n_1328),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1391),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1400),
.A2(n_1359),
.B(n_1355),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1384),
.B(n_1288),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1400),
.A2(n_1328),
.B1(n_1308),
.B2(n_1354),
.C(n_1366),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1384),
.B(n_1308),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1396),
.B(n_1283),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1408),
.A2(n_1303),
.B(n_1298),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1408),
.A2(n_1328),
.B(n_1268),
.C(n_1298),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.B(n_1298),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1429),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1438),
.B(n_1303),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1443),
.A2(n_1303),
.B(n_1268),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1415),
.B(n_1295),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1385),
.A2(n_1315),
.B1(n_1295),
.B2(n_1377),
.C(n_1362),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1415),
.B(n_1368),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1415),
.B(n_1305),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1453),
.A2(n_1450),
.B1(n_1432),
.B2(n_1395),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1385),
.A2(n_1449),
.B(n_1434),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1392),
.A2(n_1438),
.B(n_1397),
.C(n_1434),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1438),
.B(n_1446),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1410),
.A2(n_1387),
.B(n_1427),
.Y(n_1484)
);

INVx5_ASAP7_75t_L g1485 ( 
.A(n_1417),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1392),
.A2(n_1437),
.B1(n_1424),
.B2(n_1397),
.C(n_1439),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1396),
.B(n_1388),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1449),
.A2(n_1445),
.B(n_1427),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1432),
.A2(n_1430),
.B1(n_1428),
.B2(n_1437),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1391),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1431),
.B(n_1433),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1413),
.B(n_1422),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1413),
.B(n_1422),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1390),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1387),
.A2(n_1410),
.B(n_1403),
.Y(n_1497)
);

NAND4xp25_ASAP7_75t_L g1498 ( 
.A(n_1444),
.B(n_1448),
.C(n_1439),
.D(n_1451),
.Y(n_1498)
);

OAI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1417),
.A2(n_1445),
.B1(n_1432),
.B2(n_1452),
.C(n_1380),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1426),
.B(n_1435),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1435),
.B(n_1411),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1406),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1407),
.A2(n_1423),
.B(n_1382),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1482),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_1490),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1497),
.B(n_1493),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1490),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1504),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1504),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1454),
.B(n_1457),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1463),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1498),
.A2(n_1401),
.B1(n_1409),
.B2(n_1398),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1497),
.B(n_1403),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1497),
.B(n_1404),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1487),
.B(n_1404),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1493),
.B(n_1407),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1494),
.B(n_1407),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1463),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1494),
.B(n_1495),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1486),
.A2(n_1448),
.B1(n_1447),
.B2(n_1386),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1488),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1495),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1501),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1484),
.B(n_1383),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1458),
.A2(n_1447),
.B1(n_1412),
.B2(n_1419),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1484),
.B(n_1383),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1481),
.A2(n_1414),
.B1(n_1416),
.B2(n_1419),
.Y(n_1528)
);

BUFx8_ASAP7_75t_SL g1529 ( 
.A(n_1496),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1484),
.B(n_1378),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_L g1531 ( 
.A(n_1454),
.B(n_1405),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1512),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1521),
.A2(n_1481),
.B1(n_1457),
.B2(n_1480),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1525),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1505),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1521),
.B(n_1479),
.C(n_1489),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1528),
.A2(n_1476),
.B(n_1464),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1520),
.B(n_1501),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1519),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1523),
.B(n_1460),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1520),
.B(n_1483),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1509),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1506),
.B(n_1492),
.Y(n_1546)
);

AND4x1_ASAP7_75t_L g1547 ( 
.A(n_1511),
.B(n_1466),
.C(n_1455),
.D(n_1470),
.Y(n_1547)
);

OAI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1511),
.A2(n_1459),
.B1(n_1469),
.B2(n_1474),
.C(n_1499),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1508),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1528),
.B(n_1500),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1508),
.B(n_1492),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1510),
.A2(n_1462),
.B(n_1500),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1523),
.B(n_1491),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1507),
.B(n_1517),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1529),
.Y(n_1558)
);

OAI31xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1513),
.A2(n_1471),
.A3(n_1473),
.B(n_1467),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1549),
.B(n_1518),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1532),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1555),
.B(n_1514),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1555),
.B(n_1522),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1558),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1532),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1535),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1544),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1555),
.B(n_1514),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1534),
.B(n_1522),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1518),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1539),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1557),
.B(n_1517),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1536),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1522),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1534),
.B(n_1524),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.B(n_1524),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1534),
.B(n_1524),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1515),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1515),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1534),
.B(n_1505),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1536),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1477),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1546),
.B(n_1515),
.Y(n_1586)
);

INVx6_ASAP7_75t_L g1587 ( 
.A(n_1534),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1534),
.B(n_1505),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1553),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1541),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1544),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1542),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1554),
.B(n_1525),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1541),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1554),
.B(n_1525),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1587),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1593),
.B(n_1542),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1585),
.B(n_1538),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1593),
.B(n_1560),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1576),
.A2(n_1537),
.B1(n_1548),
.B2(n_1533),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1576),
.B(n_1543),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1560),
.B(n_1543),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1561),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1578),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1578),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1582),
.B(n_1550),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1564),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

AOI33xp33_ASAP7_75t_L g1621 ( 
.A1(n_1570),
.A2(n_1526),
.A3(n_1527),
.B1(n_1530),
.B2(n_1556),
.B3(n_1461),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1565),
.Y(n_1622)
);

OAI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1570),
.A2(n_1533),
.B(n_1559),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1564),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1565),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1551),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1566),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1564),
.A2(n_1548),
.B1(n_1398),
.B2(n_1467),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1586),
.B(n_1516),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1566),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1566),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_1580),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1567),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1564),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1572),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1574),
.B(n_1379),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1572),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1586),
.B(n_1516),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1572),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1602),
.B(n_1590),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1590),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1602),
.B(n_1590),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1605),
.B(n_1589),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1606),
.B(n_1580),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1607),
.B(n_1589),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1632),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1618),
.B(n_1581),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1632),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1606),
.B(n_1580),
.Y(n_1653)
);

CKINVDCx16_ASAP7_75t_R g1654 ( 
.A(n_1637),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

AND2x2_ASAP7_75t_SL g1657 ( 
.A(n_1621),
.B(n_1547),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1633),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1635),
.B(n_1529),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1634),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1634),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1619),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1613),
.B(n_1570),
.Y(n_1665)
);

AOI31xp33_ASAP7_75t_L g1666 ( 
.A1(n_1624),
.A2(n_1502),
.A3(n_1406),
.B(n_1456),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1600),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1625),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1633),
.B(n_1575),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1627),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1604),
.B(n_1573),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1621),
.B(n_1573),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1631),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1636),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1599),
.B(n_1568),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1659),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1664),
.B(n_1623),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1654),
.B(n_1628),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1654),
.B(n_1628),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1646),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1658),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1657),
.A2(n_1603),
.B1(n_1610),
.B2(n_1616),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1664),
.Y(n_1688)
);

OAI31xp33_ASAP7_75t_L g1689 ( 
.A1(n_1673),
.A2(n_1575),
.A3(n_1616),
.B(n_1610),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1616),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1672),
.A2(n_1547),
.B1(n_1559),
.B2(n_1600),
.C(n_1587),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1666),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1673),
.A2(n_1587),
.B1(n_1615),
.B2(n_1612),
.C(n_1611),
.Y(n_1694)
);

O2A1O1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1666),
.A2(n_1575),
.B(n_1574),
.C(n_1584),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1658),
.B(n_1595),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1657),
.A2(n_1587),
.B1(n_1569),
.B2(n_1562),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1646),
.B(n_1595),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1641),
.A2(n_1587),
.B1(n_1485),
.B2(n_1617),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1667),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1641),
.A2(n_1587),
.B1(n_1531),
.B2(n_1467),
.Y(n_1701)
);

AOI222xp33_ASAP7_75t_L g1702 ( 
.A1(n_1645),
.A2(n_1472),
.B1(n_1526),
.B2(n_1584),
.C1(n_1597),
.C2(n_1595),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1682),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1692),
.A2(n_1645),
.B(n_1644),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1695),
.A2(n_1649),
.B(n_1676),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1669),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1683),
.A2(n_1669),
.B1(n_1649),
.B2(n_1665),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1683),
.A2(n_1665),
.B1(n_1647),
.B2(n_1653),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1676),
.B(n_1644),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1677),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1684),
.A2(n_1653),
.B1(n_1642),
.B2(n_1647),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1681),
.B(n_1502),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1688),
.B(n_1690),
.Y(n_1717)
);

O2A1O1Ixp5_ASAP7_75t_L g1718 ( 
.A1(n_1678),
.A2(n_1675),
.B(n_1674),
.C(n_1656),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1698),
.B(n_1686),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1689),
.A2(n_1675),
.B1(n_1656),
.B2(n_1674),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1677),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1704),
.B(n_1700),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1706),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1703),
.B(n_1700),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1720),
.A2(n_1691),
.B1(n_1701),
.B2(n_1680),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1703),
.B(n_1687),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1716),
.A2(n_1702),
.B(n_1697),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1699),
.B1(n_1696),
.B2(n_1651),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1708),
.A2(n_1696),
.B1(n_1679),
.B2(n_1693),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1720),
.A2(n_1660),
.B1(n_1651),
.B2(n_1671),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_L g1731 ( 
.A(n_1717),
.B(n_1496),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1705),
.A2(n_1693),
.B(n_1679),
.Y(n_1732)
);

NAND3x1_ASAP7_75t_L g1733 ( 
.A(n_1722),
.B(n_1718),
.C(n_1714),
.Y(n_1733)
);

NAND4xp25_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1719),
.C(n_1729),
.D(n_1728),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1718),
.C(n_1707),
.D(n_1715),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1726),
.Y(n_1736)
);

AOI221x1_ASAP7_75t_SL g1737 ( 
.A1(n_1723),
.A2(n_1711),
.B1(n_1710),
.B2(n_1721),
.C(n_1668),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1732),
.Y(n_1739)
);

AOI31xp33_ASAP7_75t_SL g1740 ( 
.A1(n_1727),
.A2(n_1660),
.A3(n_1671),
.B(n_1661),
.Y(n_1740)
);

INVxp33_ASAP7_75t_L g1741 ( 
.A(n_1730),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1729),
.B(n_1712),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1722),
.B(n_1709),
.Y(n_1743)
);

AOI221x1_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1713),
.B1(n_1663),
.B2(n_1670),
.C(n_1668),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1741),
.B(n_1738),
.C(n_1742),
.Y(n_1745)
);

AOI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1740),
.A2(n_1734),
.B(n_1735),
.C(n_1743),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1670),
.B(n_1663),
.C(n_1642),
.Y(n_1747)
);

AND3x2_ASAP7_75t_L g1748 ( 
.A(n_1736),
.B(n_1655),
.C(n_1643),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1733),
.A2(n_1662),
.B1(n_1643),
.B2(n_1661),
.C(n_1655),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_L g1750 ( 
.A(n_1734),
.B(n_1662),
.C(n_1643),
.D(n_1661),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1746),
.A2(n_1749),
.B1(n_1745),
.B2(n_1747),
.C(n_1750),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1748),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1748),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1748),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1746),
.B(n_1648),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1745),
.B(n_1648),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1746),
.A2(n_1655),
.B1(n_1662),
.B2(n_1380),
.C(n_1441),
.Y(n_1757)
);

NOR2x1_ASAP7_75t_L g1758 ( 
.A(n_1752),
.B(n_1638),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1751),
.A2(n_1640),
.B(n_1478),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1755),
.B(n_1626),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1754),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1757),
.B(n_1418),
.C(n_1475),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1756),
.B1(n_1753),
.B2(n_1626),
.C(n_1608),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1758),
.B(n_1591),
.C(n_1596),
.Y(n_1764)
);

AOI21xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1760),
.A2(n_1552),
.B(n_1630),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1763),
.A2(n_1762),
.B1(n_1759),
.B2(n_1588),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1766),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1767),
.B(n_1764),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1765),
.B1(n_1583),
.B2(n_1588),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_1591),
.B(n_1567),
.Y(n_1770)
);

AOI22x1_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1594),
.B1(n_1567),
.B2(n_1592),
.Y(n_1771)
);

XOR2xp5_ASAP7_75t_L g1772 ( 
.A(n_1770),
.B(n_1465),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1596),
.B1(n_1552),
.B2(n_1592),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1772),
.A2(n_1597),
.B(n_1630),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1773),
.B1(n_1639),
.B2(n_1562),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1775),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_R g1777 ( 
.A1(n_1776),
.A2(n_1545),
.B1(n_1588),
.B2(n_1583),
.C(n_1594),
.Y(n_1777)
);

AOI211xp5_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1440),
.B(n_1436),
.C(n_1468),
.Y(n_1778)
);


endmodule