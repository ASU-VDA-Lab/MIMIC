module fake_jpeg_26838_n_243 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_65),
.B1(n_30),
.B2(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_74),
.B1(n_40),
.B2(n_69),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_35),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_31),
.Y(n_67)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_82),
.B(n_26),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_89),
.B1(n_101),
.B2(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_87),
.Y(n_111)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_29),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_95),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_21),
.A3(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_110),
.B1(n_59),
.B2(n_75),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_18),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_18),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_71),
.Y(n_127)
);

NOR2xp67_ASAP7_75t_R g101 ( 
.A(n_68),
.B(n_44),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_42),
.B1(n_25),
.B2(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_26),
.B1(n_30),
.B2(n_40),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_48),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_50),
.C(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_50),
.A2(n_47),
.B1(n_48),
.B2(n_18),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_53),
.B1(n_69),
.B2(n_70),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_47),
.B1(n_27),
.B2(n_19),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_19),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_135),
.C(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_123),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_71),
.B(n_72),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_122),
.A2(n_19),
.B(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_130),
.B1(n_92),
.B2(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_129),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_131),
.B1(n_82),
.B2(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_27),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_47),
.B1(n_60),
.B2(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_83),
.B(n_81),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_19),
.C(n_27),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_86),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_144),
.B1(n_148),
.B2(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_141),
.B(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_91),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_79),
.C(n_103),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_159),
.C(n_135),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_109),
.B1(n_94),
.B2(n_106),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_78),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_149),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_106),
.B1(n_81),
.B2(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_16),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_161),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_111),
.B(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_117),
.B1(n_134),
.B2(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_123),
.B(n_136),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_99),
.C(n_90),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_90),
.B1(n_28),
.B2(n_99),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_169),
.B1(n_179),
.B2(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_170),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_120),
.B1(n_128),
.B2(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_171),
.A2(n_172),
.B(n_174),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_129),
.B(n_114),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_130),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_150),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_126),
.B(n_124),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_162),
.B(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_125),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_181),
.B1(n_161),
.B2(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_145),
.B1(n_140),
.B2(n_139),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_159),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_199),
.C(n_202),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_192),
.B1(n_196),
.B2(n_202),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_190),
.B(n_200),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_174),
.B(n_172),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_171),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_142),
.Y(n_193)
);

AO221x1_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_156),
.B1(n_154),
.B2(n_5),
.C(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_139),
.B(n_160),
.C(n_151),
.D(n_147),
.Y(n_198)
);

NOR4xp25_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_184),
.C(n_173),
.D(n_8),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_160),
.C(n_4),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_1),
.B(n_5),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_1),
.C(n_7),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_169),
.B1(n_178),
.B2(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_208),
.B1(n_214),
.B2(n_201),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_191),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_176),
.B1(n_183),
.B2(n_167),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_167),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_215),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_195),
.B(n_186),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_1),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_7),
.B(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_200),
.Y(n_220)
);

AOI221xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_209),
.B1(n_216),
.B2(n_207),
.C(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_199),
.C(n_188),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_194),
.C(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_194),
.C(n_198),
.Y(n_227)
);

AOI31xp67_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_232),
.A3(n_229),
.B(n_12),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_207),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_217),
.B1(n_215),
.B2(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_7),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_15),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_221),
.B(n_10),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_237),
.B(n_15),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_241)
);

OAI31xp33_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_13),
.A3(n_14),
.B(n_15),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_13),
.Y(n_243)
);


endmodule