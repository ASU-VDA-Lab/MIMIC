module real_jpeg_33364_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_50;
wire n_33;
wire n_29;
wire n_49;
wire n_52;
wire n_10;
wire n_9;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_51;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_1),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NAND2x1p5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_24),
.Y(n_23)
);

BUFx2_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_49),
.A3(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

OAI211xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_25),
.B(n_29),
.C(n_48),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_16),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

AND2x4_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_13),
.B(n_15),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_15),
.B(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_20),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_19),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B1(n_42),
.B2(n_47),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule