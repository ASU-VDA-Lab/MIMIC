module real_aes_4497_n_11 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10, n_11);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
input n_10;
output n_11;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_16;
wire n_15;
wire n_20;
wire n_18;
wire n_21;
NAND2xp33_ASAP7_75t_R g11 ( .A(n_0), .B(n_12), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_2), .B(n_5), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_3), .B(n_19), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_6), .B(n_20), .C(n_21), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g13 ( .A(n_7), .B(n_8), .C(n_14), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_9), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_10), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g12 ( .A(n_13), .B(n_15), .Y(n_12) );
NAND3xp33_ASAP7_75t_SL g15 ( .A(n_16), .B(n_17), .C(n_18), .Y(n_15) );
endmodule