module fake_netlist_5_2316_n_1495 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1495);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1495;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_SL g405 ( 
.A(n_343),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_237),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_79),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_253),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_10),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_71),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_215),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_56),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_245),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_311),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_294),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_180),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_149),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_12),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_192),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_3),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_282),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_138),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_34),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_246),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_49),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_250),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_266),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_120),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_291),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_367),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_16),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_74),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_242),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_231),
.B(n_239),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_322),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_338),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_120),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_233),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_169),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_349),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_317),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_328),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_330),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_31),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_385),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_218),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_229),
.B(n_304),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_7),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_167),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_108),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_163),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_319),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_38),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_205),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_189),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_287),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_318),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_202),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_69),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_110),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_22),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_61),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_299),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_78),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_268),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_329),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_150),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_342),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_344),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_23),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_364),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_139),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_234),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_13),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_129),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_326),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_284),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_370),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_185),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_382),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_288),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_147),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_31),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_315),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_346),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_142),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_26),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_320),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_39),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_40),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_151),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_327),
.Y(n_500)
);

BUFx5_ASAP7_75t_L g501 ( 
.A(n_310),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_388),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_243),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_372),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_83),
.B(n_94),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_261),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_391),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_305),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_14),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_96),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_92),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_226),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_355),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_274),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_30),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_356),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_104),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_16),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_270),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_362),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_79),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_11),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_152),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_201),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_232),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_337),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_3),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_321),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_144),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_182),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_183),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_136),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_187),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_137),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_95),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_316),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_117),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_114),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_8),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_81),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_339),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_105),
.B(n_267),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_75),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_324),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_313),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_124),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_260),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_395),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_380),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_347),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_140),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_240),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_286),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_157),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_277),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_314),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_280),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_35),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_301),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_331),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_217),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_285),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_247),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_203),
.B(n_279),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_195),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_109),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_265),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_248),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_34),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_196),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_48),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_211),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_399),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_351),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_361),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_6),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_325),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_105),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_340),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_249),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_373),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_333),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_177),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_307),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_209),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_336),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_257),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_225),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_402),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

AOI22x1_ASAP7_75t_SL g594 ( 
.A1(n_419),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_594)
);

OA21x2_ASAP7_75t_L g595 ( 
.A1(n_421),
.A2(n_0),
.B(n_2),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_501),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_559),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_457),
.B(n_4),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_443),
.B(n_4),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g600 ( 
.A1(n_425),
.A2(n_5),
.B(n_6),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_496),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_443),
.B(n_5),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_437),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_569),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_437),
.Y(n_606)
);

CKINVDCx6p67_ASAP7_75t_R g607 ( 
.A(n_579),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_501),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_437),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_409),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_437),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_501),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_569),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_408),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_409),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_409),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_496),
.B(n_12),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_561),
.B(n_476),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_409),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_519),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_579),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_552),
.B(n_13),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_561),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_414),
.A2(n_126),
.B(n_125),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_523),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_449),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_455),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_552),
.B(n_14),
.Y(n_635)
);

BUFx12f_ASAP7_75t_L g636 ( 
.A(n_560),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_517),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_412),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_427),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_431),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_436),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_534),
.B(n_127),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_457),
.B(n_447),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_464),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_426),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

BUFx8_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_489),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_563),
.B(n_15),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_534),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_447),
.B(n_17),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_465),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_494),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_513),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_428),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_515),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_560),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_568),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_521),
.Y(n_661)
);

CKINVDCx6p67_ASAP7_75t_R g662 ( 
.A(n_539),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_562),
.B(n_128),
.Y(n_663)
);

BUFx8_ASAP7_75t_L g664 ( 
.A(n_540),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_406),
.A2(n_131),
.B(n_130),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_499),
.B(n_18),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_417),
.B(n_132),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_616),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_643),
.B(n_474),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_610),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_614),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_610),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_465),
.C(n_545),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_624),
.B(n_507),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_604),
.B(n_424),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_635),
.B(n_474),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_617),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_624),
.B(n_407),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_617),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_632),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_620),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_598),
.B(n_434),
.C(n_410),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_620),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_604),
.B(n_429),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_659),
.B(n_660),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_642),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_619),
.B(n_405),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_642),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_SL g695 ( 
.A(n_650),
.B(n_520),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_626),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_604),
.B(n_430),
.Y(n_697)
);

INVx6_ASAP7_75t_L g698 ( 
.A(n_664),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_598),
.B(n_418),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_660),
.B(n_435),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_662),
.B(n_411),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_636),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_597),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_596),
.A2(n_438),
.B(n_432),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_604),
.B(n_441),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_667),
.B(n_418),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_648),
.Y(n_708)
);

INVx11_ASAP7_75t_L g709 ( 
.A(n_648),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_652),
.B(n_460),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_628),
.Y(n_712)
);

CKINVDCx6p67_ASAP7_75t_R g713 ( 
.A(n_659),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_444),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_618),
.B(n_458),
.C(n_453),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_593),
.B(n_535),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_606),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_669),
.B(n_466),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_630),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_656),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_609),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_652),
.B(n_451),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_692),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_699),
.B(n_707),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_699),
.B(n_656),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_707),
.B(n_711),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_672),
.B(n_664),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_688),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_674),
.B(n_646),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_672),
.A2(n_669),
.B1(n_600),
.B2(n_595),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_711),
.B(n_601),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_701),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_SL g733 ( 
.A(n_702),
.B(n_413),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_679),
.B(n_656),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_688),
.B(n_599),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_722),
.A2(n_599),
.B(n_603),
.C(n_665),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_716),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_720),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_689),
.B(n_700),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_674),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_675),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_675),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_676),
.A2(n_669),
.B1(n_600),
.B2(n_595),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_721),
.B(n_657),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_704),
.B(n_603),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_674),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_721),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_681),
.B(n_677),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_715),
.B(n_602),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_677),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_713),
.B(n_627),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_704),
.B(n_459),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_681),
.A2(n_542),
.B1(n_548),
.B2(n_547),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_712),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_695),
.A2(n_588),
.B1(n_618),
.B2(n_613),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_698),
.B(n_605),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_714),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_683),
.B(n_415),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_685),
.B(n_695),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_670),
.B(n_658),
.Y(n_760)
);

OA22x2_ASAP7_75t_L g761 ( 
.A1(n_684),
.A2(n_653),
.B1(n_623),
.B2(n_631),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_671),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_671),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_691),
.B(n_416),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_686),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_678),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_696),
.B(n_658),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_698),
.B(n_607),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_698),
.B(n_625),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_687),
.B(n_653),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_680),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_719),
.B(n_634),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_708),
.A2(n_542),
.B1(n_574),
.B2(n_524),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_682),
.B(n_661),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_697),
.B(n_639),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_691),
.B(n_420),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_691),
.B(n_693),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_690),
.B(n_694),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_718),
.A2(n_629),
.B(n_669),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_703),
.B(n_422),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_710),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_706),
.B(n_634),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_693),
.B(n_595),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_717),
.B(n_609),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_717),
.B(n_609),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_726),
.A2(n_600),
.B1(n_456),
.B2(n_463),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_724),
.A2(n_452),
.B(n_567),
.C(n_439),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_740),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_740),
.B(n_621),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_732),
.B(n_621),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_757),
.B(n_734),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_732),
.B(n_709),
.Y(n_792)
);

AND2x4_ASAP7_75t_SL g793 ( 
.A(n_768),
.B(n_454),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_747),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_748),
.A2(n_473),
.B1(n_477),
.B2(n_468),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_728),
.B(n_640),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_731),
.A2(n_736),
.B(n_750),
.C(n_770),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_759),
.A2(n_647),
.B(n_649),
.C(n_645),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_750),
.A2(n_433),
.B1(n_440),
.B2(n_423),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_723),
.A2(n_655),
.B(n_654),
.C(n_641),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_737),
.B(n_638),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_737),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_783),
.A2(n_705),
.B(n_663),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_723),
.B(n_668),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_727),
.B(n_445),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_730),
.A2(n_743),
.B1(n_783),
.B2(n_766),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_735),
.A2(n_615),
.B(n_611),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_779),
.A2(n_615),
.B(n_611),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_772),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_730),
.A2(n_480),
.B1(n_481),
.B2(n_478),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_777),
.A2(n_633),
.B(n_615),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_741),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_766),
.B(n_482),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_762),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_742),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_744),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_739),
.A2(n_785),
.B(n_784),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_778),
.A2(n_743),
.B(n_774),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_733),
.B(n_483),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_740),
.B(n_446),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_753),
.B(n_467),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_749),
.B(n_448),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_755),
.A2(n_749),
.B1(n_745),
.B2(n_756),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_775),
.A2(n_486),
.B(n_487),
.C(n_485),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_760),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_751),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_781),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_782),
.B(n_488),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_781),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_769),
.B(n_479),
.C(n_475),
.Y(n_831)
);

AO22x1_ASAP7_75t_L g832 ( 
.A1(n_746),
.A2(n_511),
.B1(n_512),
.B2(n_497),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_764),
.A2(n_663),
.B(n_642),
.Y(n_833)
);

OAI321xp33_ASAP7_75t_L g834 ( 
.A1(n_773),
.A2(n_498),
.A3(n_491),
.B1(n_504),
.B2(n_500),
.C(n_490),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_763),
.A2(n_506),
.B(n_510),
.C(n_505),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_761),
.B(n_450),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_752),
.B(n_530),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_756),
.A2(n_529),
.B1(n_532),
.B2(n_526),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_776),
.A2(n_663),
.B(n_642),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_771),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_761),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_758),
.B(n_756),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_781),
.A2(n_651),
.B(n_644),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_780),
.A2(n_651),
.B(n_644),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_729),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_729),
.A2(n_554),
.B(n_555),
.C(n_553),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_746),
.B(n_558),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_724),
.B(n_566),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_724),
.B(n_570),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_748),
.A2(n_462),
.B1(n_470),
.B2(n_461),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_731),
.B(n_541),
.C(n_538),
.Y(n_852)
);

AND2x2_ASAP7_75t_SL g853 ( 
.A(n_733),
.B(n_573),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_754),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_724),
.B(n_575),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_724),
.B(n_576),
.Y(n_856)
);

AOI21xp33_ASAP7_75t_L g857 ( 
.A1(n_726),
.A2(n_581),
.B(n_572),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_724),
.B(n_577),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_725),
.A2(n_608),
.B(n_596),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_783),
.A2(n_663),
.B(n_642),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_737),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_725),
.A2(n_612),
.B(n_608),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_724),
.B(n_578),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_738),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_726),
.A2(n_586),
.B(n_584),
.C(n_612),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_724),
.B(n_663),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_L g867 ( 
.A(n_731),
.B(n_472),
.C(n_471),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_754),
.Y(n_868)
);

AOI22x1_ASAP7_75t_L g869 ( 
.A1(n_750),
.A2(n_492),
.B1(n_493),
.B2(n_484),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_724),
.B(n_495),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_724),
.B(n_502),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_740),
.B(n_666),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_726),
.B(n_503),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_724),
.B(n_509),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_724),
.B(n_516),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_725),
.A2(n_522),
.B(n_518),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_726),
.A2(n_527),
.B1(n_531),
.B2(n_525),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_724),
.B(n_533),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_819),
.A2(n_537),
.B(n_536),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_873),
.B(n_544),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_818),
.A2(n_637),
.B(n_133),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_807),
.A2(n_550),
.B(n_549),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_795),
.B(n_637),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_791),
.A2(n_556),
.B(n_551),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_861),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_804),
.A2(n_564),
.B(n_557),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_866),
.A2(n_571),
.B(n_565),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_860),
.A2(n_582),
.B(n_580),
.Y(n_888)
);

AO31x2_ASAP7_75t_L g889 ( 
.A1(n_811),
.A2(n_21),
.A3(n_19),
.B(n_20),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_815),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_809),
.A2(n_585),
.B(n_583),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_864),
.B(n_870),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_817),
.A2(n_589),
.B(n_587),
.Y(n_893)
);

OA21x2_ASAP7_75t_L g894 ( 
.A1(n_859),
.A2(n_591),
.B(n_590),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_827),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_795),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_822),
.A2(n_592),
.B(n_594),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_826),
.A2(n_135),
.B(n_134),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_798),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_839),
.A2(n_143),
.B(n_141),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_862),
.A2(n_404),
.B(n_146),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_829),
.A2(n_148),
.B(n_145),
.Y(n_902)
);

NOR2x1_ASAP7_75t_SL g903 ( 
.A(n_788),
.B(n_153),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_878),
.A2(n_155),
.B(n_154),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_857),
.A2(n_837),
.B(n_787),
.C(n_849),
.Y(n_905)
);

OAI21x1_ASAP7_75t_SL g906 ( 
.A1(n_833),
.A2(n_158),
.B(n_156),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_841),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_810),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_795),
.B(n_159),
.Y(n_909)
);

AO31x2_ASAP7_75t_L g910 ( 
.A1(n_865),
.A2(n_25),
.A3(n_23),
.B(n_24),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_850),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_828),
.Y(n_912)
);

NOR2x1_ASAP7_75t_SL g913 ( 
.A(n_788),
.B(n_164),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_871),
.B(n_25),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_802),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_872),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_874),
.A2(n_166),
.B(n_165),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_SL g918 ( 
.A1(n_824),
.A2(n_26),
.B(n_27),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_875),
.B(n_28),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_797),
.Y(n_920)
);

OAI21x1_ASAP7_75t_SL g921 ( 
.A1(n_840),
.A2(n_170),
.B(n_168),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_846),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_855),
.A2(n_172),
.B1(n_173),
.B2(n_171),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_790),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_856),
.A2(n_863),
.B(n_858),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_L g926 ( 
.A(n_803),
.B(n_852),
.C(n_877),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_786),
.A2(n_175),
.B(n_174),
.Y(n_927)
);

CKINVDCx11_ASAP7_75t_R g928 ( 
.A(n_872),
.Y(n_928)
);

BUFx10_ASAP7_75t_L g929 ( 
.A(n_792),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_797),
.Y(n_930)
);

OA22x2_ASAP7_75t_L g931 ( 
.A1(n_842),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_820),
.A2(n_178),
.B1(n_179),
.B2(n_176),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_813),
.B(n_181),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_843),
.A2(n_33),
.B(n_29),
.C(n_32),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_805),
.B(n_814),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_794),
.A2(n_403),
.B(n_184),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_854),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_796),
.A2(n_35),
.B(n_32),
.C(n_33),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_828),
.A2(n_188),
.B(n_186),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_853),
.A2(n_191),
.B1(n_193),
.B2(n_190),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_851),
.A2(n_197),
.B1(n_198),
.B2(n_194),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_868),
.B(n_36),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_867),
.A2(n_200),
.B(n_199),
.Y(n_943)
);

OAI21xp33_ASAP7_75t_L g944 ( 
.A1(n_800),
.A2(n_36),
.B(n_37),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_834),
.B(n_37),
.C(n_38),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_SL g946 ( 
.A1(n_838),
.A2(n_39),
.B(n_40),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_SL g947 ( 
.A1(n_828),
.A2(n_830),
.B(n_788),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_808),
.A2(n_816),
.B(n_812),
.Y(n_948)
);

BUFx12f_ASAP7_75t_L g949 ( 
.A(n_848),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_789),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_830),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_793),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_41),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_836),
.Y(n_954)
);

OAI21xp33_ASAP7_75t_L g955 ( 
.A1(n_806),
.A2(n_42),
.B(n_43),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_869),
.Y(n_956)
);

AOI221x1_ASAP7_75t_L g957 ( 
.A1(n_825),
.A2(n_244),
.B1(n_400),
.B2(n_398),
.C(n_396),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_831),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_799),
.Y(n_959)
);

OAI21x1_ASAP7_75t_SL g960 ( 
.A1(n_801),
.A2(n_206),
.B(n_204),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_844),
.A2(n_208),
.B(n_207),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_847),
.A2(n_44),
.A3(n_42),
.B(n_43),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_832),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_876),
.B(n_44),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_845),
.A2(n_401),
.B(n_210),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_821),
.Y(n_966)
);

AO31x2_ASAP7_75t_L g967 ( 
.A1(n_835),
.A2(n_47),
.A3(n_45),
.B(n_46),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_861),
.B(n_45),
.Y(n_968)
);

AO31x2_ASAP7_75t_L g969 ( 
.A1(n_807),
.A2(n_50),
.A3(n_46),
.B(n_47),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_872),
.Y(n_970)
);

OAI22x1_ASAP7_75t_L g971 ( 
.A1(n_822),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_795),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_815),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_873),
.B(n_51),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_798),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_819),
.A2(n_213),
.B(n_212),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_873),
.B(n_53),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_819),
.A2(n_216),
.B(n_214),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_798),
.A2(n_220),
.B1(n_221),
.B2(n_219),
.Y(n_979)
);

OA21x2_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_223),
.B(n_222),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_819),
.A2(n_227),
.B(n_224),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_828),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_788),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_802),
.B(n_54),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_819),
.A2(n_230),
.B(n_228),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_815),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_819),
.A2(n_236),
.B(n_235),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_822),
.A2(n_55),
.B(n_56),
.Y(n_989)
);

AO31x2_ASAP7_75t_L g990 ( 
.A1(n_807),
.A2(n_55),
.A3(n_57),
.B(n_58),
.Y(n_990)
);

AO31x2_ASAP7_75t_L g991 ( 
.A1(n_807),
.A2(n_57),
.A3(n_58),
.B(n_59),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_873),
.B(n_59),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_820),
.B(n_238),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_861),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_873),
.B(n_60),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_815),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_802),
.B(n_60),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_798),
.A2(n_276),
.B1(n_393),
.B2(n_390),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_827),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_792),
.B(n_241),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_788),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_873),
.B(n_61),
.Y(n_1002)
);

BUFx2_ASAP7_75t_SL g1003 ( 
.A(n_788),
.Y(n_1003)
);

AO22x2_ASAP7_75t_L g1004 ( 
.A1(n_824),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_820),
.B(n_251),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_819),
.A2(n_254),
.B(n_252),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_795),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_873),
.A2(n_292),
.B1(n_389),
.B2(n_387),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_873),
.B(n_63),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_872),
.B(n_64),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_798),
.A2(n_290),
.B1(n_386),
.B2(n_384),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_819),
.A2(n_256),
.B(n_255),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_860),
.A2(n_259),
.B(n_258),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_873),
.B(n_65),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_861),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_820),
.B(n_262),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_807),
.A2(n_65),
.A3(n_66),
.B(n_67),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_798),
.A2(n_296),
.B1(n_383),
.B2(n_376),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_822),
.A2(n_66),
.B(n_67),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_819),
.A2(n_264),
.B(n_263),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_827),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_873),
.B(n_68),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_861),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_873),
.B(n_68),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_819),
.A2(n_271),
.B(n_269),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_792),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_896),
.B(n_972),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_994),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_892),
.A2(n_298),
.B1(n_375),
.B2(n_374),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_924),
.B(n_69),
.C(n_70),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_972),
.B(n_272),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_925),
.A2(n_297),
.B(n_371),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_937),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_930),
.B(n_273),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_948),
.A2(n_295),
.B(n_369),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_905),
.A2(n_293),
.B1(n_368),
.B2(n_366),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_881),
.A2(n_289),
.B(n_365),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_951),
.Y(n_1038)
);

INVx8_ASAP7_75t_L g1039 ( 
.A(n_970),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_915),
.B(n_70),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_974),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_1010),
.B(n_72),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_890),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_895),
.B(n_73),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_977),
.A2(n_283),
.B1(n_360),
.B2(n_359),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_992),
.A2(n_281),
.B(n_357),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_985),
.A2(n_278),
.B(n_354),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_R g1048 ( 
.A(n_949),
.B(n_74),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_928),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_935),
.B(n_75),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1007),
.B(n_275),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_1007),
.B(n_300),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_995),
.A2(n_394),
.B(n_353),
.Y(n_1053)
);

O2A1O1Ixp5_ASAP7_75t_L g1054 ( 
.A1(n_1002),
.A2(n_352),
.B(n_350),
.C(n_348),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_899),
.A2(n_76),
.A3(n_77),
.B(n_78),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_1015),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_1010),
.B(n_76),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_996),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_984),
.B(n_997),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_999),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_930),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_975),
.A2(n_80),
.A3(n_81),
.B(n_82),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_880),
.B(n_80),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1009),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_1023),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1021),
.B(n_885),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1014),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_920),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_883),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1022),
.A2(n_85),
.B(n_87),
.C(n_88),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_1024),
.B(n_87),
.C(n_88),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_897),
.B(n_89),
.C(n_90),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_916),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_883),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_SL g1075 ( 
.A1(n_927),
.A2(n_89),
.B(n_90),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_968),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_914),
.A2(n_335),
.B(n_334),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_922),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_983),
.B(n_332),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_970),
.B(n_312),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_907),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_SL g1082 ( 
.A(n_922),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_973),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_908),
.B(n_91),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_919),
.A2(n_309),
.B(n_308),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_1001),
.B(n_306),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_916),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_953),
.B(n_91),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_986),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_987),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_947),
.A2(n_303),
.B(n_302),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_936),
.A2(n_92),
.B(n_93),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_957),
.A2(n_93),
.A3(n_94),
.B(n_95),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_959),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_969),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_901),
.A2(n_96),
.B(n_97),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_926),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_942),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_882),
.A2(n_886),
.B(n_888),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_909),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_950),
.B(n_98),
.Y(n_1101)
);

CKINVDCx11_ASAP7_75t_R g1102 ( 
.A(n_929),
.Y(n_1102)
);

OAI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_918),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_963),
.B(n_102),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_L g1105 ( 
.A(n_944),
.B(n_103),
.C(n_104),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_917),
.A2(n_106),
.B(n_107),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_1003),
.B(n_106),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_879),
.A2(n_107),
.B(n_108),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_909),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_952),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_945),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_933),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_989),
.B(n_113),
.C(n_114),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_933),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_969),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_969),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_958),
.B(n_115),
.Y(n_1117)
);

BUFx8_ASAP7_75t_SL g1118 ( 
.A(n_966),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_SL g1119 ( 
.A1(n_903),
.A2(n_116),
.B(n_117),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_993),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_954),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_SL g1122 ( 
.A(n_1013),
.B(n_122),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_887),
.A2(n_123),
.B(n_906),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_954),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_956),
.A2(n_123),
.B1(n_912),
.B2(n_982),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_976),
.A2(n_981),
.B(n_1020),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1026),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_966),
.B(n_1000),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1005),
.B(n_1016),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_990),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_990),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_884),
.B(n_955),
.Y(n_1132)
);

INVx8_ASAP7_75t_L g1133 ( 
.A(n_931),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1019),
.A2(n_943),
.B(n_946),
.C(n_1006),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_893),
.B(n_964),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_971),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_934),
.B(n_1004),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_978),
.A2(n_1012),
.B(n_988),
.C(n_1011),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_965),
.A2(n_961),
.B(n_921),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1004),
.A2(n_1018),
.B1(n_979),
.B2(n_998),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_1017),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_980),
.B(n_940),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_980),
.B(n_932),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_941),
.A2(n_923),
.B1(n_911),
.B2(n_1008),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_938),
.A2(n_898),
.B1(n_900),
.B2(n_904),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_991),
.B(n_1017),
.Y(n_1146)
);

CKINVDCx16_ASAP7_75t_R g1147 ( 
.A(n_960),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_902),
.A2(n_913),
.B(n_891),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_SL g1149 ( 
.A(n_939),
.B(n_889),
.C(n_991),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1017),
.B(n_889),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_962),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_962),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_889),
.B(n_962),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_910),
.B(n_967),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_894),
.A2(n_905),
.B(n_977),
.C(n_974),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_894),
.A2(n_974),
.B1(n_992),
.B2(n_977),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_967),
.A2(n_974),
.B1(n_992),
.B2(n_977),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_974),
.A2(n_977),
.B1(n_995),
.B2(n_992),
.Y(n_1158)
);

AO21x2_ASAP7_75t_L g1159 ( 
.A1(n_985),
.A2(n_1025),
.B(n_925),
.Y(n_1159)
);

AOI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_989),
.A2(n_731),
.B1(n_672),
.B2(n_822),
.C(n_753),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_951),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_892),
.A2(n_783),
.B(n_807),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_937),
.Y(n_1163)
);

CKINVDCx12_ASAP7_75t_R g1164 ( 
.A(n_1066),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_1039),
.B(n_1133),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1081),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1100),
.B(n_1059),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1153),
.A2(n_1141),
.B(n_1154),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1094),
.B(n_1160),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1083),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1095),
.A2(n_1116),
.B(n_1115),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1083),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1118),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1089),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1039),
.B(n_1133),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1068),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1056),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1073),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1065),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1110),
.B(n_1127),
.Y(n_1180)
);

INVx4_ASAP7_75t_SL g1181 ( 
.A(n_1055),
.Y(n_1181)
);

AO21x2_ASAP7_75t_L g1182 ( 
.A1(n_1099),
.A2(n_1149),
.B(n_1159),
.Y(n_1182)
);

OAI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1111),
.A2(n_1064),
.B(n_1041),
.C(n_1075),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1033),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1088),
.B(n_1109),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1028),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1060),
.B(n_1050),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1090),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1136),
.A2(n_1113),
.B1(n_1097),
.B2(n_1105),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1031),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1073),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1076),
.B(n_1069),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1074),
.B(n_1114),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1049),
.Y(n_1194)
);

BUFx2_ASAP7_75t_SL g1195 ( 
.A(n_1110),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1121),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1163),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1043),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1058),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1112),
.B(n_1040),
.Y(n_1200)
);

AO21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1140),
.A2(n_1108),
.B(n_1137),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1104),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1102),
.Y(n_1203)
);

BUFx4f_ASAP7_75t_L g1204 ( 
.A(n_1073),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1087),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_R g1206 ( 
.A(n_1078),
.B(n_1061),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1087),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1063),
.B(n_1098),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1044),
.B(n_1128),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1027),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1084),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1038),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1117),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1095),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1152),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1115),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1124),
.B(n_1158),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1042),
.A2(n_1057),
.B1(n_1103),
.B2(n_1071),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1037),
.A2(n_1035),
.B(n_1126),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1161),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1130),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1162),
.B(n_1129),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1082),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1129),
.B(n_1061),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1138),
.A2(n_1134),
.B(n_1155),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1130),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1042),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1057),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1135),
.B(n_1157),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1080),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1131),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1131),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1107),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1031),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1132),
.B(n_1125),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1055),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1142),
.B(n_1143),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1072),
.B(n_1051),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1055),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_1156),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1146),
.B(n_1150),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1120),
.B(n_1106),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1062),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1034),
.B(n_1079),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1062),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1101),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1107),
.B(n_1070),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1052),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1067),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1046),
.A2(n_1053),
.B1(n_1036),
.B2(n_1045),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1119),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1086),
.B(n_1091),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1123),
.B(n_1148),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1030),
.B(n_1147),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1077),
.B(n_1085),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1093),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1093),
.B(n_1122),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1096),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1092),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1122),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1208),
.B(n_1032),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1242),
.B(n_1047),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1208),
.B(n_1048),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1242),
.B(n_1047),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1187),
.B(n_1029),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1204),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1166),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1169),
.B(n_1054),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1177),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1169),
.B(n_1139),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1170),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1204),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1250),
.B(n_1201),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1172),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1174),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1164),
.Y(n_1277)
);

NOR2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1190),
.B(n_1249),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1247),
.B(n_1202),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1176),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1176),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1202),
.B(n_1211),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1179),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1239),
.B(n_1184),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1196),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1217),
.B(n_1167),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1197),
.B(n_1189),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1214),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1171),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1179),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1189),
.B(n_1222),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1216),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_1215),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1196),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1186),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1253),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1185),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1229),
.B(n_1248),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1221),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1192),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1241),
.A2(n_1251),
.B(n_1219),
.Y(n_1302)
);

AO22x1_ASAP7_75t_L g1303 ( 
.A1(n_1255),
.A2(n_1203),
.B1(n_1209),
.B2(n_1224),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1213),
.B(n_1238),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1200),
.B(n_1213),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1173),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1226),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1235),
.B(n_1193),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1231),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1173),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1238),
.B(n_1188),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1168),
.B(n_1244),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1232),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1246),
.B(n_1258),
.Y(n_1315)
);

INVx11_ASAP7_75t_L g1316 ( 
.A(n_1194),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1207),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1253),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1198),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1199),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1218),
.B(n_1256),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1253),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1165),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1234),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1178),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1230),
.B(n_1210),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1212),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1249),
.B(n_1245),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1181),
.B(n_1241),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1285),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1281),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1289),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1289),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1286),
.B(n_1257),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1288),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1294),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1280),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1292),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1283),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1322),
.A2(n_1228),
.B1(n_1227),
.B2(n_1245),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1297),
.B(n_1291),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1297),
.B(n_1182),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1291),
.B(n_1182),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1279),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1296),
.B(n_1252),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1273),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1299),
.B(n_1225),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_1310),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1300),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1304),
.B(n_1305),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1307),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1322),
.B(n_1183),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1330),
.B(n_1261),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1264),
.A2(n_1165),
.B1(n_1175),
.B2(n_1195),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1330),
.B(n_1254),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1290),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1309),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1314),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1315),
.B(n_1243),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1262),
.A2(n_1183),
.B(n_1287),
.C(n_1269),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1284),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1263),
.B(n_1259),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1325),
.B(n_1220),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1263),
.B(n_1259),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1265),
.B(n_1260),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1268),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1272),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1278),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1275),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1301),
.B(n_1180),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1276),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1336),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1333),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1353),
.A2(n_1274),
.B1(n_1266),
.B2(n_1298),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1344),
.B(n_1317),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1344),
.B(n_1313),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1345),
.B(n_1351),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1346),
.B(n_1319),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1343),
.B(n_1313),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1357),
.B(n_1293),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1339),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1340),
.Y(n_1384)
);

NOR2x1_ASAP7_75t_L g1385 ( 
.A(n_1355),
.B(n_1323),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1343),
.B(n_1311),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1334),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1388)
);

BUFx2_ASAP7_75t_SL g1389 ( 
.A(n_1370),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1346),
.B(n_1323),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1364),
.B(n_1271),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1353),
.B(n_1274),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1342),
.B(n_1320),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1335),
.B(n_1282),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1350),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1362),
.B(n_1323),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1352),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1359),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1342),
.B(n_1321),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1358),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1349),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1363),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1360),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1368),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1367),
.B(n_1302),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1338),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1406),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1379),
.B(n_1337),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1375),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1377),
.B(n_1402),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1374),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1382),
.B(n_1332),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1400),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1388),
.B(n_1386),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1394),
.B(n_1332),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1393),
.B(n_1362),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1399),
.B(n_1348),
.Y(n_1417)
);

OAI33xp33_ASAP7_75t_L g1418 ( 
.A1(n_1392),
.A2(n_1331),
.A3(n_1373),
.B1(n_1371),
.B2(n_1369),
.B3(n_1365),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1396),
.A2(n_1392),
.B(n_1376),
.C(n_1385),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1381),
.B(n_1361),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1377),
.B(n_1356),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1383),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1378),
.B(n_1361),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1384),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1387),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1411),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1419),
.A2(n_1396),
.B1(n_1376),
.B2(n_1380),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1409),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1416),
.B(n_1401),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1413),
.B(n_1380),
.Y(n_1430)
);

INVxp33_ASAP7_75t_L g1431 ( 
.A(n_1407),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1422),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1425),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1410),
.B(n_1391),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1414),
.B(n_1405),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1409),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1418),
.B(n_1389),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1419),
.A2(n_1405),
.B(n_1404),
.Y(n_1438)
);

AO22x1_ASAP7_75t_L g1439 ( 
.A1(n_1424),
.A2(n_1407),
.B1(n_1306),
.B2(n_1203),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1425),
.Y(n_1440)
);

OAI21xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1417),
.A2(n_1395),
.B(n_1397),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1421),
.B(n_1391),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1429),
.B(n_1408),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1436),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1427),
.A2(n_1341),
.B1(n_1412),
.B2(n_1390),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1426),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1437),
.B(n_1420),
.Y(n_1447)
);

OAI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1438),
.A2(n_1233),
.B(n_1415),
.C(n_1372),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1437),
.B(n_1423),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1448),
.A2(n_1438),
.B(n_1429),
.C(n_1441),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1447),
.A2(n_1438),
.B1(n_1430),
.B2(n_1354),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1449),
.B(n_1442),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1445),
.Y(n_1453)
);

OAI211xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1443),
.A2(n_1233),
.B(n_1432),
.C(n_1277),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1450),
.A2(n_1439),
.B(n_1431),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1452),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1453),
.A2(n_1446),
.B(n_1431),
.C(n_1295),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1451),
.B(n_1430),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1454),
.B(n_1306),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1450),
.A2(n_1303),
.B(n_1310),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1450),
.A2(n_1370),
.B(n_1329),
.C(n_1444),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_L g1462 ( 
.A(n_1454),
.B(n_1324),
.C(n_1347),
.Y(n_1462)
);

AND2x2_ASAP7_75t_SL g1463 ( 
.A(n_1462),
.B(n_1270),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1460),
.B(n_1403),
.C(n_1398),
.Y(n_1464)
);

XNOR2xp5_ASAP7_75t_L g1465 ( 
.A(n_1455),
.B(n_1223),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1456),
.B(n_1434),
.Y(n_1466)
);

NOR3xp33_ASAP7_75t_L g1467 ( 
.A(n_1461),
.B(n_1206),
.C(n_1347),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1468)
);

NAND4xp75_ASAP7_75t_L g1469 ( 
.A(n_1459),
.B(n_1267),
.C(n_1191),
.D(n_1316),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1457),
.B(n_1440),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1466),
.B(n_1435),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1465),
.B(n_1428),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1470),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1464),
.B(n_1223),
.C(n_1273),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1463),
.B(n_1273),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1475),
.B(n_1468),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1471),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1473),
.B(n_1469),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1472),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1476),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1478),
.A2(n_1165),
.B1(n_1175),
.B2(n_1326),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1477),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1478),
.A2(n_1474),
.B1(n_1467),
.B2(n_1428),
.C(n_1346),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1482),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1480),
.B(n_1479),
.C(n_1327),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1481),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1484),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1485),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1486),
.A2(n_1483),
.B(n_1175),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1487),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1489),
.A2(n_1267),
.B(n_1205),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1490),
.A2(n_1488),
.B(n_1318),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1492),
.A2(n_1491),
.B(n_1178),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1493),
.B(n_1308),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1494),
.A2(n_1205),
.B(n_1328),
.Y(n_1495)
);


endmodule