module real_jpeg_5287_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_0),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_0),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_0),
.B(n_210),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_0),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_0),
.B(n_306),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_1),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_1),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_3),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_3),
.B(n_215),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_3),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_3),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_3),
.B(n_180),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_4),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_4),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_4),
.B(n_214),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_6),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_7),
.Y(n_513)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_8),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_8),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_8),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_9),
.B(n_93),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_9),
.B(n_109),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_9),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_9),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_9),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_9),
.B(n_415),
.Y(n_414)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_11),
.B(n_82),
.Y(n_201)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_11),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_11),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_11),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_11),
.B(n_409),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_12),
.Y(n_129)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_12),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_13),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_13),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_13),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_13),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_15),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_15),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_15),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_15),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_15),
.B(n_113),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_15),
.B(n_398),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_16),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_16),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_16),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_16),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_16),
.B(n_355),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_17),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_17),
.B(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_17),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_17),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_18),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_18),
.B(n_67),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_18),
.B(n_123),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_18),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_18),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_18),
.B(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_18),
.B(n_381),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_18),
.B(n_406),
.Y(n_405)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_508),
.B(n_511),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_159),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_158),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_98),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_25),
.B(n_98),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_75),
.B1(n_76),
.B2(n_97),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_48),
.C(n_64),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_27),
.A2(n_28),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_32),
.C(n_36),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_34),
.Y(n_221)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_35),
.Y(n_148)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_35),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.C(n_46),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_37),
.B(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_132)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_43),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_44),
.Y(n_353)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_45),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_45),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_45),
.Y(n_406)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_48),
.A2(n_64),
.B1(n_65),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_49),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_51),
.Y(n_259)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_55),
.B1(n_127),
.B2(n_130),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_151)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_55),
.B(n_122),
.C(n_127),
.Y(n_152)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_58),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_72),
.C(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_63),
.Y(n_333)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_63),
.Y(n_410)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_73),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_96),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_86),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_84),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_149),
.C(n_154),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_99),
.A2(n_100),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_131),
.C(n_133),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_101),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.C(n_121),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_102),
.A2(n_103),
.B1(n_115),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_106),
.C(n_112),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_116),
.B(n_120),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_117),
.B(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_121),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_136),
.C(n_140),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_127),
.A2(n_130),
.B1(n_140),
.B2(n_141),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_129),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_131),
.Y(n_497)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.C(n_145),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_136),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_140),
.A2(n_141),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_141),
.B(n_192),
.C(n_194),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_231)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_146),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_202),
.C(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_148),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_149),
.B(n_154),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_153),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g498 ( 
.A(n_150),
.B(n_152),
.CI(n_153),
.CON(n_498),
.SN(n_498)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_488),
.B(n_505),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_289),
.B(n_487),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_238),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_163),
.B(n_238),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_222),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_164),
.B(n_223),
.C(n_226),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_199),
.C(n_204),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_165),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.C(n_191),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_166),
.B(n_473),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_173),
.C(n_174),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_171),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_177),
.A2(n_178),
.B1(n_191),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_187),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_179),
.B(n_187),
.Y(n_463)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_182),
.B(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_191),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_196),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_197),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_204),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_216),
.C(n_218),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_205),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_213),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_206),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_213),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_215),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_216),
.B(n_218),
.Y(n_267)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_221),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_245),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_240),
.B(n_243),
.Y(n_483)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_245),
.B(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_265),
.C(n_268),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_247),
.B(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_256),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_248),
.A2(n_249),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_251),
.A2(n_252),
.B(n_255),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_251),
.B(n_256),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_431)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_262),
.B(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_263),
.B(n_366),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_268),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_280),
.C(n_285),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_270),
.B(n_465),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_277),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_271),
.B(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_273),
.A2(n_277),
.B1(n_278),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_273),
.Y(n_444)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_280),
.B(n_285),
.Y(n_465)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_481),
.B(n_486),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_468),
.B(n_480),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_450),
.B(n_467),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_424),
.B(n_449),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_392),
.B(n_423),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_358),
.B(n_391),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_335),
.B(n_357),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_313),
.B(n_334),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_310),
.B(n_312),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_308),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_308),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_315),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_323),
.B2(n_324),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_326),
.C(n_330),
.Y(n_356)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_321),
.Y(n_346)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_330),
.B2(n_331),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_356),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_347),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_346),
.C(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_343),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_377),
.C(n_378),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_354),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_361),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_375),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_376),
.C(n_379),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_365),
.C(n_368),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_371),
.B1(n_372),
.B2(n_374),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_369),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_386),
.C(n_389),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_386),
.B1(n_389),
.B2(n_390),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_383),
.Y(n_389)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_386),
.Y(n_390)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_422),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_422),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_403),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_402),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_395),
.B(n_402),
.C(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_438),
.C(n_439),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_411),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_413),
.C(n_420),
.Y(n_427)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_404),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_407),
.CI(n_408),
.CON(n_404),
.SN(n_404)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_407),
.C(n_408),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_420),
.B2(n_421),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_419),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_419),
.Y(n_434)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_447),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_447),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_436),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_428),
.C(n_436),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_433),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_459),
.C(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_441),
.C(n_446),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_445),
.B2(n_446),
.Y(n_440)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_442),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_466),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_466),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_456),
.C(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_462),
.C(n_464),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_478),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_478),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_475),
.C(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_484),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_500),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_493),
.Y(n_507)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_491),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_498),
.C(n_499),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_494),
.A2(n_495),
.B1(n_498),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_498),
.Y(n_503)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_498),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_504),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_509),
.Y(n_512)
);

INVx13_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);


endmodule