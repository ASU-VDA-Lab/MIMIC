module real_aes_1461_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g575 ( .A(n_0), .B(n_183), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_1), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g141 ( .A(n_2), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_3), .B(n_537), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g618 ( .A(n_4), .B(n_170), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_5), .B(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g611 ( .A(n_6), .Y(n_611) );
INVx1_ASAP7_75t_L g196 ( .A(n_7), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_8), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_9), .Y(n_212) );
AND2x2_ASAP7_75t_L g534 ( .A(n_10), .B(n_227), .Y(n_534) );
INVx2_ASAP7_75t_L g149 ( .A(n_11), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_12), .Y(n_113) );
INVx1_ASAP7_75t_L g184 ( .A(n_13), .Y(n_184) );
AOI221x1_ASAP7_75t_L g614 ( .A1(n_14), .A2(n_201), .B1(n_539), .B2(n_615), .C(n_617), .Y(n_614) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_15), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_16), .B(n_537), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_17), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g508 ( .A(n_17), .Y(n_508) );
INVx1_ASAP7_75t_L g181 ( .A(n_18), .Y(n_181) );
INVx1_ASAP7_75t_SL g256 ( .A(n_19), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_20), .B(n_161), .Y(n_160) );
AOI33xp33_ASAP7_75t_L g233 ( .A1(n_21), .A2(n_50), .A3(n_138), .B1(n_156), .B2(n_234), .B3(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_22), .A2(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_23), .B(n_183), .Y(n_541) );
AOI221xp5_ASAP7_75t_SL g585 ( .A1(n_24), .A2(n_40), .B1(n_537), .B2(n_539), .C(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g205 ( .A(n_25), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_26), .A2(n_117), .B1(n_118), .B2(n_498), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_26), .Y(n_117) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_27), .A2(n_92), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g151 ( .A(n_27), .B(n_92), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_28), .B(n_186), .Y(n_602) );
INVxp67_ASAP7_75t_L g613 ( .A(n_29), .Y(n_613) );
AND2x2_ASAP7_75t_L g560 ( .A(n_30), .B(n_226), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_31), .B(n_194), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_32), .A2(n_539), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_33), .B(n_186), .Y(n_587) );
AND2x2_ASAP7_75t_L g144 ( .A(n_34), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g155 ( .A(n_34), .Y(n_155) );
AND2x2_ASAP7_75t_L g170 ( .A(n_34), .B(n_141), .Y(n_170) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_35), .B(n_111), .C(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g506 ( .A(n_35), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_36), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_37), .B(n_194), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_38), .A2(n_135), .B1(n_147), .B2(n_150), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_39), .B(n_167), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_41), .A2(n_82), .B1(n_153), .B2(n_539), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_42), .B(n_161), .Y(n_257) );
AOI22xp5_ASAP7_75t_SL g812 ( .A1(n_43), .A2(n_73), .B1(n_813), .B2(n_814), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_43), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_44), .B(n_183), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_45), .B(n_172), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_46), .B(n_161), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_47), .Y(n_146) );
AND2x2_ASAP7_75t_L g578 ( .A(n_48), .B(n_226), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_49), .B(n_226), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_51), .B(n_161), .Y(n_224) );
INVx1_ASAP7_75t_L g139 ( .A(n_52), .Y(n_139) );
INVx1_ASAP7_75t_L g163 ( .A(n_52), .Y(n_163) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_53), .B(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g225 ( .A(n_54), .B(n_226), .Y(n_225) );
AOI221xp5_ASAP7_75t_L g193 ( .A1(n_55), .A2(n_75), .B1(n_153), .B2(n_194), .C(n_195), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_56), .B(n_194), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_57), .B(n_537), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_58), .B(n_147), .Y(n_214) );
AOI21xp5_ASAP7_75t_SL g244 ( .A1(n_59), .A2(n_153), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g551 ( .A(n_60), .B(n_226), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_61), .B(n_186), .Y(n_576) );
INVx1_ASAP7_75t_L g177 ( .A(n_62), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_63), .B(n_183), .Y(n_549) );
AND2x2_ASAP7_75t_SL g603 ( .A(n_64), .B(n_227), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_65), .A2(n_539), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g223 ( .A(n_66), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_67), .B(n_186), .Y(n_542) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_68), .B(n_172), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_69), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_70), .A2(n_153), .B(n_222), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_71), .A2(n_90), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
INVx1_ASAP7_75t_L g145 ( .A(n_72), .Y(n_145) );
INVx1_ASAP7_75t_L g165 ( .A(n_72), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_73), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_74), .B(n_194), .Y(n_236) );
AND2x2_ASAP7_75t_L g258 ( .A(n_76), .B(n_201), .Y(n_258) );
INVx1_ASAP7_75t_L g178 ( .A(n_77), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_78), .A2(n_153), .B(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_79), .A2(n_153), .B(n_159), .C(n_171), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_80), .B(n_537), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_81), .A2(n_85), .B1(n_194), .B2(n_537), .Y(n_565) );
INVx1_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_84), .B(n_201), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_86), .A2(n_153), .B1(n_231), .B2(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_87), .B(n_183), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_88), .B(n_183), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_89), .A2(n_121), .B1(n_122), .B2(n_125), .Y(n_120) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_90), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_90), .B(n_128), .C(n_469), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_91), .A2(n_539), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g246 ( .A(n_93), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_94), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_95), .B(n_186), .Y(n_548) );
AND2x2_ASAP7_75t_L g237 ( .A(n_96), .B(n_201), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_97), .A2(n_203), .B(n_204), .C(n_206), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_98), .B(n_537), .Y(n_577) );
INVxp67_ASAP7_75t_L g616 ( .A(n_99), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_100), .B(n_186), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_101), .A2(n_539), .B(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g500 ( .A(n_102), .Y(n_500) );
BUFx2_ASAP7_75t_SL g826 ( .A(n_102), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_103), .B(n_161), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B(n_827), .Y(n_104) );
INVx3_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g829 ( .A(n_106), .Y(n_829) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_109), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_113), .B(n_505), .Y(n_504) );
AND2x6_ASAP7_75t_SL g526 ( .A(n_113), .B(n_506), .Y(n_526) );
OR2x6_ASAP7_75t_SL g810 ( .A(n_113), .B(n_505), .Y(n_810) );
OR2x2_ASAP7_75t_L g822 ( .A(n_113), .B(n_506), .Y(n_822) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_511), .Y(n_114) );
AOI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_499), .B1(n_509), .B2(n_510), .Y(n_115) );
INVx2_ASAP7_75t_L g498 ( .A(n_118), .Y(n_498) );
XNOR2x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_126), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_123), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_SL g520 ( .A1(n_123), .A2(n_521), .B(n_522), .Y(n_520) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_432), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_355), .Y(n_127) );
INVxp67_ASAP7_75t_L g519 ( .A(n_128), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_302), .C(n_335), .Y(n_128) );
AOI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_259), .B(n_268), .C(n_292), .Y(n_129) );
OAI21xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_188), .B(n_238), .Y(n_130) );
OR2x2_ASAP7_75t_L g312 ( .A(n_131), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g467 ( .A(n_131), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_132), .A2(n_358), .B1(n_362), .B2(n_364), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_132), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_173), .Y(n_132) );
INVx1_ASAP7_75t_L g291 ( .A(n_133), .Y(n_291) );
AND2x4_ASAP7_75t_L g308 ( .A(n_133), .B(n_289), .Y(n_308) );
INVx2_ASAP7_75t_L g330 ( .A(n_133), .Y(n_330) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_133), .Y(n_413) );
AND2x2_ASAP7_75t_L g484 ( .A(n_133), .B(n_241), .Y(n_484) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_152), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_142), .C(n_146), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g194 ( .A(n_137), .B(n_143), .Y(n_194) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
OR2x6_ASAP7_75t_L g168 ( .A(n_138), .B(n_157), .Y(n_168) );
INVxp33_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g158 ( .A(n_139), .B(n_141), .Y(n_158) );
AND2x4_ASAP7_75t_L g186 ( .A(n_139), .B(n_164), .Y(n_186) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g539 ( .A(n_144), .B(n_158), .Y(n_539) );
INVx2_ASAP7_75t_L g157 ( .A(n_145), .Y(n_157) );
AND2x6_ASAP7_75t_L g183 ( .A(n_145), .B(n_162), .Y(n_183) );
INVx4_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_147), .B(n_211), .Y(n_210) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_147), .A2(n_572), .B(n_578), .Y(n_571) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x4_ASAP7_75t_L g150 ( .A(n_149), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_149), .B(n_151), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_150), .B(n_169), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_150), .A2(n_244), .B(n_248), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_150), .A2(n_536), .B(n_538), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_150), .B(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_150), .B(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_150), .B(n_616), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_150), .B(n_179), .C(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_153), .A2(n_194), .B1(n_610), .B2(n_612), .Y(n_609) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_158), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g235 ( .A(n_156), .Y(n_235) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_166), .B(n_169), .Y(n_159) );
INVx1_ASAP7_75t_L g179 ( .A(n_161), .Y(n_179) );
AND2x4_ASAP7_75t_L g537 ( .A(n_161), .B(n_170), .Y(n_537) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_168), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_168), .A2(n_169), .B(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_168), .A2(n_169), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_168), .A2(n_169), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_168), .A2(n_169), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_169), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_169), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_169), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_169), .A2(n_575), .B(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_169), .A2(n_587), .B(n_588), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_169), .A2(n_601), .B(n_602), .Y(n_600) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_229), .B(n_237), .Y(n_228) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_171), .A2(n_229), .B(n_237), .Y(n_273) );
AOI21x1_ASAP7_75t_L g563 ( .A1(n_171), .A2(n_564), .B(n_567), .Y(n_563) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_172), .A2(n_193), .B(n_198), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_172), .A2(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g249 ( .A(n_173), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
INVx3_ASAP7_75t_L g289 ( .A(n_173), .Y(n_289) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_180), .B(n_187), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_179), .B(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B1(n_184), .B2(n_185), .Y(n_180) );
INVxp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVxp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_188), .A2(n_479), .B1(n_481), .B2(n_483), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_188), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_216), .Y(n_189) );
INVx3_ASAP7_75t_L g262 ( .A(n_190), .Y(n_262) );
AND2x2_ASAP7_75t_L g270 ( .A(n_190), .B(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_190), .Y(n_300) );
NAND2x1_ASAP7_75t_SL g494 ( .A(n_190), .B(n_261), .Y(n_494) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_199), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_192), .B(n_273), .Y(n_285) );
AND2x2_ASAP7_75t_L g298 ( .A(n_192), .B(n_199), .Y(n_298) );
AND2x4_ASAP7_75t_L g305 ( .A(n_192), .B(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_192), .Y(n_354) );
INVxp67_ASAP7_75t_L g361 ( .A(n_192), .Y(n_361) );
INVx1_ASAP7_75t_L g366 ( .A(n_192), .Y(n_366) );
INVx1_ASAP7_75t_L g215 ( .A(n_194), .Y(n_215) );
INVx1_ASAP7_75t_L g265 ( .A(n_199), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_199), .B(n_275), .Y(n_284) );
INVx2_ASAP7_75t_L g352 ( .A(n_199), .Y(n_352) );
INVx1_ASAP7_75t_L g391 ( .A(n_199), .Y(n_391) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B1(n_207), .B2(n_208), .Y(n_200) );
INVx3_ASAP7_75t_L g208 ( .A(n_201), .Y(n_208) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_225), .Y(n_218) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_208), .A2(n_219), .B(n_225), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_213), .B1(n_214), .B2(n_215), .Y(n_209) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g321 ( .A(n_216), .B(n_298), .Y(n_321) );
AND2x2_ASAP7_75t_L g389 ( .A(n_216), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g403 ( .A(n_216), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_216), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_218), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g359 ( .A(n_218), .B(n_352), .Y(n_359) );
AND2x2_ASAP7_75t_L g450 ( .A(n_218), .B(n_272), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_226), .Y(n_251) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_226), .A2(n_585), .B(n_589), .Y(n_584) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
INVx2_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
AND2x2_ASAP7_75t_L g351 ( .A(n_228), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_230), .B(n_236), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
AND2x2_ASAP7_75t_L g393 ( .A(n_240), .B(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g452 ( .A(n_240), .B(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx4_ASAP7_75t_L g282 ( .A(n_241), .Y(n_282) );
AND2x4_ASAP7_75t_L g290 ( .A(n_241), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g325 ( .A(n_241), .B(n_250), .Y(n_325) );
INVx2_ASAP7_75t_L g374 ( .A(n_241), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_241), .B(n_348), .Y(n_423) );
AND2x2_ASAP7_75t_L g460 ( .A(n_241), .B(n_278), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_241), .B(n_343), .Y(n_468) );
OR2x6_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g301 ( .A(n_249), .B(n_290), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_249), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_249), .B(n_328), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_249), .B(n_341), .Y(n_462) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_250), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_250), .B(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_250), .Y(n_311) );
INVx2_ASAP7_75t_L g314 ( .A(n_250), .Y(n_314) );
INVx1_ASAP7_75t_L g347 ( .A(n_250), .Y(n_347) );
INVx1_ASAP7_75t_L g395 ( .A(n_250), .Y(n_395) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_258), .Y(n_250) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_251), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_251), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g592 ( .A1(n_251), .A2(n_554), .B(n_560), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_261), .B(n_264), .Y(n_337) );
OR2x2_ASAP7_75t_L g409 ( .A(n_261), .B(n_410), .Y(n_409) );
AND4x1_ASAP7_75t_SL g455 ( .A(n_261), .B(n_437), .C(n_456), .D(n_457), .Y(n_455) );
OR2x2_ASAP7_75t_L g479 ( .A(n_262), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g316 ( .A(n_265), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_265), .B(n_274), .Y(n_466) );
AND2x2_ASAP7_75t_L g491 ( .A(n_266), .B(n_351), .Y(n_491) );
OAI32xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_276), .A3(n_281), .B1(n_283), .B2(n_286), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g364 ( .A(n_271), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g464 ( .A(n_271), .B(n_418), .Y(n_464) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AND2x2_ASAP7_75t_L g360 ( .A(n_272), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g446 ( .A(n_272), .Y(n_446) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_273), .B(n_275), .Y(n_480) );
INVx3_ASAP7_75t_L g297 ( .A(n_274), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_274), .B(n_402), .Y(n_475) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_275), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g487 ( .A(n_277), .Y(n_487) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g327 ( .A(n_278), .Y(n_327) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_278), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_281), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_287), .Y(n_319) );
AND2x4_ASAP7_75t_L g341 ( .A(n_282), .B(n_291), .Y(n_341) );
AND2x4_ASAP7_75t_SL g412 ( .A(n_282), .B(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_282), .B(n_363), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_283), .A2(n_406), .B1(n_409), .B2(n_411), .Y(n_405) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_SL g425 ( .A(n_284), .Y(n_425) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_288), .B(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_288), .A2(n_424), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
AND2x2_ASAP7_75t_L g371 ( .A(n_289), .B(n_330), .Y(n_371) );
INVx2_ASAP7_75t_L g294 ( .A(n_290), .Y(n_294) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_299), .Y(n_292) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_296), .A2(n_368), .B1(n_372), .B2(n_373), .Y(n_367) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_297), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_297), .B(n_365), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_297), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_318), .C(n_322), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B1(n_312), .B2(n_315), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g372 ( .A(n_305), .B(n_359), .Y(n_372) );
AND2x2_ASAP7_75t_L g424 ( .A(n_305), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g441 ( .A(n_305), .B(n_391), .Y(n_441) );
AND2x2_ASAP7_75t_L g496 ( .A(n_305), .B(n_390), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx4_ASAP7_75t_L g363 ( .A(n_308), .Y(n_363) );
AND2x2_ASAP7_75t_L g373 ( .A(n_308), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g378 ( .A(n_311), .Y(n_378) );
AND2x2_ASAP7_75t_L g387 ( .A(n_311), .B(n_371), .Y(n_387) );
INVx1_ASAP7_75t_L g422 ( .A(n_313), .Y(n_422) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_316), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_317), .B(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B(n_331), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_324), .B(n_363), .Y(n_472) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AOI21xp33_ASAP7_75t_SL g335 ( .A1(n_327), .A2(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g482 ( .A(n_327), .B(n_341), .Y(n_482) );
AND2x4_ASAP7_75t_L g345 ( .A(n_328), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g379 ( .A(n_328), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_328), .B(n_395), .Y(n_461) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_344), .B(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_341), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_341), .B(n_346), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_342), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g404 ( .A(n_342), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_342), .Y(n_408) );
AND2x2_ASAP7_75t_L g492 ( .A(n_342), .B(n_460), .Y(n_492) );
AND2x2_ASAP7_75t_L g495 ( .A(n_342), .B(n_412), .Y(n_495) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_347), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g474 ( .A(n_351), .Y(n_474) );
AND2x2_ASAP7_75t_L g365 ( .A(n_352), .B(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_355), .B(n_433), .Y(n_516) );
INVxp67_ASAP7_75t_L g518 ( .A(n_355), .Y(n_518) );
NAND4xp75_ASAP7_75t_L g355 ( .A(n_356), .B(n_375), .C(n_396), .D(n_414), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_367), .Y(n_356) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_359), .B(n_446), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_360), .B(n_425), .Y(n_431) );
NAND2xp5_ASAP7_75t_R g447 ( .A(n_363), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g497 ( .A(n_363), .Y(n_497) );
INVx2_ASAP7_75t_L g410 ( .A(n_365), .Y(n_410) );
BUFx3_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g453 ( .A(n_371), .Y(n_453) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_380), .B(n_382), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_378), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_379), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_381), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_388), .B2(n_392), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_390), .A2(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g418 ( .A(n_390), .Y(n_418) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g449 ( .A(n_391), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g457 ( .A(n_391), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_392), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g427 ( .A(n_395), .B(n_428), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_403), .B(n_405), .Y(n_396) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g444 ( .A(n_401), .B(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
INVx2_ASAP7_75t_SL g448 ( .A(n_412), .Y(n_448) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_426), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B1(n_421), .B2(n_424), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_469), .Y(n_432) );
INVxp67_ASAP7_75t_L g522 ( .A(n_433), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_442), .C(n_454), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_447), .B1(n_449), .B2(n_451), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .C(n_465), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_463), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_488), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_478), .C(n_485), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_476), .B2(n_477), .Y(n_471) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g485 ( .A(n_479), .B(n_484), .C(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B1(n_493), .B2(n_495), .C1(n_496), .C2(n_497), .Y(n_488) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NOR2x1_ASAP7_75t_R g509 ( .A(n_500), .B(n_504), .Y(n_509) );
CKINVDCx14_ASAP7_75t_R g510 ( .A(n_501), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_501), .B(n_819), .C(n_823), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_815), .C(n_818), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_811), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_523), .B1(n_527), .B2(n_808), .Y(n_513) );
AO22x2_ASAP7_75t_L g817 ( .A1(n_514), .A2(n_524), .B1(n_527), .B2(n_809), .Y(n_817) );
AOI211x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .C(n_520), .Y(n_514) );
INVx4_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_738), .Y(n_528) );
NOR4xp25_ASAP7_75t_SL g529 ( .A(n_530), .B(n_631), .C(n_675), .D(n_702), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_594), .B1(n_604), .B2(n_619), .C(n_621), .Y(n_530) );
AOI32xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_561), .A3(n_568), .B1(n_579), .B2(n_590), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_532), .B(n_774), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_532), .A2(n_744), .B1(n_802), .B2(n_805), .Y(n_801) );
AND2x4_ASAP7_75t_SL g532 ( .A(n_533), .B(n_543), .Y(n_532) );
INVx5_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
OR2x2_ASAP7_75t_L g620 ( .A(n_533), .B(n_592), .Y(n_620) );
AND2x4_ASAP7_75t_L g622 ( .A(n_533), .B(n_553), .Y(n_622) );
INVx2_ASAP7_75t_L g637 ( .A(n_533), .Y(n_637) );
OR2x2_ASAP7_75t_L g649 ( .A(n_533), .B(n_562), .Y(n_649) );
AND2x2_ASAP7_75t_L g656 ( .A(n_533), .B(n_552), .Y(n_656) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_533), .B(n_581), .Y(n_698) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_533), .Y(n_755) );
OR2x6_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx3_ASAP7_75t_SL g650 ( .A(n_543), .Y(n_650) );
AND2x2_ASAP7_75t_L g669 ( .A(n_543), .B(n_593), .Y(n_669) );
AOI32xp33_ASAP7_75t_L g784 ( .A1(n_543), .A2(n_655), .A3(n_685), .B1(n_715), .B2(n_750), .Y(n_784) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_552), .Y(n_543) );
AND2x2_ASAP7_75t_L g624 ( .A(n_544), .B(n_562), .Y(n_624) );
OR2x2_ASAP7_75t_L g640 ( .A(n_544), .B(n_553), .Y(n_640) );
INVx1_ASAP7_75t_L g663 ( .A(n_544), .Y(n_663) );
INVx2_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
AND2x2_ASAP7_75t_L g716 ( .A(n_544), .B(n_581), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_544), .B(n_553), .Y(n_735) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_544), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g771 ( .A(n_553), .B(n_562), .Y(n_771) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_553), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
OR2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_561), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g638 ( .A(n_561), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g800 ( .A(n_561), .B(n_669), .Y(n_800) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g729 ( .A(n_562), .B(n_679), .Y(n_729) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_563), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_568), .B(n_696), .Y(n_798) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_569), .B(n_746), .Y(n_745) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g583 ( .A(n_570), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
AND2x2_ASAP7_75t_L g629 ( .A(n_570), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_570), .B(n_607), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_570), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
OR2x2_ASAP7_75t_L g706 ( .A(n_570), .B(n_633), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_570), .Y(n_713) );
NOR2xp33_ASAP7_75t_R g765 ( .A(n_570), .B(n_596), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_570), .B(n_608), .Y(n_769) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
AOI32xp33_ASAP7_75t_L g792 ( .A1(n_579), .A2(n_628), .A3(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
AND2x4_ASAP7_75t_L g678 ( .A(n_581), .B(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_581), .B(n_650), .Y(n_707) );
OR2x2_ASAP7_75t_L g761 ( .A(n_581), .B(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g719 ( .A(n_582), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g777 ( .A(n_582), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_583), .B(n_596), .Y(n_743) );
AND2x2_ASAP7_75t_L g780 ( .A(n_583), .B(n_746), .Y(n_780) );
INVx2_ASAP7_75t_L g630 ( .A(n_584), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_584), .B(n_596), .Y(n_653) );
INVx1_ASAP7_75t_L g684 ( .A(n_584), .Y(n_684) );
OR2x2_ASAP7_75t_L g710 ( .A(n_584), .B(n_596), .Y(n_710) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_584), .Y(n_762) );
BUFx3_ASAP7_75t_L g791 ( .A(n_584), .Y(n_791) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g660 ( .A(n_591), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_591), .B(n_678), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_591), .B(n_749), .Y(n_748) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_592), .B(n_663), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g692 ( .A1(n_592), .A2(n_659), .B(n_677), .Y(n_692) );
OAI32xp33_ASAP7_75t_L g714 ( .A1(n_593), .A2(n_715), .A3(n_717), .B1(n_719), .B2(n_721), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_593), .B(n_678), .Y(n_787) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g720 ( .A(n_595), .Y(n_720) );
NOR2x1p5_ASAP7_75t_L g790 ( .A(n_595), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g606 ( .A(n_596), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_596), .B(n_608), .Y(n_628) );
OR2x2_ASAP7_75t_L g632 ( .A(n_596), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g667 ( .A(n_596), .Y(n_667) );
AND2x2_ASAP7_75t_L g685 ( .A(n_596), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g696 ( .A(n_596), .B(n_608), .Y(n_696) );
OR2x2_ASAP7_75t_L g758 ( .A(n_596), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g775 ( .A(n_596), .B(n_706), .Y(n_775) );
INVx1_ASAP7_75t_L g807 ( .A(n_596), .Y(n_807) );
OR2x6_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_605), .B(n_684), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_606), .B(n_718), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_606), .A2(n_723), .B1(n_728), .B2(n_730), .C1(n_733), .C2(n_736), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_606), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g750 ( .A(n_606), .B(n_629), .Y(n_750) );
AND2x2_ASAP7_75t_L g712 ( .A(n_607), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g727 ( .A(n_607), .B(n_632), .Y(n_727) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_608), .B(n_633), .Y(n_665) );
AND2x4_ASAP7_75t_L g686 ( .A(n_608), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g746 ( .A(n_608), .B(n_667), .Y(n_746) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_614), .Y(n_608) );
INVx1_ASAP7_75t_SL g626 ( .A(n_620), .Y(n_626) );
NAND2xp33_ASAP7_75t_SL g795 ( .A(n_620), .B(n_650), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B(n_625), .C(n_627), .Y(n_621) );
INVx2_ASAP7_75t_SL g672 ( .A(n_622), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_623), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_624), .B(n_672), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_624), .A2(n_662), .B(n_698), .C(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g774 ( .A(n_624), .B(n_755), .Y(n_774) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x4_ASAP7_75t_L g673 ( .A(n_628), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g778 ( .A(n_628), .Y(n_778) );
OAI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_641), .C(n_668), .Y(n_631) );
INVx2_ASAP7_75t_L g643 ( .A(n_632), .Y(n_643) );
OR2x2_ASAP7_75t_L g690 ( .A(n_632), .B(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_633), .Y(n_674) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_636), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g728 ( .A(n_636), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_636), .B(n_716), .Y(n_782) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g740 ( .A1(n_638), .A2(n_741), .B1(n_742), .B2(n_744), .C1(n_747), .C2(n_750), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_639), .A2(n_704), .B1(n_707), .B2(n_708), .C(n_714), .Y(n_703) );
AND2x2_ASAP7_75t_L g741 ( .A(n_639), .B(n_698), .Y(n_741) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp33_ASAP7_75t_SL g654 ( .A(n_640), .B(n_655), .Y(n_654) );
AOI221x1_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_646), .B1(n_651), .B2(n_654), .C(n_657), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g794 ( .A(n_644), .B(n_732), .Y(n_794) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g652 ( .A(n_645), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
OAI32xp33_ASAP7_75t_L g760 ( .A1(n_650), .A2(n_691), .A3(n_761), .B1(n_763), .B2(n_767), .Y(n_760) );
OAI21xp33_ASAP7_75t_SL g779 ( .A1(n_651), .A2(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_664), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
OR2x2_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g734 ( .A(n_659), .B(n_735), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_663), .A2(n_689), .B1(n_692), .B2(n_693), .C(n_697), .Y(n_688) );
INVx1_ASAP7_75t_L g764 ( .A(n_663), .Y(n_764) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_663), .Y(n_770) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_673), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_672), .B(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_680), .B(n_688), .Y(n_675) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_679), .Y(n_749) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_682), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g701 ( .A(n_684), .Y(n_701) );
INVx1_ASAP7_75t_L g691 ( .A(n_686), .Y(n_691) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_686), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_686), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_686), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g705 ( .A(n_696), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_701), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_703), .B(n_722), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g718 ( .A(n_706), .Y(n_718) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_SL g732 ( .A(n_710), .Y(n_732) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_712), .B(n_790), .Y(n_789) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_713), .Y(n_726) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_724), .B(n_727), .Y(n_723) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g756 ( .A(n_735), .Y(n_756) );
NOR4xp25_ASAP7_75t_L g738 ( .A(n_739), .B(n_772), .C(n_783), .D(n_796), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_751), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_741), .A2(n_752), .B(n_757), .C(n_760), .Y(n_751) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_756), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g763 ( .A1(n_754), .A2(n_764), .B(n_765), .C(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
OAI21xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_770), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_SL g802 ( .A(n_771), .B(n_803), .Y(n_802) );
OAI221xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_775), .B1(n_776), .B2(n_777), .C(n_779), .Y(n_772) );
INVx1_ASAP7_75t_SL g776 ( .A(n_774), .Y(n_776) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND3xp33_ASAP7_75t_SL g783 ( .A(n_784), .B(n_785), .C(n_792), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_799), .B(n_801), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVxp33_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_811), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
BUFx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
CKINVDCx11_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
CKINVDCx8_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
endmodule