module real_aes_616_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_496;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_310;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_0), .A2(n_94), .B1(n_395), .B2(n_606), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_1), .A2(n_5), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_2), .A2(n_114), .B1(n_440), .B2(n_550), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_3), .A2(n_46), .B1(n_370), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_4), .A2(n_244), .B1(n_307), .B2(n_324), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_6), .A2(n_150), .B1(n_355), .B2(n_462), .Y(n_518) );
AO22x2_ASAP7_75t_L g314 ( .A1(n_7), .A2(n_198), .B1(n_311), .B2(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g734 ( .A(n_7), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_8), .A2(n_259), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_9), .A2(n_204), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_10), .A2(n_43), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_11), .A2(n_134), .B1(n_359), .B2(n_360), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_12), .A2(n_274), .B1(n_537), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_13), .A2(n_241), .B1(n_403), .B2(n_487), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_14), .A2(n_64), .B1(n_553), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_15), .A2(n_137), .B1(n_376), .B2(n_378), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_16), .A2(n_269), .B1(n_335), .B2(n_337), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_17), .A2(n_106), .B1(n_380), .B2(n_588), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_18), .A2(n_69), .B1(n_324), .B2(n_470), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_19), .A2(n_72), .B1(n_501), .B2(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_20), .A2(n_31), .B1(n_577), .B2(n_627), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_21), .A2(n_57), .B1(n_399), .B2(n_403), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_22), .A2(n_90), .B1(n_435), .B2(n_437), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_23), .A2(n_100), .B1(n_307), .B2(n_324), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_24), .A2(n_201), .B1(n_330), .B2(n_331), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_25), .A2(n_34), .B1(n_337), .B2(n_470), .Y(n_749) );
AO22x2_ASAP7_75t_L g310 ( .A1(n_26), .A2(n_65), .B1(n_311), .B2(n_312), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_26), .B(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_27), .A2(n_49), .B1(n_307), .B2(n_337), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_28), .A2(n_163), .B1(n_324), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_29), .A2(n_58), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_30), .A2(n_215), .B1(n_330), .B2(n_331), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_32), .A2(n_264), .B1(n_407), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_33), .A2(n_62), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_35), .A2(n_111), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_36), .A2(n_60), .B1(n_335), .B2(n_343), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g742 ( .A1(n_37), .A2(n_243), .B1(n_278), .B2(n_356), .C1(n_443), .C2(n_457), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_38), .A2(n_182), .B1(n_548), .B2(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_39), .A2(n_220), .B1(n_330), .B2(n_331), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_40), .A2(n_247), .B1(n_307), .B2(n_337), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_41), .A2(n_130), .B1(n_307), .B2(n_324), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_42), .A2(n_170), .B1(n_543), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_44), .A2(n_125), .B1(n_443), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_45), .A2(n_200), .B1(n_324), .B2(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_47), .A2(n_188), .B1(n_359), .B2(n_360), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_48), .A2(n_113), .B1(n_493), .B2(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_50), .B(n_457), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_51), .A2(n_283), .B1(n_351), .B2(n_352), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_52), .A2(n_223), .B1(n_542), .B2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_53), .A2(n_207), .B1(n_670), .B2(n_671), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_54), .A2(n_222), .B1(n_343), .B2(n_470), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_55), .A2(n_145), .B1(n_403), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_56), .A2(n_74), .B1(n_405), .B2(n_634), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_59), .A2(n_218), .B1(n_307), .B2(n_413), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_61), .A2(n_142), .B1(n_340), .B2(n_343), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_63), .A2(n_85), .B1(n_351), .B2(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_66), .A2(n_149), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI222xp33_ASAP7_75t_SL g495 ( .A1(n_67), .A2(n_185), .B1(n_270), .B2(n_378), .C1(n_433), .C2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_68), .A2(n_126), .B1(n_355), .B2(n_462), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_70), .A2(n_194), .B1(n_370), .B2(n_372), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_71), .A2(n_262), .B1(n_351), .B2(n_455), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_73), .A2(n_144), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_75), .A2(n_738), .B1(n_739), .B2(n_750), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_75), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_76), .A2(n_171), .B1(n_343), .B2(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_77), .A2(n_281), .B1(n_330), .B2(n_331), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_78), .A2(n_110), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx3_ASAP7_75t_L g311 ( .A(n_79), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_80), .A2(n_141), .B1(n_392), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_81), .A2(n_165), .B1(n_370), .B2(n_566), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_82), .A2(n_98), .B1(n_588), .B2(n_589), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_83), .A2(n_208), .B1(n_543), .B2(n_640), .Y(n_639) );
AO22x2_ASAP7_75t_L g706 ( .A1(n_84), .A2(n_707), .B1(n_719), .B2(n_720), .Y(n_706) );
INVx1_ASAP7_75t_L g719 ( .A(n_84), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_86), .A2(n_151), .B1(n_409), .B2(n_571), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_87), .A2(n_154), .B1(n_414), .B2(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_88), .A2(n_186), .B1(n_565), .B2(n_594), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_89), .A2(n_181), .B1(n_385), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_91), .A2(n_169), .B1(n_411), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_92), .A2(n_184), .B1(n_335), .B2(n_343), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_93), .A2(n_180), .B1(n_550), .B2(n_553), .Y(n_549) );
XOR2x2_ASAP7_75t_L g513 ( .A(n_95), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_96), .B(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_97), .A2(n_221), .B1(n_351), .B2(n_455), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_99), .A2(n_129), .B1(n_408), .B2(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g322 ( .A(n_101), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_101), .B(n_135), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_102), .A2(n_231), .B1(n_492), .B2(n_769), .Y(n_768) );
XNOR2x1_ASAP7_75t_L g527 ( .A(n_103), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_104), .A2(n_143), .B1(n_399), .B2(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g296 ( .A(n_105), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_107), .A2(n_287), .B(n_297), .C(n_736), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_108), .A2(n_237), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_109), .A2(n_282), .B1(n_343), .B2(n_425), .Y(n_466) );
XOR2x2_ASAP7_75t_L g366 ( .A(n_112), .B(n_367), .Y(n_366) );
XOR2x2_ASAP7_75t_L g652 ( .A(n_115), .B(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_116), .A2(n_203), .B1(n_258), .B2(n_385), .C1(n_638), .C2(n_642), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_117), .A2(n_133), .B1(n_337), .B2(n_425), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_118), .A2(n_147), .B1(n_477), .B2(n_479), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_119), .A2(n_132), .B1(n_324), .B2(n_492), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_120), .A2(n_263), .B1(n_504), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_121), .A2(n_229), .B1(n_571), .B2(n_572), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_122), .A2(n_148), .B1(n_603), .B2(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_123), .A2(n_159), .B1(n_411), .B2(n_414), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_124), .A2(n_277), .B1(n_370), .B2(n_548), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_127), .A2(n_666), .B1(n_682), .B2(n_683), .Y(n_665) );
INVx1_ASAP7_75t_L g683 ( .A(n_127), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_128), .A2(n_251), .B1(n_359), .B2(n_360), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_131), .A2(n_240), .B1(n_335), .B2(n_343), .Y(n_619) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_135), .A2(n_209), .B1(n_311), .B2(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_136), .B(n_457), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_138), .A2(n_206), .B1(n_385), .B2(n_439), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_139), .A2(n_235), .B1(n_385), .B2(n_439), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_140), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_146), .B(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_152), .A2(n_266), .B1(n_634), .B2(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_153), .B(n_433), .Y(n_713) );
INVx1_ASAP7_75t_L g323 ( .A(n_155), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_156), .A2(n_160), .B1(n_490), .B2(n_493), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_157), .A2(n_179), .B1(n_412), .B2(n_503), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_158), .A2(n_195), .B1(n_477), .B2(n_479), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_161), .A2(n_239), .B1(n_640), .B2(n_711), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_162), .A2(n_192), .B1(n_330), .B2(n_331), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_164), .A2(n_246), .B1(n_360), .B2(n_435), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_166), .A2(n_276), .B1(n_427), .B2(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_167), .B(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_168), .A2(n_234), .B1(n_413), .B2(n_576), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_172), .A2(n_211), .B1(n_330), .B2(n_331), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_173), .A2(n_197), .B1(n_330), .B2(n_331), .Y(n_656) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_174), .B(n_755), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_174), .Y(n_776) );
INVx1_ASAP7_75t_L g583 ( .A(n_175), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_176), .A2(n_265), .B1(n_382), .B2(n_385), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_177), .A2(n_232), .B1(n_490), .B2(n_607), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_178), .A2(n_191), .B1(n_392), .B2(n_395), .Y(n_391) );
XNOR2x1_ASAP7_75t_L g610 ( .A(n_183), .B(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_187), .A2(n_213), .B1(n_576), .B2(n_577), .Y(n_575) );
XNOR2x1_ASAP7_75t_L g473 ( .A(n_189), .B(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_189), .A2(n_474), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_189), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_190), .A2(n_224), .B1(n_359), .B2(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_193), .A2(n_267), .B1(n_359), .B2(n_460), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_196), .A2(n_268), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_199), .A2(n_254), .B1(n_382), .B2(n_484), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_202), .A2(n_261), .B1(n_405), .B2(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g471 ( .A(n_205), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_210), .A2(n_219), .B1(n_598), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_212), .A2(n_252), .B1(n_351), .B2(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_214), .B(n_346), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_216), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_217), .B(n_388), .Y(n_387) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_225), .B(n_688), .Y(n_687) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_226), .A2(n_304), .B1(n_363), .B2(n_364), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_226), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_227), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g730 ( .A(n_227), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_228), .A2(n_255), .B1(n_356), .B2(n_443), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_230), .A2(n_271), .B1(n_439), .B2(n_440), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_233), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
AND2x2_ASAP7_75t_R g752 ( .A(n_236), .B(n_730), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_238), .B(n_638), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_242), .A2(n_256), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_245), .A2(n_257), .B1(n_428), .B2(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_L g294 ( .A(n_248), .Y(n_294) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_249), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_250), .B(n_388), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_253), .A2(n_285), .B1(n_356), .B2(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_260), .A2(n_273), .B1(n_307), .B2(n_324), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_272), .B(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_275), .A2(n_280), .B1(n_355), .B2(n_356), .Y(n_354) );
XNOR2xp5_ASAP7_75t_L g623 ( .A(n_279), .B(n_624), .Y(n_623) );
OA22x2_ASAP7_75t_L g418 ( .A1(n_284), .A2(n_419), .B1(n_420), .B2(n_444), .Y(n_418) );
INVx1_ASAP7_75t_L g444 ( .A(n_284), .Y(n_444) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g775 ( .A(n_291), .B(n_293), .Y(n_775) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_292), .B(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_649), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_297) );
INVx1_ASAP7_75t_L g725 ( .A(n_298), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_509), .B1(n_510), .B2(n_648), .Y(n_298) );
INVx1_ASAP7_75t_L g648 ( .A(n_299), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_447), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_417), .B1(n_445), .B2(n_446), .Y(n_300) );
INVx1_ASAP7_75t_L g446 ( .A(n_301), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_365), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g364 ( .A(n_304), .Y(n_364) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_305), .B(n_344), .Y(n_304) );
NAND4xp25_ASAP7_75t_L g305 ( .A(n_306), .B(n_329), .C(n_334), .D(n_339), .Y(n_305) );
AND2x6_ASAP7_75t_L g307 ( .A(n_308), .B(n_316), .Y(n_307) );
AND2x2_ASAP7_75t_L g335 ( .A(n_308), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g342 ( .A(n_308), .B(n_325), .Y(n_342) );
AND2x2_ASAP7_75t_L g348 ( .A(n_308), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g394 ( .A(n_308), .B(n_316), .Y(n_394) );
AND2x4_ASAP7_75t_L g416 ( .A(n_308), .B(n_336), .Y(n_416) );
AND2x2_ASAP7_75t_L g425 ( .A(n_308), .B(n_336), .Y(n_425) );
AND2x4_ASAP7_75t_L g457 ( .A(n_308), .B(n_349), .Y(n_457) );
AND2x2_ASAP7_75t_L g470 ( .A(n_308), .B(n_325), .Y(n_470) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g328 ( .A(n_310), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_310), .B(n_314), .Y(n_333) );
AND2x4_ASAP7_75t_L g338 ( .A(n_310), .B(n_313), .Y(n_338) );
INVx2_ASAP7_75t_L g312 ( .A(n_311), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_311), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
OAI22x1_ASAP7_75t_L g320 ( .A1(n_311), .A2(n_321), .B1(n_322), .B2(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_311), .Y(n_321) );
INVxp67_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g327 ( .A(n_314), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g330 ( .A(n_316), .B(n_327), .Y(n_330) );
AND2x2_ASAP7_75t_L g355 ( .A(n_316), .B(n_338), .Y(n_355) );
AND2x4_ASAP7_75t_L g377 ( .A(n_316), .B(n_338), .Y(n_377) );
AND2x2_ASAP7_75t_L g402 ( .A(n_316), .B(n_327), .Y(n_402) );
AND2x2_ASAP7_75t_L g443 ( .A(n_316), .B(n_338), .Y(n_443) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx2_ASAP7_75t_L g326 ( .A(n_317), .Y(n_326) );
BUFx2_ASAP7_75t_L g332 ( .A(n_317), .Y(n_332) );
AND2x2_ASAP7_75t_L g349 ( .A(n_317), .B(n_320), .Y(n_349) );
AND2x4_ASAP7_75t_L g325 ( .A(n_319), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g336 ( .A(n_320), .B(n_326), .Y(n_336) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_320), .Y(n_353) );
AND2x6_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_325), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g343 ( .A(n_325), .B(n_333), .Y(n_343) );
AND2x4_ASAP7_75t_L g397 ( .A(n_325), .B(n_327), .Y(n_397) );
AND2x4_ASAP7_75t_L g409 ( .A(n_325), .B(n_333), .Y(n_409) );
AND2x4_ASAP7_75t_L g413 ( .A(n_325), .B(n_338), .Y(n_413) );
AND2x4_ASAP7_75t_L g359 ( .A(n_327), .B(n_336), .Y(n_359) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_336), .Y(n_371) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x4_ASAP7_75t_L g405 ( .A(n_332), .B(n_333), .Y(n_405) );
AND2x2_ASAP7_75t_SL g352 ( .A(n_333), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g386 ( .A(n_333), .B(n_353), .Y(n_386) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_333), .B(n_353), .Y(n_455) );
AND2x4_ASAP7_75t_L g351 ( .A(n_336), .B(n_338), .Y(n_351) );
AND2x2_ASAP7_75t_L g384 ( .A(n_336), .B(n_338), .Y(n_384) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_340), .Y(n_407) );
INVx2_ASAP7_75t_L g604 ( .A(n_340), .Y(n_604) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_SL g430 ( .A(n_341), .Y(n_430) );
INVx2_ASAP7_75t_L g503 ( .A(n_341), .Y(n_503) );
INVx3_ASAP7_75t_L g576 ( .A(n_341), .Y(n_576) );
INVx2_ASAP7_75t_SL g627 ( .A(n_341), .Y(n_627) );
INVx2_ASAP7_75t_SL g680 ( .A(n_341), .Y(n_680) );
INVx8_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND4xp25_ASAP7_75t_SL g344 ( .A(n_345), .B(n_350), .C(n_354), .D(n_358), .Y(n_344) );
INVx4_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_SL g389 ( .A(n_347), .Y(n_389) );
INVx3_ASAP7_75t_L g433 ( .A(n_347), .Y(n_433) );
BUFx2_ASAP7_75t_L g546 ( .A(n_347), .Y(n_546) );
INVx4_ASAP7_75t_SL g560 ( .A(n_347), .Y(n_560) );
INVx3_ASAP7_75t_L g638 ( .A(n_347), .Y(n_638) );
INVx6_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_349), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g360 ( .A(n_349), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g374 ( .A(n_349), .B(n_361), .Y(n_374) );
AND2x4_ASAP7_75t_L g380 ( .A(n_349), .B(n_357), .Y(n_380) );
AND2x2_ASAP7_75t_L g460 ( .A(n_349), .B(n_361), .Y(n_460) );
AND2x2_ASAP7_75t_L g462 ( .A(n_349), .B(n_357), .Y(n_462) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_368), .B(n_390), .Y(n_367) );
NAND4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_375), .C(n_381), .D(n_387), .Y(n_368) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g436 ( .A(n_371), .Y(n_436) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_371), .Y(n_565) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g595 ( .A(n_373), .Y(n_595) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_SL g437 ( .A(n_374), .Y(n_437) );
BUFx3_ASAP7_75t_L g480 ( .A(n_374), .Y(n_480) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_374), .Y(n_548) );
INVx1_ASAP7_75t_L g567 ( .A(n_374), .Y(n_567) );
BUFx2_ASAP7_75t_L g496 ( .A(n_376), .Y(n_496) );
BUFx2_ASAP7_75t_L g588 ( .A(n_376), .Y(n_588) );
BUFx4f_ASAP7_75t_SL g670 ( .A(n_376), .Y(n_670) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g542 ( .A(n_377), .Y(n_542) );
BUFx2_ASAP7_75t_L g563 ( .A(n_377), .Y(n_563) );
BUFx2_ASAP7_75t_L g640 ( .A(n_377), .Y(n_640) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_SL g543 ( .A(n_379), .Y(n_543) );
INVx2_ASAP7_75t_L g589 ( .A(n_379), .Y(n_589) );
INVx2_ASAP7_75t_SL g671 ( .A(n_379), .Y(n_671) );
INVx2_ASAP7_75t_L g711 ( .A(n_379), .Y(n_711) );
INVx6_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx3_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
BUFx3_ASAP7_75t_L g552 ( .A(n_384), .Y(n_552) );
BUFx5_ASAP7_75t_L g642 ( .A(n_384), .Y(n_642) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g696 ( .A(n_389), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_398), .C(n_406), .D(n_410), .Y(n_390) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g574 ( .A(n_393), .Y(n_574) );
INVx2_ASAP7_75t_SL g606 ( .A(n_393), .Y(n_606) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g492 ( .A(n_394), .Y(n_492) );
BUFx2_ASAP7_75t_L g630 ( .A(n_394), .Y(n_630) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g504 ( .A(n_396), .Y(n_504) );
INVx2_ASAP7_75t_SL g533 ( .A(n_396), .Y(n_533) );
INVx2_ASAP7_75t_L g577 ( .A(n_396), .Y(n_577) );
INVx2_ASAP7_75t_L g607 ( .A(n_396), .Y(n_607) );
INVx8_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g601 ( .A(n_400), .Y(n_601) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g488 ( .A(n_401), .Y(n_488) );
INVx1_ASAP7_75t_L g761 ( .A(n_401), .Y(n_761) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx3_ASAP7_75t_L g427 ( .A(n_402), .Y(n_427) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_402), .Y(n_634) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g535 ( .A(n_404), .Y(n_535) );
INVx2_ASAP7_75t_L g675 ( .A(n_404), .Y(n_675) );
INVx5_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g428 ( .A(n_405), .Y(n_428) );
BUFx3_ASAP7_75t_L g635 ( .A(n_405), .Y(n_635) );
BUFx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g501 ( .A(n_409), .Y(n_501) );
INVx2_ASAP7_75t_L g539 ( .A(n_409), .Y(n_539) );
BUFx3_ASAP7_75t_L g572 ( .A(n_409), .Y(n_572) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_409), .Y(n_598) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g702 ( .A(n_412), .Y(n_702) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g494 ( .A(n_413), .Y(n_494) );
BUFx3_ASAP7_75t_L g678 ( .A(n_413), .Y(n_678) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_413), .Y(n_769) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
INVx2_ASAP7_75t_L g537 ( .A(n_415), .Y(n_537) );
INVx3_ASAP7_75t_L g632 ( .A(n_415), .Y(n_632) );
INVx1_ASAP7_75t_SL g704 ( .A(n_415), .Y(n_704) );
INVx6_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g571 ( .A(n_416), .Y(n_571) );
INVx1_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR2xp67_ASAP7_75t_L g420 ( .A(n_421), .B(n_431), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_426), .C(n_429), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .C(n_438), .D(n_442), .Y(n_431) );
INVx2_ASAP7_75t_SL g593 ( .A(n_435), .Y(n_593) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g478 ( .A(n_436), .Y(n_478) );
INVx2_ASAP7_75t_L g644 ( .A(n_436), .Y(n_644) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_440), .Y(n_553) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g484 ( .A(n_441), .Y(n_484) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_472), .B(n_505), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_450), .B(n_506), .Y(n_505) );
XOR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_471), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_458), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_456), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g508 ( .A(n_474), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .C(n_495), .D(n_497), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_481), .Y(n_475) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .Y(n_485) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g531 ( .A(n_494), .Y(n_531) );
INVx2_ASAP7_75t_L g628 ( .A(n_494), .Y(n_628) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_498), .B(n_502), .Y(n_497) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_580), .B2(n_581), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_525), .B1(n_578), .B2(n_579), .Y(n_512) );
INVx2_ASAP7_75t_L g578 ( .A(n_513), .Y(n_578) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
NAND4xp25_ASAP7_75t_SL g515 ( .A(n_516), .B(n_517), .C(n_518), .D(n_519), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .C(n_523), .D(n_524), .Y(n_520) );
INVx2_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
OA22x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_554), .B2(n_555), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .C(n_534), .D(n_536), .Y(n_529) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .C(n_547), .D(n_549), .Y(n_540) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_SL g693 ( .A(n_552), .Y(n_693) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_568), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .C(n_562), .D(n_564), .Y(n_558) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .C(n_573), .D(n_575), .Y(n_568) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_608), .B1(n_646), .B2(n_647), .Y(n_581) );
INVx2_ASAP7_75t_L g646 ( .A(n_582), .Y(n_646) );
XNOR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_596), .Y(n_584) );
NAND4xp25_ASAP7_75t_SL g585 ( .A(n_586), .B(n_587), .C(n_590), .D(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .C(n_602), .D(n_605), .Y(n_596) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g647 ( .A(n_608), .Y(n_647) );
OA22x2_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_622), .B1(n_623), .B2(n_645), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_610), .Y(n_645) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_614), .C(n_615), .D(n_616), .Y(n_612) );
NAND4xp25_ASAP7_75t_SL g617 ( .A(n_618), .B(n_619), .C(n_620), .D(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_625), .B(n_636), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .C(n_631), .D(n_633), .Y(n_625) );
NAND4xp25_ASAP7_75t_SL g636 ( .A(n_637), .B(n_639), .C(n_641), .D(n_643), .Y(n_636) );
INVx1_ASAP7_75t_L g726 ( .A(n_649), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_685), .B1(n_722), .B2(n_724), .Y(n_649) );
INVx2_ASAP7_75t_SL g723 ( .A(n_650), .Y(n_723) );
AO22x2_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_665), .B2(n_684), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_659), .C(n_662), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_657), .D(n_658), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g684 ( .A(n_665), .Y(n_684) );
INVx1_ASAP7_75t_L g682 ( .A(n_666), .Y(n_682) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_667), .B(n_672), .C(n_676), .D(n_681), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_SL g724 ( .A(n_685), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B1(n_705), .B2(n_721), .Y(n_685) );
INVx4_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_697), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_692), .D(n_694), .Y(n_689) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .C(n_700), .D(n_703), .Y(n_697) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g721 ( .A(n_705), .Y(n_721) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g720 ( .A(n_707), .Y(n_720) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_714), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_712), .D(n_713), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .C(n_717), .D(n_718), .Y(n_714) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_729), .B(n_732), .Y(n_772) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
OAI222xp33_ASAP7_75t_R g736 ( .A1(n_737), .A2(n_751), .B1(n_753), .B2(n_770), .C1(n_773), .C2(n_776), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .C(n_744), .Y(n_741) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .C(n_748), .D(n_749), .Y(n_745) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND4xp75_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .C(n_763), .D(n_766), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx6p67_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
endmodule