module fake_netlist_6_784_n_1841 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1841);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1841;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_46),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_32),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_32),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_76),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_30),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_84),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_39),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_71),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_116),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_98),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_51),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_29),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_33),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_119),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_83),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_165),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_56),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_27),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_80),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_105),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_52),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_156),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_89),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_20),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_30),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_111),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_13),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_24),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_150),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_110),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_69),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_40),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_55),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_60),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_141),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_53),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_87),
.Y(n_268)
);

BUFx8_ASAP7_75t_SL g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_97),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_57),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_46),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_106),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_74),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_61),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_168),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_65),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_67),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_57),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_14),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_11),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_50),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_130),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_96),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_129),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_17),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_115),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_59),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_55),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_77),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_164),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_128),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_134),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_47),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_2),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_149),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_53),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_60),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_16),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_6),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_37),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_33),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_104),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_155),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_37),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_28),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_45),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_152),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_86),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_120),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_138),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_11),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_36),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_9),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_127),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_28),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_21),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_68),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_117),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_9),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_20),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_58),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_26),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_269),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_190),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_169),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_267),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_176),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_267),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_175),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_175),
.B(n_0),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_249),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_229),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_185),
.B(n_0),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_328),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_291),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_171),
.B(n_1),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_171),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_217),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_232),
.B(n_3),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_300),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_250),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_191),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_182),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_174),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_174),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_178),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_288),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_178),
.B(n_5),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_191),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_209),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_209),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_183),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_195),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_211),
.B(n_5),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_172),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_211),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_298),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_200),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_214),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_202),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_205),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_206),
.B(n_166),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_214),
.B(n_6),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_215),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_207),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_208),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_221),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_170),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_232),
.B(n_7),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_221),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_249),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_225),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_225),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_212),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_233),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_216),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_268),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_172),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_245),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_327),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_173),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_219),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_220),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_249),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_245),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_203),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_184),
.B(n_7),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_226),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_227),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_228),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_414),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_351),
.B(n_179),
.Y(n_420)
);

OA22x2_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_272),
.B1(n_329),
.B2(n_251),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_414),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_192),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_184),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_382),
.B(n_391),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_344),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_344),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_346),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_347),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_192),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_363),
.B(n_235),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_213),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_396),
.B(n_179),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_369),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_373),
.B(n_186),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_373),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_349),
.B(n_374),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_374),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_377),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_238),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_405),
.B(n_240),
.Y(n_487)
);

XNOR2x2_ASAP7_75t_R g488 ( 
.A(n_356),
.B(n_8),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_399),
.B(n_186),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_400),
.B(n_241),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_447),
.B(n_342),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

CKINVDCx6p67_ASAP7_75t_R g495 ( 
.A(n_475),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_187),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_395),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_345),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_422),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_431),
.A2(n_379),
.B(n_372),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_468),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_470),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_429),
.B(n_409),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_487),
.B(n_348),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_367),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_464),
.B(n_378),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_445),
.B(n_385),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_487),
.B(n_386),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_429),
.B(n_390),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_401),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_469),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_448),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_468),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_468),
.B(n_404),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

AND3x4_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_379),
.C(n_372),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_480),
.B(n_416),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_456),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_468),
.B(n_417),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_462),
.A2(n_356),
.B1(n_333),
.B2(n_358),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_473),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_468),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_402),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_420),
.B(n_383),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_472),
.B(n_418),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_448),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_435),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_426),
.A2(n_339),
.B1(n_251),
.B2(n_254),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_425),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_472),
.B(n_426),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_420),
.B(n_393),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_425),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_480),
.B(n_371),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_461),
.B(n_402),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_197),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_462),
.A2(n_260),
.B1(n_371),
.B2(n_375),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_465),
.B(n_314),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_465),
.B(n_461),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_423),
.Y(n_560)
);

NOR2x1p5_ASAP7_75t_L g561 ( 
.A(n_491),
.B(n_338),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_410),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_437),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_465),
.B(n_441),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_435),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_480),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_490),
.B(n_187),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_421),
.A2(n_276),
.B1(n_272),
.B2(n_329),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_438),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_421),
.B(n_189),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_480),
.B(n_375),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_439),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_476),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_419),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_441),
.B(n_242),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_419),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_425),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_441),
.B(n_247),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_421),
.B(n_189),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_475),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_462),
.A2(n_302),
.B1(n_243),
.B2(n_239),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_477),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_478),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_478),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_490),
.B(n_403),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_439),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_423),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_430),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_440),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_441),
.B(n_257),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_479),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_421),
.A2(n_276),
.B1(n_292),
.B2(n_271),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_441),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_423),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_441),
.B(n_261),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_480),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_480),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_490),
.B(n_403),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_419),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_421),
.A2(n_446),
.B1(n_283),
.B2(n_188),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_419),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_428),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_428),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_436),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_430),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_467),
.B(n_411),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_428),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_492),
.B(n_407),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_428),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_435),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_456),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_492),
.B(n_352),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_440),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_428),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_446),
.B(n_387),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_492),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_419),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_446),
.B(n_362),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_435),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_440),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_442),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_446),
.A2(n_442),
.B1(n_458),
.B2(n_459),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_433),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_459),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_444),
.B(n_407),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_446),
.B(n_265),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_520),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_580),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_559),
.A2(n_463),
.B(n_484),
.C(n_446),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_541),
.B(n_456),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_518),
.B(n_456),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_548),
.B(n_456),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_497),
.B(n_196),
.C(n_181),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_506),
.B(n_408),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_520),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_515),
.B(n_341),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_475),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_359),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_564),
.B(n_457),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_457),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_562),
.B(n_364),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_595),
.B(n_457),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_521),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_636),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_198),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_595),
.B(n_457),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_201),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_576),
.A2(n_266),
.B1(n_213),
.B2(n_234),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_484),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_527),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_611),
.B(n_457),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_611),
.B(n_457),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_504),
.B(n_457),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_504),
.B(n_203),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_583),
.B(n_457),
.Y(n_672)
);

INVx8_ASAP7_75t_L g673 ( 
.A(n_604),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_614),
.B(n_532),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_532),
.B(n_466),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_576),
.A2(n_234),
.B1(n_282),
.B2(n_275),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_534),
.B(n_536),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_534),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_525),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_545),
.B(n_466),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_636),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_545),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_539),
.B(n_454),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_618),
.B(n_508),
.Y(n_687)
);

BUFx6f_ASAP7_75t_SL g688 ( 
.A(n_576),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_555),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_560),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_539),
.B(n_454),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_639),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_575),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_509),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_527),
.B(n_203),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_576),
.A2(n_586),
.B1(n_570),
.B2(n_613),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_575),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_466),
.Y(n_699)
);

NAND2x1p5_ASAP7_75t_L g700 ( 
.A(n_568),
.B(n_193),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_579),
.B(n_466),
.Y(n_701)
);

BUFx6f_ASAP7_75t_SL g702 ( 
.A(n_576),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_517),
.B(n_218),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_193),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_527),
.B(n_203),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_632),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_586),
.A2(n_282),
.B1(n_252),
.B2(n_266),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_581),
.B(n_466),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_639),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_640),
.Y(n_710)
);

INVxp33_ASAP7_75t_SL g711 ( 
.A(n_505),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_581),
.B(n_466),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_598),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_466),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_580),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_591),
.B(n_466),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_592),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_586),
.A2(n_252),
.B1(n_275),
.B2(n_489),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_586),
.A2(n_489),
.B1(n_471),
.B2(n_481),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_471),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_640),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_530),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_550),
.A2(n_318),
.B1(n_319),
.B2(n_279),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_593),
.B(n_471),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_527),
.B(n_203),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_509),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_503),
.A2(n_433),
.B(n_224),
.C(n_320),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_537),
.B(n_237),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_613),
.A2(n_280),
.B1(n_281),
.B2(n_259),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_593),
.B(n_594),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_641),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_572),
.A2(n_303),
.B1(n_301),
.B2(n_312),
.C(n_311),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_594),
.B(n_471),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_596),
.B(n_471),
.Y(n_734)
);

BUFx12f_ASAP7_75t_SL g735 ( 
.A(n_586),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_596),
.B(n_471),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_537),
.B(n_237),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_602),
.B(n_471),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_554),
.A2(n_304),
.B1(n_259),
.B2(n_256),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_543),
.B(n_222),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_471),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_537),
.B(n_237),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_543),
.B(n_523),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_553),
.B(n_570),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_537),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_606),
.B(n_481),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_526),
.B(n_237),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_568),
.B(n_237),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_493),
.B(n_231),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_641),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_622),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_622),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_557),
.B(n_236),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_533),
.B(n_255),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_606),
.B(n_481),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_609),
.B(n_481),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_570),
.A2(n_489),
.B1(n_481),
.B2(n_482),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_540),
.A2(n_273),
.B1(n_274),
.B2(n_297),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_509),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_498),
.B(n_244),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_612),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_496),
.B(n_194),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_642),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_612),
.B(n_255),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_609),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_630),
.B(n_481),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_570),
.B(n_642),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_630),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_612),
.B(n_255),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_496),
.B(n_481),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_502),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_510),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_511),
.B(n_246),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_496),
.B(n_481),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_512),
.B(n_248),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_502),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_509),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_510),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_629),
.A2(n_313),
.B1(n_331),
.B2(n_299),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_631),
.B(n_255),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_631),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_507),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_631),
.B(n_255),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_513),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_605),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_582),
.A2(n_256),
.B1(n_304),
.B2(n_230),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_507),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_496),
.B(n_585),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_634),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_601),
.B(n_482),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_607),
.B(n_482),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_643),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_634),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_626),
.B(n_482),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_587),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_513),
.B(n_482),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_514),
.B(n_482),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_556),
.B(n_258),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_514),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_516),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_620),
.B(n_284),
.C(n_307),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_590),
.B(n_262),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_516),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_501),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_608),
.B(n_424),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_608),
.B(n_610),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_531),
.B(n_482),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_610),
.A2(n_230),
.B1(n_224),
.B2(n_223),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_635),
.B(n_482),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_531),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_546),
.B(n_413),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_563),
.B(n_565),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_635),
.B(n_489),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_563),
.B(n_489),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_565),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_667),
.A2(n_599),
.B(n_574),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_729),
.A2(n_529),
.B(n_577),
.C(n_552),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_697),
.B(n_616),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_667),
.B(n_616),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_667),
.A2(n_599),
.B(n_574),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_745),
.A2(n_599),
.B(n_574),
.Y(n_821)
);

BUFx4f_ASAP7_75t_L g822 ( 
.A(n_654),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_745),
.A2(n_599),
.B(n_574),
.Y(n_823)
);

AO21x1_ASAP7_75t_L g824 ( 
.A1(n_747),
.A2(n_199),
.B(n_194),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_753),
.B(n_603),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_561),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_652),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_739),
.A2(n_567),
.B(n_569),
.C(n_571),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_767),
.B(n_567),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_660),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_745),
.A2(n_619),
.B(n_604),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_660),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_767),
.B(n_569),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_706),
.B(n_528),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_744),
.B(n_571),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_656),
.A2(n_619),
.B(n_604),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_696),
.A2(n_503),
.B(n_573),
.Y(n_839)
);

OR2x2_ASAP7_75t_SL g840 ( 
.A(n_654),
.B(n_528),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_713),
.Y(n_841)
);

NAND2x1_ASAP7_75t_L g842 ( 
.A(n_677),
.B(n_619),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_647),
.A2(n_619),
.B(n_604),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_792),
.B(n_616),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_649),
.A2(n_621),
.B(n_617),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_792),
.B(n_666),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_648),
.A2(n_788),
.B(n_790),
.Y(n_847)
);

AO21x1_ASAP7_75t_L g848 ( 
.A1(n_747),
.A2(n_204),
.B(n_199),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_732),
.A2(n_597),
.B(n_573),
.C(n_627),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_791),
.A2(n_538),
.B(n_530),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_722),
.A2(n_538),
.B(n_530),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_715),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_657),
.A2(n_621),
.B(n_617),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_696),
.A2(n_725),
.B(n_705),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_706),
.B(n_528),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_680),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_659),
.A2(n_621),
.B(n_617),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_743),
.B(n_535),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_744),
.B(n_578),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_705),
.A2(n_538),
.B(n_530),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_760),
.B(n_578),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_773),
.B(n_588),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_715),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_751),
.A2(n_600),
.B(n_588),
.C(n_597),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_653),
.B(n_535),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_725),
.A2(n_737),
.B(n_728),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_681),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_775),
.B(n_600),
.Y(n_869)
);

O2A1O1Ixp5_ASAP7_75t_L g870 ( 
.A1(n_754),
.A2(n_627),
.B(n_623),
.C(n_628),
.Y(n_870)
);

NOR3xp33_ASAP7_75t_L g871 ( 
.A(n_658),
.B(n_294),
.C(n_210),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_802),
.B(n_264),
.C(n_263),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_686),
.B(n_623),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_686),
.B(n_691),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_798),
.B(n_278),
.C(n_277),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_728),
.A2(n_615),
.B(n_538),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_690),
.B(n_785),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_666),
.B(n_623),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_754),
.A2(n_638),
.B(n_628),
.C(n_499),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_663),
.A2(n_669),
.B(n_668),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_740),
.A2(n_305),
.B(n_285),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_737),
.A2(n_530),
.B(n_538),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_688),
.A2(n_561),
.B1(n_210),
.B2(n_223),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_655),
.B(n_495),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_742),
.A2(n_615),
.B(n_530),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_770),
.A2(n_633),
.B(n_522),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_742),
.A2(n_615),
.B(n_538),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_670),
.A2(n_615),
.B(n_625),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_804),
.B(n_495),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_727),
.A2(n_638),
.B(n_628),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_748),
.A2(n_615),
.B(n_625),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_687),
.B(n_638),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_795),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_662),
.B(n_253),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_685),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_752),
.A2(n_271),
.B(n_254),
.C(n_323),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_748),
.A2(n_615),
.B(n_625),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_735),
.B(n_286),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_691),
.B(n_522),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_672),
.A2(n_625),
.B(n_633),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_646),
.A2(n_812),
.B(n_774),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_674),
.A2(n_625),
.B(n_633),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_685),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_763),
.B(n_413),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_735),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_689),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_688),
.Y(n_907)
);

AO21x1_ASAP7_75t_L g908 ( 
.A1(n_808),
.A2(n_204),
.B(n_330),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_677),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_664),
.B(n_444),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_679),
.A2(n_547),
.B(n_500),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_794),
.A2(n_625),
.B(n_633),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_703),
.A2(n_323),
.B(n_322),
.C(n_292),
.Y(n_914)
);

BUFx8_ASAP7_75t_L g915 ( 
.A(n_688),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_661),
.B(n_287),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_749),
.A2(n_693),
.B(n_709),
.C(n_684),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_702),
.A2(n_666),
.B1(n_762),
.B2(n_704),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_689),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_730),
.A2(n_683),
.B(n_675),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_758),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_710),
.B(n_522),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_645),
.A2(n_624),
.B(n_522),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_702),
.A2(n_330),
.B1(n_280),
.B2(n_281),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_645),
.A2(n_761),
.B(n_678),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_692),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_721),
.B(n_293),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_699),
.A2(n_542),
.B(n_584),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_711),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_692),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_786),
.A2(n_320),
.B(n_321),
.C(n_325),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_702),
.A2(n_325),
.B1(n_321),
.B2(n_290),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_731),
.B(n_544),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_694),
.A2(n_765),
.B(n_698),
.C(n_768),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_694),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_704),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_715),
.B(n_544),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_677),
.Y(n_938)
);

INVxp33_ASAP7_75t_L g939 ( 
.A(n_801),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_781),
.B(n_544),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_750),
.B(n_544),
.Y(n_941)
);

BUFx12f_ASAP7_75t_L g942 ( 
.A(n_811),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_665),
.A2(n_270),
.B1(n_289),
.B2(n_624),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_SL g944 ( 
.A(n_723),
.B(n_316),
.C(n_296),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_701),
.A2(n_499),
.B(n_584),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_645),
.A2(n_624),
.B(n_566),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_678),
.A2(n_624),
.B(n_566),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_708),
.A2(n_714),
.B(n_712),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_781),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_678),
.A2(n_566),
.B(n_524),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_789),
.A2(n_309),
.B(n_310),
.C(n_311),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_761),
.A2(n_566),
.B(n_524),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_695),
.B(n_444),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_698),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_717),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_677),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_811),
.B(n_253),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_781),
.B(n_524),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_704),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_761),
.A2(n_524),
.B(n_558),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_781),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_771),
.B(n_776),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_800),
.A2(n_524),
.B(n_558),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_762),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_782),
.B(n_489),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_787),
.B(n_489),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_793),
.B(n_489),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_682),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_800),
.B(n_494),
.Y(n_969)
);

INVx3_ASAP7_75t_SL g970 ( 
.A(n_762),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_717),
.B(n_494),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_695),
.B(n_494),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_676),
.A2(n_309),
.B(n_322),
.C(n_317),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_650),
.B(n_253),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_765),
.B(n_499),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_671),
.A2(n_524),
.B(n_558),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_700),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_768),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_772),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_779),
.B(n_451),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_671),
.A2(n_584),
.B(n_551),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_707),
.A2(n_718),
.B(n_784),
.C(n_772),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_805),
.A2(n_682),
.B(n_741),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_778),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_306),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_716),
.A2(n_720),
.B(n_724),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_764),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_682),
.B(n_500),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_726),
.B(n_759),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_700),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_682),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_778),
.B(n_500),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_810),
.B(n_315),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_805),
.A2(n_551),
.B(n_547),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_726),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_784),
.B(n_803),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_803),
.B(n_542),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_806),
.A2(n_551),
.B1(n_547),
.B2(n_542),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_673),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_815),
.B(n_454),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_796),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_797),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_719),
.B(n_430),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_999),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_911),
.B(n_673),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_866),
.A2(n_806),
.B(n_733),
.C(n_734),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_892),
.B(n_759),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_999),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_909),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_847),
.A2(n_673),
.B(n_777),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_877),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_866),
.A2(n_746),
.B(n_755),
.C(n_736),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_859),
.A2(n_766),
.B(n_738),
.C(n_756),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_871),
.A2(n_777),
.B1(n_673),
.B2(n_780),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_874),
.B(n_807),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_929),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_892),
.B(n_814),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_859),
.B(n_764),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_871),
.A2(n_783),
.B(n_780),
.C(n_769),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_884),
.B(n_769),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_909),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_999),
.B(n_809),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_942),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_841),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_880),
.A2(n_757),
.B(n_809),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_910),
.B(n_783),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_826),
.B(n_813),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_962),
.B(n_813),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_838),
.B(n_820),
.Y(n_1031)
);

AO22x1_ASAP7_75t_L g1032 ( 
.A1(n_884),
.A2(n_336),
.B1(n_335),
.B2(n_334),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_825),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_841),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_816),
.A2(n_823),
.B(n_821),
.Y(n_1035)
);

AO32x1_ASAP7_75t_L g1036 ( 
.A1(n_998),
.A2(n_317),
.A3(n_312),
.B1(n_310),
.B2(n_451),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_819),
.A2(n_432),
.B(n_430),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_827),
.A2(n_179),
.B1(n_326),
.B2(n_451),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_822),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_934),
.A2(n_486),
.B(n_485),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_939),
.B(n_324),
.Y(n_1041)
);

BUFx2_ASAP7_75t_R g1042 ( 
.A(n_970),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_822),
.Y(n_1043)
);

CKINVDCx8_ASAP7_75t_R g1044 ( 
.A(n_835),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_819),
.A2(n_432),
.B(n_430),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_925),
.A2(n_432),
.B(n_430),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_977),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_828),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_914),
.A2(n_486),
.B(n_485),
.C(n_483),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_983),
.A2(n_432),
.B(n_430),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_862),
.A2(n_432),
.B(n_485),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_835),
.B(n_326),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_959),
.B(n_486),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_432),
.B(n_485),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_855),
.B(n_894),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_869),
.A2(n_432),
.B(n_483),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_959),
.B(n_486),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_944),
.B(n_454),
.C(n_474),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_855),
.B(n_326),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_SL g1060 ( 
.A(n_904),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_833),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_936),
.B(n_483),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_921),
.A2(n_483),
.B1(n_474),
.B2(n_460),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_920),
.A2(n_432),
.B(n_460),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_918),
.B(n_474),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_914),
.A2(n_474),
.B(n_460),
.C(n_455),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_L g1067 ( 
.A(n_949),
.B(n_889),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_893),
.B(n_8),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_840),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_917),
.A2(n_460),
.B1(n_455),
.B2(n_454),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_957),
.B(n_455),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_917),
.A2(n_896),
.B(n_817),
.C(n_881),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_836),
.B(n_455),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_SL g1074 ( 
.A1(n_818),
.A2(n_846),
.B(n_1003),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_990),
.B(n_75),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_916),
.B(n_452),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_SL g1077 ( 
.A(n_909),
.B(n_453),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_SL g1078 ( 
.A1(n_924),
.A2(n_433),
.B(n_12),
.C(n_14),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_938),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_982),
.A2(n_452),
.B1(n_450),
.B2(n_449),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_988),
.A2(n_433),
.B(n_452),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_982),
.A2(n_452),
.B1(n_450),
.B2(n_449),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_875),
.B(n_450),
.C(n_449),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_850),
.A2(n_433),
.B(n_443),
.Y(n_1084)
);

AO32x2_ASAP7_75t_L g1085 ( 
.A1(n_932),
.A2(n_10),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_970),
.B(n_453),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_SL g1087 ( 
.A(n_964),
.B(n_453),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_872),
.B(n_453),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_898),
.B(n_15),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_846),
.B(n_453),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_905),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_818),
.A2(n_443),
.B(n_435),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_868),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_856),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_860),
.A2(n_443),
.B1(n_453),
.B2(n_435),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_904),
.B(n_453),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_907),
.B(n_424),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_938),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_903),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_916),
.A2(n_424),
.B(n_78),
.C(n_162),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_905),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_938),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_907),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_832),
.A2(n_435),
.B(n_453),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_873),
.A2(n_424),
.B(n_73),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_938),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_883),
.A2(n_25),
.B(n_26),
.C(n_31),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_830),
.B(n_35),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_915),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_989),
.B(n_90),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_834),
.B(n_35),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_901),
.A2(n_424),
.B(n_93),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_837),
.B(n_99),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1003),
.A2(n_38),
.B(n_41),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_956),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_898),
.B(n_107),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_927),
.B(n_108),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_927),
.B(n_42),
.C(n_43),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_956),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1001),
.B(n_424),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_985),
.B(n_81),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_985),
.B(n_112),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_926),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_980),
.A2(n_424),
.B1(n_43),
.B2(n_44),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_857),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_953),
.A2(n_424),
.B1(n_44),
.B2(n_45),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_865),
.A2(n_42),
.B(n_48),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_949),
.B(n_123),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_930),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_SL g1130 ( 
.A(n_993),
.B(n_49),
.C(n_56),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_953),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_974),
.B(n_993),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_915),
.Y(n_1133)
);

INVx6_ASAP7_75t_L g1134 ( 
.A(n_956),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_895),
.A2(n_49),
.B1(n_59),
.B2(n_62),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_956),
.B(n_72),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_934),
.A2(n_113),
.B(n_121),
.C(n_124),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_935),
.B(n_137),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1002),
.B(n_906),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_991),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_954),
.B(n_140),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_951),
.A2(n_424),
.B(n_142),
.C(n_151),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_919),
.B(n_424),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_931),
.A2(n_844),
.B(n_973),
.C(n_978),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_844),
.A2(n_973),
.B(n_922),
.C(n_941),
.Y(n_1145)
);

AND2x4_ASAP7_75t_SL g1146 ( 
.A(n_968),
.B(n_991),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_899),
.B(n_955),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_837),
.B(n_852),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_SL g1149 ( 
.A1(n_987),
.A2(n_852),
.B1(n_961),
.B2(n_864),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_854),
.A2(n_867),
.B(n_965),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_979),
.B(n_984),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_991),
.B(n_968),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_864),
.B(n_961),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_908),
.A2(n_878),
.B1(n_995),
.B2(n_943),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_996),
.B(n_969),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_948),
.B(n_986),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_913),
.B(n_845),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1132),
.B(n_995),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1005),
.B(n_991),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1089),
.A2(n_1020),
.B1(n_1055),
.B2(n_1059),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1048),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1109),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1061),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1156),
.A2(n_902),
.B(n_900),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1012),
.B(n_878),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1150),
.A2(n_1031),
.A3(n_1127),
.B(n_1082),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1035),
.A2(n_886),
.B(n_870),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1012),
.B(n_853),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_L g1169 ( 
.A1(n_1052),
.A2(n_824),
.B(n_848),
.C(n_870),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1043),
.B(n_937),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1104),
.A2(n_879),
.B(n_888),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1017),
.B(n_975),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1011),
.A2(n_851),
.B(n_897),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_L g1174 ( 
.A(n_1004),
.B(n_972),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1080),
.A2(n_891),
.A3(n_967),
.B(n_966),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1117),
.A2(n_958),
.B(n_940),
.C(n_933),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1007),
.A2(n_842),
.B(n_858),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1034),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1019),
.A2(n_912),
.B(n_994),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1040),
.A2(n_879),
.B(n_839),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1040),
.A2(n_1050),
.B(n_1046),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1027),
.A2(n_971),
.B(n_945),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1064),
.A2(n_890),
.B(n_885),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1131),
.B(n_997),
.Y(n_1184)
);

CKINVDCx11_ASAP7_75t_R g1185 ( 
.A(n_1133),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_SL g1186 ( 
.A1(n_1107),
.A2(n_849),
.B1(n_829),
.B2(n_1000),
.C(n_947),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1017),
.A2(n_928),
.B(n_940),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1094),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1038),
.B(n_861),
.C(n_876),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1098),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1034),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1041),
.B(n_958),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1092),
.A2(n_923),
.B(n_946),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1074),
.A2(n_981),
.B(n_882),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1022),
.A2(n_992),
.B1(n_887),
.B2(n_963),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_972),
.B1(n_952),
.B2(n_950),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1125),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1072),
.A2(n_960),
.B1(n_972),
.B2(n_976),
.C(n_1135),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1121),
.A2(n_972),
.B(n_1122),
.C(n_1112),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1084),
.A2(n_972),
.B(n_1037),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1130),
.A2(n_1118),
.B(n_1068),
.C(n_1135),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1155),
.A2(n_1071),
.B(n_1073),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1131),
.B(n_1028),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1005),
.B(n_1067),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1124),
.A2(n_1139),
.B1(n_1044),
.B2(n_1155),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1013),
.A2(n_1015),
.B(n_1006),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1091),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1042),
.B(n_1047),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1076),
.B(n_1147),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1073),
.A2(n_1029),
.B(n_1145),
.Y(n_1210)
);

AO22x2_ASAP7_75t_L g1211 ( 
.A1(n_1085),
.A2(n_1116),
.B1(n_1111),
.B2(n_1108),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1030),
.A2(n_1154),
.B1(n_1110),
.B2(n_1016),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1147),
.A2(n_1088),
.B(n_1077),
.Y(n_1213)
);

AND2x2_ASAP7_75t_SL g1214 ( 
.A(n_1047),
.B(n_1128),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1032),
.B(n_1078),
.C(n_1114),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1018),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1051),
.A2(n_1054),
.B(n_1056),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1110),
.A2(n_1063),
.B1(n_1126),
.B2(n_1151),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1045),
.A2(n_1081),
.B(n_1080),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1137),
.A2(n_1136),
.B(n_1100),
.C(n_1152),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1101),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1026),
.B(n_1039),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1144),
.A2(n_1103),
.B1(n_1065),
.B2(n_1021),
.C(n_1057),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1014),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1082),
.A2(n_1070),
.B(n_1024),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1090),
.A2(n_1095),
.B(n_1070),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1025),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1004),
.A2(n_1096),
.B(n_1105),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1093),
.B(n_1099),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1095),
.A2(n_1036),
.A3(n_1143),
.B(n_1120),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1004),
.A2(n_1146),
.B(n_1120),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1138),
.A2(n_1141),
.B(n_1142),
.C(n_1083),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1024),
.A2(n_1066),
.B(n_1049),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1036),
.A2(n_1123),
.A3(n_1106),
.B(n_1115),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1004),
.A2(n_1086),
.B(n_1128),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1149),
.A2(n_1005),
.B1(n_1060),
.B2(n_1134),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1148),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1148),
.A2(n_1153),
.B(n_1097),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1134),
.A2(n_1140),
.B1(n_1098),
.B2(n_1119),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1008),
.B(n_1010),
.Y(n_1241)
);

NAND3x1_ASAP7_75t_L g1242 ( 
.A(n_1085),
.B(n_1075),
.C(n_1009),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1097),
.A2(n_1087),
.B1(n_1119),
.B2(n_1023),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1008),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1079),
.A2(n_1102),
.B(n_1036),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1098),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1102),
.B(n_1106),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1010),
.A2(n_1115),
.B(n_1140),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1140),
.B(n_1085),
.C(n_1113),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1008),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1109),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1055),
.B(n_651),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1020),
.B(n_874),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1012),
.B(n_822),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1074),
.A2(n_1156),
.B(n_1072),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1035),
.A2(n_886),
.B(n_1031),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1132),
.A2(n_651),
.B(n_866),
.Y(n_1258)
);

AOI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_866),
.B1(n_651),
.B2(n_859),
.C(n_798),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1150),
.A2(n_1031),
.A3(n_917),
.B(n_1127),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1117),
.A2(n_1122),
.B(n_1121),
.C(n_917),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1132),
.A2(n_651),
.B(n_866),
.C(n_497),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1132),
.A2(n_1020),
.B(n_866),
.C(n_497),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1034),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1132),
.A2(n_1020),
.B(n_866),
.C(n_497),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1034),
.Y(n_1269)
);

AOI211xp5_ASAP7_75t_L g1270 ( 
.A1(n_1132),
.A2(n_651),
.B(n_866),
.C(n_859),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1150),
.A2(n_1031),
.A3(n_917),
.B(n_1127),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1020),
.A2(n_1132),
.B1(n_826),
.B2(n_859),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1132),
.A2(n_866),
.B1(n_651),
.B2(n_859),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1132),
.A2(n_1020),
.B(n_866),
.C(n_497),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1132),
.A2(n_1020),
.B(n_866),
.C(n_497),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1035),
.A2(n_886),
.B(n_1031),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1040),
.A2(n_1031),
.B(n_1156),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1033),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1035),
.A2(n_886),
.B(n_1031),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1132),
.A2(n_866),
.B1(n_651),
.B2(n_658),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1008),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1012),
.B(n_840),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1035),
.A2(n_886),
.B(n_1031),
.Y(n_1286)
);

AO32x2_ASAP7_75t_L g1287 ( 
.A1(n_1080),
.A2(n_1082),
.A3(n_1070),
.B1(n_1135),
.B2(n_924),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1132),
.A2(n_871),
.B1(n_1089),
.B2(n_1112),
.C(n_1031),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1109),
.Y(n_1290)
);

AND2x6_ASAP7_75t_L g1291 ( 
.A(n_1128),
.B(n_999),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1132),
.A2(n_1020),
.B(n_866),
.C(n_497),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1108),
.A2(n_827),
.B(n_1111),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1132),
.B(n_822),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1018),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1008),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1020),
.A2(n_1132),
.B1(n_826),
.B2(n_859),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1055),
.B(n_651),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1132),
.B(n_1055),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1156),
.A2(n_745),
.B(n_667),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1035),
.A2(n_886),
.B(n_1031),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1020),
.B(n_874),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1207),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1281),
.A2(n_1270),
.B1(n_1274),
.B2(n_1292),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1270),
.A2(n_1265),
.B1(n_1268),
.B2(n_1275),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1216),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1253),
.B(n_1302),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1262),
.B(n_1266),
.Y(n_1314)
);

INVx8_ASAP7_75t_L g1315 ( 
.A(n_1291),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1272),
.A2(n_1301),
.B1(n_1160),
.B2(n_1282),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1162),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1228),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1301),
.A2(n_1264),
.B1(n_1303),
.B2(n_1300),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1291),
.Y(n_1320)
);

INVx11_ASAP7_75t_L g1321 ( 
.A(n_1244),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1296),
.A2(n_1295),
.B1(n_1192),
.B2(n_1205),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1249),
.A2(n_1206),
.B1(n_1218),
.B2(n_1212),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_1307),
.B1(n_1254),
.B2(n_1256),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1190),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1291),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1190),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1254),
.A2(n_1307),
.B1(n_1256),
.B2(n_1205),
.Y(n_1328)
);

INVx3_ASAP7_75t_SL g1329 ( 
.A(n_1214),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1159),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1211),
.A2(n_1215),
.B1(n_1212),
.B2(n_1249),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1269),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1269),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1251),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1185),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1285),
.A2(n_1218),
.B1(n_1158),
.B2(n_1209),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1222),
.A2(n_1203),
.B1(n_1233),
.B2(n_1178),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1190),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1290),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1191),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1208),
.A2(n_1289),
.B1(n_1165),
.B2(n_1267),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1208),
.A2(n_1172),
.B1(n_1279),
.B2(n_1163),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1298),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1211),
.A2(n_1215),
.B1(n_1168),
.B2(n_1188),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1237),
.A2(n_1197),
.B1(n_1242),
.B2(n_1287),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1287),
.A2(n_1201),
.B1(n_1225),
.B2(n_1172),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1246),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1224),
.A2(n_1210),
.B1(n_1184),
.B2(n_1202),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1221),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1230),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1243),
.A2(n_1236),
.B1(n_1159),
.B2(n_1204),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1189),
.A2(n_1170),
.B1(n_1227),
.B2(n_1187),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1241),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1250),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1250),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1284),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1287),
.A2(n_1194),
.B1(n_1174),
.B2(n_1223),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1240),
.Y(n_1358)
);

BUFx2_ASAP7_75t_SL g1359 ( 
.A(n_1284),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1299),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1194),
.A2(n_1223),
.B1(n_1278),
.B2(n_1179),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1196),
.A2(n_1239),
.B1(n_1238),
.B2(n_1213),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1299),
.A2(n_1247),
.B1(n_1232),
.B2(n_1229),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1226),
.A2(n_1177),
.B(n_1157),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1240),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1195),
.Y(n_1366)
);

BUFx8_ASAP7_75t_L g1367 ( 
.A(n_1294),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1278),
.A2(n_1195),
.B1(n_1183),
.B2(n_1182),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1248),
.A2(n_1252),
.B1(n_1263),
.B2(n_1305),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1235),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1261),
.B(n_1271),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1183),
.A2(n_1164),
.B1(n_1234),
.B2(n_1181),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1235),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1245),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1260),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1198),
.A2(n_1219),
.B1(n_1199),
.B2(n_1180),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1276),
.A2(n_1293),
.B1(n_1304),
.B2(n_1288),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1283),
.A2(n_1297),
.B1(n_1173),
.B2(n_1217),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1198),
.A2(n_1166),
.B1(n_1200),
.B2(n_1171),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1193),
.A2(n_1167),
.B1(n_1306),
.B2(n_1286),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1220),
.A2(n_1176),
.B1(n_1186),
.B2(n_1169),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1280),
.A2(n_1257),
.B1(n_1277),
.B2(n_1186),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1166),
.A2(n_1272),
.B1(n_1301),
.B2(n_866),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1166),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1231),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1175),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1231),
.A2(n_1259),
.B1(n_1273),
.B2(n_1258),
.Y(n_1387)
);

BUFx8_ASAP7_75t_L g1388 ( 
.A(n_1231),
.Y(n_1388)
);

INVx6_ASAP7_75t_L g1389 ( 
.A(n_1244),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1216),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1162),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1161),
.Y(n_1392)
);

CKINVDCx12_ASAP7_75t_R g1393 ( 
.A(n_1222),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1255),
.B(n_1069),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1161),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1281),
.A2(n_1270),
.B1(n_1265),
.B2(n_1268),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1281),
.A2(n_1259),
.B(n_866),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1281),
.A2(n_1273),
.B1(n_1259),
.B2(n_1272),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1281),
.A2(n_1270),
.B1(n_1265),
.B2(n_1268),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1244),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_866),
.B1(n_1273),
.B2(n_1281),
.Y(n_1405)
);

BUFx2_ASAP7_75t_SL g1406 ( 
.A(n_1228),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1259),
.A2(n_866),
.B1(n_1273),
.B2(n_1281),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1281),
.A2(n_1259),
.B(n_866),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1272),
.A2(n_1301),
.B1(n_866),
.B2(n_1253),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1162),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1207),
.Y(n_1412)
);

INVx4_ASAP7_75t_SL g1413 ( 
.A(n_1291),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1281),
.A2(n_1270),
.B1(n_1265),
.B2(n_1268),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1161),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1161),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1161),
.Y(n_1418)
);

BUFx4_ASAP7_75t_R g1419 ( 
.A(n_1208),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1244),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1255),
.B(n_1069),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1161),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1244),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1185),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1258),
.B2(n_1272),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1388),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1375),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1378),
.A2(n_1364),
.B(n_1377),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1330),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1386),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1369),
.A2(n_1380),
.B(n_1382),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1318),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1374),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1340),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1388),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1384),
.Y(n_1436)
);

AOI21xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1399),
.A2(n_1408),
.B(n_1398),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1371),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1384),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1370),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1373),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1313),
.B(n_1314),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1344),
.B(n_1331),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1346),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1346),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1365),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1383),
.B(n_1344),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1399),
.A2(n_1410),
.B1(n_1407),
.B2(n_1405),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1410),
.A2(n_1403),
.B(n_1308),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1330),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1392),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1357),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1395),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1382),
.A2(n_1380),
.B(n_1372),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1357),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1372),
.A2(n_1368),
.B(n_1381),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1362),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1415),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1310),
.A2(n_1396),
.B1(n_1401),
.B2(n_1414),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1417),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1406),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1331),
.B(n_1311),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1368),
.A2(n_1363),
.B(n_1348),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1418),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1332),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1385),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1348),
.A2(n_1352),
.B(n_1351),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1336),
.B(n_1316),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1333),
.Y(n_1469)
);

CKINVDCx6p67_ASAP7_75t_R g1470 ( 
.A(n_1335),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1393),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1309),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1315),
.B(n_1330),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1383),
.B(n_1323),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1379),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1379),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1323),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1326),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1352),
.A2(n_1324),
.B(n_1387),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1342),
.A2(n_1341),
.B(n_1319),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1308),
.A2(n_1409),
.B1(n_1397),
.B2(n_1416),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1322),
.A2(n_1329),
.B1(n_1358),
.B2(n_1342),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1422),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1337),
.A2(n_1360),
.B(n_1350),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1361),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_SL g1486 ( 
.A(n_1391),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1334),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1361),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1376),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1376),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1324),
.B(n_1328),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1345),
.B(n_1387),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1345),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1328),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1316),
.B(n_1425),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1397),
.B(n_1425),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1400),
.B(n_1409),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1366),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1367),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1355),
.Y(n_1500)
);

CKINVDCx9p33_ASAP7_75t_R g1501 ( 
.A(n_1419),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1400),
.B(n_1402),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1367),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1341),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1359),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1355),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1413),
.B(n_1320),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1437),
.A2(n_1419),
.B(n_1315),
.C(n_1394),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1466),
.B(n_1412),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1432),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1437),
.A2(n_1312),
.B(n_1390),
.C(n_1349),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1459),
.B(n_1347),
.C(n_1356),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1466),
.B(n_1347),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1481),
.A2(n_1329),
.B1(n_1354),
.B2(n_1343),
.C(n_1411),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1481),
.A2(n_1317),
.B1(n_1339),
.B2(n_1356),
.C(n_1338),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1448),
.A2(n_1338),
.B(n_1413),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1449),
.A2(n_1389),
.B1(n_1420),
.B2(n_1404),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1462),
.A2(n_1389),
.B1(n_1420),
.B2(n_1404),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1469),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1506),
.B(n_1325),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_SL g1524 ( 
.A1(n_1484),
.A2(n_1391),
.B(n_1423),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1462),
.A2(n_1474),
.B1(n_1477),
.B2(n_1493),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1474),
.A2(n_1325),
.B(n_1327),
.C(n_1423),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1389),
.C(n_1420),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1506),
.B(n_1327),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1457),
.B(n_1355),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1428),
.A2(n_1353),
.B(n_1404),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1434),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1467),
.A2(n_1423),
.B(n_1321),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1467),
.A2(n_1479),
.B(n_1468),
.C(n_1496),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1457),
.B(n_1446),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_SL g1535 ( 
.A1(n_1499),
.A2(n_1503),
.B(n_1498),
.C(n_1442),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1496),
.A2(n_1504),
.B1(n_1502),
.B2(n_1497),
.Y(n_1536)
);

AO32x2_ASAP7_75t_L g1537 ( 
.A1(n_1429),
.A2(n_1450),
.A3(n_1445),
.B1(n_1444),
.B2(n_1508),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1497),
.A2(n_1504),
.B1(n_1502),
.B2(n_1495),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1492),
.A2(n_1447),
.B(n_1477),
.Y(n_1539)
);

AO32x1_ASAP7_75t_L g1540 ( 
.A1(n_1505),
.A2(n_1492),
.A3(n_1495),
.B1(n_1447),
.B2(n_1490),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1471),
.B(n_1461),
.Y(n_1541)
);

NOR2x1_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1428),
.A2(n_1463),
.B(n_1467),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1465),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1487),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1472),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_SL g1547 ( 
.A1(n_1498),
.A2(n_1507),
.B(n_1443),
.C(n_1468),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1479),
.A2(n_1491),
.B(n_1443),
.C(n_1505),
.Y(n_1548)
);

AO32x2_ASAP7_75t_L g1549 ( 
.A1(n_1429),
.A2(n_1450),
.A3(n_1444),
.B1(n_1445),
.B2(n_1500),
.Y(n_1549)
);

AND2x4_ASAP7_75t_SL g1550 ( 
.A(n_1470),
.B(n_1473),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1427),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1491),
.A2(n_1494),
.B1(n_1480),
.B2(n_1493),
.C(n_1455),
.Y(n_1552)
);

BUFx5_ASAP7_75t_L g1553 ( 
.A(n_1439),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1454),
.A2(n_1431),
.B(n_1456),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1463),
.A2(n_1494),
.B(n_1498),
.C(n_1456),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1452),
.A2(n_1455),
.B1(n_1485),
.B2(n_1488),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1438),
.B(n_1452),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1485),
.A2(n_1489),
.B1(n_1426),
.B2(n_1435),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_L g1561 ( 
.A1(n_1484),
.A2(n_1476),
.B(n_1475),
.C(n_1426),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1480),
.A2(n_1460),
.B1(n_1458),
.B2(n_1464),
.C(n_1483),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1538),
.A2(n_1536),
.B1(n_1552),
.B2(n_1514),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1559),
.B(n_1438),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1554),
.B(n_1433),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1559),
.B(n_1480),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1544),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1519),
.A2(n_1435),
.B1(n_1473),
.B2(n_1501),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1554),
.B(n_1440),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1480),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1551),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1441),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1553),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1524),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1555),
.B(n_1456),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1537),
.B(n_1428),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1534),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1533),
.A2(n_1431),
.B(n_1454),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1544),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1428),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1433),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1534),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1454),
.Y(n_1583)
);

BUFx8_ASAP7_75t_SL g1584 ( 
.A(n_1545),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1557),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1550),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1436),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1430),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1549),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1531),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1516),
.A2(n_1464),
.B1(n_1460),
.B2(n_1458),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1571),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1565),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1591),
.B(n_1522),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1516),
.C(n_1513),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1577),
.B(n_1582),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1562),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1563),
.A2(n_1570),
.B1(n_1527),
.B2(n_1517),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1581),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1517),
.B1(n_1520),
.B2(n_1518),
.C(n_1532),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1583),
.B(n_1532),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1582),
.B(n_1566),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1608)
);

INVx5_ASAP7_75t_L g1609 ( 
.A(n_1575),
.Y(n_1609)
);

OAI31xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1568),
.A2(n_1561),
.A3(n_1525),
.B(n_1518),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1593),
.B(n_1548),
.C(n_1547),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1430),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1593),
.A2(n_1525),
.B1(n_1558),
.B2(n_1560),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1558),
.Y(n_1616)
);

AOI322xp5_ASAP7_75t_L g1617 ( 
.A1(n_1568),
.A2(n_1510),
.A3(n_1556),
.B1(n_1542),
.B2(n_1526),
.C1(n_1540),
.C2(n_1511),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1581),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1587),
.B(n_1553),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1572),
.B(n_1560),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1589),
.A2(n_1515),
.B1(n_1521),
.B2(n_1528),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1569),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1523),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_SL g1627 ( 
.A(n_1609),
.B(n_1576),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1611),
.B(n_1618),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1614),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1609),
.B(n_1573),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1619),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1619),
.B(n_1576),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1609),
.B(n_1573),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1595),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1623),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1580),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1569),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1595),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1595),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1608),
.B(n_1580),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1596),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1569),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1600),
.B(n_1572),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1609),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1592),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1597),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.B(n_1578),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1573),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1609),
.B(n_1594),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1620),
.B(n_1585),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1598),
.B(n_1589),
.C(n_1535),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1609),
.B(n_1594),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1597),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1612),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1636),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1636),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1650),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1649),
.B(n_1600),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1648),
.B(n_1609),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1629),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1648),
.B(n_1605),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1605),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1653),
.B(n_1605),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1625),
.B(n_1601),
.Y(n_1671)
);

NOR2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1598),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1625),
.B(n_1601),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1649),
.B(n_1651),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1628),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1597),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1643),
.B(n_1592),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1642),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1652),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1590),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1657),
.B(n_1584),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1628),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1599),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1652),
.B(n_1590),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1641),
.B(n_1613),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1606),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1606),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1660),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1629),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1644),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1644),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1641),
.B(n_1613),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1633),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1679),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1674),
.B(n_1621),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1617),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1685),
.B(n_1673),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1664),
.B(n_1641),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1664),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1691),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1682),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1617),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1680),
.B(n_1684),
.Y(n_1715)
);

AOI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1675),
.A2(n_1610),
.B(n_1611),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1694),
.B(n_1627),
.Y(n_1717)
);

O2A1O1Ixp5_ASAP7_75t_R g1718 ( 
.A1(n_1690),
.A2(n_1529),
.B(n_1564),
.C(n_1610),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1674),
.B(n_1621),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1567),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1695),
.B(n_1567),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1688),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1486),
.Y(n_1723)
);

INVxp33_ASAP7_75t_L g1724 ( 
.A(n_1699),
.Y(n_1724)
);

OAI31xp33_ASAP7_75t_L g1725 ( 
.A1(n_1665),
.A2(n_1603),
.A3(n_1615),
.B(n_1630),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1683),
.B(n_1579),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1668),
.B(n_1579),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1698),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1698),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1668),
.B(n_1624),
.Y(n_1731)
);

AOI211x1_ASAP7_75t_SL g1732 ( 
.A1(n_1667),
.A2(n_1633),
.B(n_1521),
.C(n_1623),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1689),
.B(n_1678),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1669),
.B(n_1624),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1669),
.B(n_1670),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1679),
.B(n_1618),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1701),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1678),
.B(n_1621),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1701),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1714),
.A2(n_1615),
.B(n_1665),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1663),
.C(n_1603),
.Y(n_1741)
);

AOI222xp33_ASAP7_75t_L g1742 ( 
.A1(n_1707),
.A2(n_1670),
.B1(n_1622),
.B2(n_1637),
.C1(n_1639),
.C2(n_1632),
.Y(n_1742)
);

AOI222xp33_ASAP7_75t_L g1743 ( 
.A1(n_1718),
.A2(n_1622),
.B1(n_1639),
.B2(n_1637),
.C1(n_1631),
.C2(n_1632),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1712),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1722),
.A2(n_1618),
.B1(n_1663),
.B2(n_1574),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1713),
.B(n_1679),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1728),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1708),
.A2(n_1725),
.B1(n_1723),
.B2(n_1710),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1730),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1737),
.Y(n_1751)
);

NAND4xp25_ASAP7_75t_SL g1752 ( 
.A(n_1736),
.B(n_1735),
.C(n_1711),
.D(n_1717),
.Y(n_1752)
);

AOI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1708),
.A2(n_1639),
.B1(n_1637),
.B2(n_1631),
.C1(n_1632),
.C2(n_1626),
.Y(n_1753)
);

OAI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1724),
.A2(n_1618),
.B1(n_1574),
.B2(n_1586),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1723),
.B(n_1630),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1732),
.A2(n_1530),
.B(n_1646),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1711),
.A2(n_1635),
.B1(n_1654),
.B2(n_1630),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1704),
.B(n_1656),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1739),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1724),
.A2(n_1635),
.B1(n_1630),
.B2(n_1654),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1704),
.A2(n_1541),
.B1(n_1512),
.B2(n_1584),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1715),
.A2(n_1635),
.B(n_1654),
.C(n_1630),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1733),
.A2(n_1726),
.B1(n_1720),
.B2(n_1721),
.C(n_1727),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1731),
.B(n_1692),
.Y(n_1764)
);

AOI21xp33_ASAP7_75t_L g1765 ( 
.A1(n_1709),
.A2(n_1702),
.B(n_1692),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1748),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1750),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1751),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1744),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1749),
.A2(n_1709),
.B1(n_1729),
.B2(n_1705),
.C(n_1719),
.Y(n_1770)
);

OAI31xp33_ASAP7_75t_L g1771 ( 
.A1(n_1741),
.A2(n_1717),
.A3(n_1729),
.B(n_1738),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1759),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1747),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1749),
.A2(n_1740),
.B1(n_1752),
.B2(n_1746),
.C(n_1765),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1764),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1758),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1763),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1761),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1755),
.Y(n_1779)
);

AOI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1754),
.A2(n_1734),
.B(n_1706),
.C(n_1646),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1742),
.B(n_1627),
.Y(n_1781)
);

OAI311xp33_ASAP7_75t_L g1782 ( 
.A1(n_1743),
.A2(n_1702),
.A3(n_1647),
.B1(n_1661),
.C1(n_1696),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1627),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1756),
.B(n_1706),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1745),
.B(n_1626),
.Y(n_1785)
);

AOI32xp33_ASAP7_75t_L g1786 ( 
.A1(n_1774),
.A2(n_1745),
.A3(n_1754),
.B1(n_1760),
.B2(n_1646),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1778),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1769),
.B(n_1757),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1773),
.B(n_1762),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1771),
.A2(n_1654),
.B(n_1630),
.C(n_1635),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1777),
.A2(n_1646),
.B1(n_1574),
.B2(n_1635),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1776),
.Y(n_1792)
);

OAI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1779),
.A2(n_1666),
.B(n_1661),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1770),
.A2(n_1776),
.B1(n_1781),
.B2(n_1780),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1775),
.B(n_1626),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1782),
.A2(n_1784),
.B(n_1781),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1766),
.Y(n_1797)
);

XNOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1767),
.B(n_1574),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1787),
.B(n_1784),
.C(n_1772),
.D(n_1766),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1792),
.Y(n_1800)
);

NAND4xp25_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1768),
.C(n_1785),
.D(n_1783),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1788),
.B(n_1789),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1797),
.Y(n_1803)
);

AOI322xp5_ASAP7_75t_L g1804 ( 
.A1(n_1793),
.A2(n_1783),
.A3(n_1768),
.B1(n_1640),
.B2(n_1645),
.C1(n_1631),
.C2(n_1634),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1798),
.B(n_1640),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1794),
.B(n_1647),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1796),
.B(n_1662),
.C(n_1666),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_L g1808 ( 
.A(n_1786),
.B(n_1703),
.C(n_1687),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1795),
.Y(n_1809)
);

OAI222xp33_ASAP7_75t_L g1810 ( 
.A1(n_1806),
.A2(n_1791),
.B1(n_1790),
.B2(n_1646),
.C1(n_1703),
.C2(n_1700),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1799),
.B(n_1802),
.Y(n_1811)
);

OAI211xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1809),
.A2(n_1681),
.B(n_1662),
.C(n_1676),
.Y(n_1812)
);

AOI211x1_ASAP7_75t_L g1813 ( 
.A1(n_1801),
.A2(n_1677),
.B(n_1676),
.C(n_1687),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1808),
.A2(n_1646),
.B(n_1654),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1811),
.B(n_1799),
.C(n_1800),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1812),
.A2(n_1805),
.B1(n_1807),
.B2(n_1803),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1813),
.B(n_1804),
.Y(n_1817)
);

AOI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1810),
.A2(n_1814),
.B1(n_1681),
.B2(n_1677),
.C(n_1696),
.Y(n_1818)
);

AOI21xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1811),
.A2(n_1693),
.B(n_1654),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1813),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.B(n_1693),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1820),
.B(n_1686),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1817),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1640),
.Y(n_1824)
);

NAND4xp75_ASAP7_75t_L g1825 ( 
.A(n_1818),
.B(n_1700),
.C(n_1697),
.D(n_1686),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1823),
.A2(n_1819),
.B(n_1697),
.C(n_1633),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1824),
.B(n_1633),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1822),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1828),
.Y(n_1829)
);

OAI22x1_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1821),
.B1(n_1827),
.B2(n_1826),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1825),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1830),
.A2(n_1635),
.B1(n_1658),
.B2(n_1655),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_R g1833 ( 
.A(n_1831),
.B(n_1832),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1831),
.A2(n_1638),
.B(n_1658),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1833),
.A2(n_1638),
.B(n_1655),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1638),
.B(n_1655),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1837),
.A2(n_1836),
.B(n_1658),
.Y(n_1838)
);

XNOR2xp5_ASAP7_75t_L g1839 ( 
.A(n_1838),
.B(n_1509),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1638),
.B1(n_1655),
.B2(n_1658),
.C(n_1604),
.Y(n_1840)
);

AOI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1508),
.B(n_1500),
.C(n_1478),
.Y(n_1841)
);


endmodule