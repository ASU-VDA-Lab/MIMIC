module real_jpeg_16678_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_463),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_0),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_1),
.B(n_89),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_1),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_2),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_3),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_3),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_4),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_4),
.B(n_34),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_4),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_4),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_54),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_5),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_5),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_5),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_5),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_5),
.B(n_431),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_6),
.Y(n_464)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_7),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_8),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_8),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_9),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_9),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_9),
.B(n_173),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_9),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_9),
.B(n_408),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_9),
.B(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_10),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_12),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_12),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_12),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_12),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_12),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_12),
.B(n_188),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_14),
.B(n_102),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_14),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_14),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_14),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_14),
.B(n_383),
.Y(n_382)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_15),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_54),
.Y(n_53)
);

AND2x4_ASAP7_75t_SL g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_16),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_16),
.B(n_172),
.Y(n_171)
);

NAND2x2_ASAP7_75t_SL g197 ( 
.A(n_16),
.B(n_198),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_201),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_200),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_155),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_23),
.B(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_130),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_72),
.B2(n_73),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_44),
.C(n_52),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_33),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_33),
.B(n_230),
.C(n_232),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_33),
.A2(n_41),
.B1(n_230),
.B2(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_36),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_37),
.B(n_84),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_38),
.B(n_85),
.C(n_241),
.Y(n_240)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_39),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_56),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_50),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_50),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_97),
.C(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_52),
.A2(n_53),
.B1(n_97),
.B2(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_53),
.B(n_187),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_55),
.Y(n_377)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_55),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.C(n_66),
.Y(n_56)
);

INVxp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_63),
.B(n_166),
.C(n_171),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_63),
.A2(n_77),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_65),
.Y(n_361)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_92),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_90),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_78),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.C(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_79),
.A2(n_80),
.B1(n_86),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_83),
.Y(n_231)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_88),
.Y(n_233)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2x2_ASAP7_75t_SL g158 ( 
.A(n_90),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_112),
.B2(n_113),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_107),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_97),
.A2(n_137),
.B1(n_145),
.B2(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_97),
.B(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_103),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_150),
.C(n_153),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_108),
.B1(n_153),
.B2(n_154),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_111),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_111),
.Y(n_260)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_122),
.B(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_125),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_151),
.C(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_128),
.B1(n_152),
.B2(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_146),
.C(n_149),
.Y(n_130)
);

XOR2x1_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_143),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_132),
.B(n_135),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_137),
.A2(n_164),
.B1(n_222),
.B2(n_223),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_142),
.A2(n_266),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_143),
.B(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_145),
.B(n_382),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_156),
.B(n_158),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_160),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_178),
.C(n_181),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_161),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_175),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_162),
.B(n_165),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_166),
.A2(n_167),
.B1(n_171),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

XOR2x2_ASAP7_75t_L g284 ( 
.A(n_175),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_331)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.C(n_197),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_183),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_191),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_184),
.B(n_187),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_189),
.Y(n_379)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_193),
.A2(n_197),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_193),
.Y(n_291)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_195),
.Y(n_417)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_347),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_324),
.B(n_338),
.C(n_339),
.D(n_346),
.Y(n_203)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_296),
.B(n_323),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_281),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_206),
.B(n_281),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_253),
.C(n_274),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_207),
.B(n_298),
.Y(n_297)
);

XOR2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_234),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_208),
.B(n_235),
.C(n_239),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.C(n_229),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_209),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJx3_ASAP7_75t_L g280 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_213),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_217),
.B(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_220),
.A2(n_221),
.B1(n_229),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_230),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_245),
.C(n_250),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.C(n_265),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_256),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_264),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_450),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_284),
.C(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_287),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_294),
.C(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_299),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.C(n_307),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_300),
.A2(n_301),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_307),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.C(n_312),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_308),
.B(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_311),
.B(n_312),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.C(n_322),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2x2_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_401),
.Y(n_400)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_322),
.Y(n_402)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_325),
.B(n_340),
.Y(n_349)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_336),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_336),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_342),
.C(n_343),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_344),
.Y(n_346)
);

NAND4xp25_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.C(n_350),
.D(n_351),
.Y(n_347)
);

OAI21x1_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_456),
.B(n_462),
.Y(n_351)
);

AOI21x1_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_444),
.B(n_455),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_403),
.B(n_443),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_387),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_355),
.B(n_387),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_373),
.C(n_380),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_440),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_369),
.C(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_369),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_373),
.A2(n_380),
.B1(n_381),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_378),
.Y(n_413)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_397),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_398),
.C(n_400),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_392),
.C(n_395),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_392),
.B1(n_395),
.B2(n_396),
.Y(n_390)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_391),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_392),
.Y(n_396)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_437),
.B(n_442),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_424),
.B(n_436),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_412),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_406),
.B(n_412),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_411),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_411),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_416),
.C(n_418),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_418),
.B2(n_419),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_429),
.B(n_435),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_428),
.Y(n_435)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_439),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_454),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_SL g455 ( 
.A(n_445),
.B(n_454),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_452),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_457)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_458),
.Y(n_462)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);


endmodule