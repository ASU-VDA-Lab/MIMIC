module fake_jpeg_3804_n_79 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_20),
.B1(n_0),
.B2(n_8),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_51),
.B(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_32),
.B1(n_45),
.B2(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_57),
.B(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_62),
.B1(n_48),
.B2(n_30),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_46),
.C(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_56),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_54),
.B1(n_30),
.B2(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_40),
.B1(n_36),
.B2(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_47),
.C(n_25),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_35),
.B(n_28),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_59),
.B(n_54),
.C(n_58),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_63),
.A3(n_26),
.B1(n_34),
.B2(n_41),
.C1(n_23),
.C2(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_49),
.B1(n_26),
.B2(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_76),
.B1(n_34),
.B2(n_41),
.C(n_23),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_55),
.Y(n_79)
);


endmodule