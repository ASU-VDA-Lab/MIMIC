module fake_jpeg_12007_n_182 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_5),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_0),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_69),
.B(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_64),
.B1(n_62),
.B2(n_68),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_78),
.B1(n_64),
.B2(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_76),
.B1(n_78),
.B2(n_73),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_R g100 ( 
.A(n_83),
.B(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_75),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_115),
.B1(n_118),
.B2(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_125),
.B1(n_11),
.B2(n_51),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_7),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_67),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_113),
.B(n_10),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_77),
.C(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_60),
.B1(n_66),
.B2(n_59),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_120),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_32),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_60),
.B1(n_65),
.B2(n_72),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_37),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_60),
.B1(n_67),
.B2(n_57),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_139),
.B(n_145),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_9),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_142),
.B(n_146),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_42),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_132),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_16),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_152),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_29),
.B(n_30),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_157),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_35),
.B(n_38),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_39),
.C(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_143),
.B(n_49),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_46),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_147),
.B(n_155),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_173),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_169),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_177),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.A3(n_174),
.B1(n_168),
.B2(n_170),
.C1(n_161),
.C2(n_163),
.Y(n_179)
);

AOI21x1_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_159),
.B(n_157),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_180),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_167),
.Y(n_182)
);


endmodule