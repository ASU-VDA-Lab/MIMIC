module real_aes_10105_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_315;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1162;
wire n_762;
wire n_325;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_304;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_0), .A2(n_204), .B1(n_325), .B2(n_327), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_0), .A2(n_204), .B1(n_342), .B2(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_1), .A2(n_15), .B1(n_762), .B2(n_771), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_1), .A2(n_218), .B1(n_397), .B2(n_811), .Y(n_991) );
INVx1_ASAP7_75t_L g1022 ( .A(n_2), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_3), .A2(n_100), .B1(n_451), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_3), .A2(n_100), .B1(n_624), .B2(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_SL g827 ( .A(n_4), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_4), .A2(n_17), .B1(n_451), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g1242 ( .A(n_5), .Y(n_1242) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_6), .Y(n_246) );
INVx1_ASAP7_75t_L g350 ( .A(n_6), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_7), .A2(n_84), .B1(n_534), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_7), .A2(n_84), .B1(n_571), .B2(n_573), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_8), .A2(n_192), .B1(n_329), .B2(n_334), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_8), .A2(n_192), .B1(n_361), .B2(n_799), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_9), .A2(n_158), .B1(n_329), .B2(n_334), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_9), .A2(n_158), .B1(n_799), .B2(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_10), .A2(n_226), .B1(n_361), .B2(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_10), .A2(n_226), .B1(n_807), .B2(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g1115 ( .A(n_11), .Y(n_1115) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_11), .A2(n_1226), .B1(n_1284), .B2(n_1286), .C1(n_1290), .C2(n_1294), .Y(n_1225) );
AO22x2_ASAP7_75t_L g1229 ( .A1(n_11), .A2(n_1115), .B1(n_1230), .B2(n_1283), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_12), .A2(n_116), .B1(n_571), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_12), .A2(n_116), .B1(n_534), .B2(n_544), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_13), .Y(n_938) );
INVx1_ASAP7_75t_L g821 ( .A(n_14), .Y(n_821) );
INVx1_ASAP7_75t_L g979 ( .A(n_15), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g1259 ( .A1(n_16), .A2(n_225), .B1(n_724), .B2(n_1260), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_16), .A2(n_225), .B1(n_678), .B2(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g826 ( .A(n_17), .Y(n_826) );
INVx1_ASAP7_75t_L g859 ( .A(n_18), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_18), .A2(n_113), .B1(n_338), .B2(n_457), .Y(n_883) );
XNOR2xp5_ASAP7_75t_L g947 ( .A(n_19), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1063 ( .A(n_19), .Y(n_1063) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_20), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_20), .A2(n_181), .B1(n_632), .B2(n_634), .Y(n_631) );
INVxp33_ASAP7_75t_L g700 ( .A(n_21), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_21), .A2(n_201), .B1(n_737), .B2(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g267 ( .A(n_22), .Y(n_267) );
INVx1_ASAP7_75t_L g816 ( .A(n_23), .Y(n_816) );
AO221x2_ASAP7_75t_L g1044 ( .A1(n_24), .A2(n_48), .B1(n_1020), .B2(n_1035), .C(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1046 ( .A(n_25), .Y(n_1046) );
INVx1_ASAP7_75t_L g519 ( .A(n_26), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_26), .A2(n_103), .B1(n_539), .B2(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g429 ( .A(n_27), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_27), .A2(n_194), .B1(n_456), .B2(n_457), .Y(n_455) );
BUFx2_ASAP7_75t_L g313 ( .A(n_28), .Y(n_313) );
BUFx2_ASAP7_75t_L g353 ( .A(n_28), .Y(n_353) );
INVx1_ASAP7_75t_L g551 ( .A(n_28), .Y(n_551) );
INVx1_ASAP7_75t_L g512 ( .A(n_29), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_29), .A2(n_90), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g1113 ( .A(n_30), .Y(n_1113) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_31), .A2(n_98), .B1(n_361), .B2(n_362), .Y(n_360) );
INVxp67_ASAP7_75t_L g392 ( .A(n_31), .Y(n_392) );
INVx1_ASAP7_75t_L g528 ( .A(n_32), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_32), .A2(n_40), .B1(n_534), .B2(n_536), .Y(n_533) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_33), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_33), .A2(n_108), .B1(n_415), .B2(n_599), .Y(n_598) );
INVxp33_ASAP7_75t_L g658 ( .A(n_34), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_34), .A2(n_138), .B1(n_556), .B2(n_670), .Y(n_669) );
AO22x2_ASAP7_75t_L g498 ( .A1(n_35), .A2(n_499), .B1(n_500), .B2(n_575), .Y(n_498) );
INVx1_ASAP7_75t_L g575 ( .A(n_35), .Y(n_575) );
INVx1_ASAP7_75t_L g989 ( .A(n_36), .Y(n_989) );
INVx1_ASAP7_75t_L g709 ( .A(n_37), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_37), .A2(n_126), .B1(n_723), .B2(n_733), .Y(n_732) );
CKINVDCx16_ASAP7_75t_R g1060 ( .A(n_38), .Y(n_1060) );
INVx1_ASAP7_75t_L g1109 ( .A(n_39), .Y(n_1109) );
INVx1_ASAP7_75t_L g521 ( .A(n_40), .Y(n_521) );
INVx1_ASAP7_75t_L g862 ( .A(n_41), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_41), .A2(n_215), .B1(n_334), .B2(n_718), .Y(n_882) );
INVx1_ASAP7_75t_L g820 ( .A(n_42), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_42), .A2(n_174), .B1(n_457), .B2(n_667), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_43), .A2(n_223), .B1(n_675), .B2(n_799), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_43), .A2(n_159), .B1(n_397), .B2(n_811), .Y(n_941) );
INVx1_ASAP7_75t_L g1236 ( .A(n_44), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_45), .A2(n_127), .B1(n_411), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_45), .A2(n_127), .B1(n_358), .B2(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g511 ( .A(n_46), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_46), .A2(n_62), .B1(n_559), .B2(n_562), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_47), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_49), .A2(n_206), .B1(n_357), .B2(n_358), .Y(n_356) );
INVxp33_ASAP7_75t_L g395 ( .A(n_49), .Y(n_395) );
INVxp33_ASAP7_75t_L g650 ( .A(n_50), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_50), .A2(n_82), .B1(n_357), .B2(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_51), .A2(n_73), .B1(n_759), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g782 ( .A(n_51), .Y(n_782) );
INVx1_ASAP7_75t_L g914 ( .A(n_52), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_52), .A2(n_159), .B1(n_759), .B2(n_762), .Y(n_933) );
INVx1_ASAP7_75t_L g1074 ( .A(n_53), .Y(n_1074) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_54), .A2(n_216), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_54), .A2(n_216), .B1(n_716), .B2(n_730), .C(n_781), .Y(n_780) );
CKINVDCx16_ASAP7_75t_R g1077 ( .A(n_55), .Y(n_1077) );
INVx1_ASAP7_75t_L g988 ( .A(n_56), .Y(n_988) );
INVx1_ASAP7_75t_L g960 ( .A(n_57), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_58), .A2(n_211), .B1(n_716), .B2(n_719), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_58), .A2(n_211), .B1(n_740), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g647 ( .A(n_59), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_60), .A2(n_230), .B1(n_329), .B2(n_334), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_60), .A2(n_230), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g1026 ( .A(n_61), .Y(n_1026) );
OAI222xp33_ASAP7_75t_L g503 ( .A1(n_62), .A2(n_141), .B1(n_220), .B2(n_504), .C1(n_507), .C2(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g698 ( .A(n_63), .Y(n_698) );
INVx1_ASAP7_75t_L g876 ( .A(n_64), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_64), .A2(n_74), .B1(n_323), .B2(n_361), .Y(n_889) );
INVx1_ASAP7_75t_L g910 ( .A(n_65), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_65), .A2(n_150), .B1(n_770), .B2(n_771), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_66), .A2(n_133), .B1(n_338), .B2(n_457), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_66), .A2(n_133), .B1(n_325), .B2(n_327), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_67), .A2(n_93), .B1(n_509), .B2(n_867), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_67), .A2(n_93), .B1(n_485), .B2(n_599), .Y(n_871) );
INVx1_ASAP7_75t_L g834 ( .A(n_68), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_68), .A2(n_87), .B1(n_323), .B2(n_361), .Y(n_853) );
INVx1_ASAP7_75t_L g965 ( .A(n_69), .Y(n_965) );
OAI211xp5_ASAP7_75t_SL g992 ( .A1(n_69), .A2(n_424), .B(n_943), .C(n_993), .Y(n_992) );
AO22x2_ASAP7_75t_L g639 ( .A1(n_70), .A2(n_640), .B1(n_681), .B2(n_682), .Y(n_639) );
INVx1_ASAP7_75t_L g681 ( .A(n_70), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g1079 ( .A(n_71), .Y(n_1079) );
AO22x2_ASAP7_75t_L g402 ( .A1(n_72), .A2(n_403), .B1(n_473), .B2(n_474), .Y(n_402) );
INVxp67_ASAP7_75t_L g473 ( .A(n_72), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_72), .A2(n_123), .B1(n_1029), .B2(n_1032), .Y(n_1041) );
INVx1_ASAP7_75t_L g805 ( .A(n_73), .Y(n_805) );
INVx1_ASAP7_75t_L g874 ( .A(n_74), .Y(n_874) );
INVx1_ASAP7_75t_L g291 ( .A(n_75), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_75), .A2(n_81), .B1(n_378), .B2(n_381), .Y(n_377) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_76), .Y(n_1237) );
AOI22xp33_ASAP7_75t_SL g1262 ( .A1(n_76), .A2(n_180), .B1(n_553), .B2(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g311 ( .A(n_77), .Y(n_311) );
INVxp33_ASAP7_75t_SL g1247 ( .A(n_78), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_78), .A2(n_173), .B1(n_546), .B2(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1239 ( .A(n_79), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_79), .A2(n_165), .B1(n_1260), .B2(n_1266), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_80), .A2(n_111), .B1(n_553), .B2(n_1257), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_80), .A2(n_111), .B1(n_1272), .B2(n_1274), .Y(n_1271) );
INVx1_ASAP7_75t_L g298 ( .A(n_81), .Y(n_298) );
INVx1_ASAP7_75t_L g646 ( .A(n_82), .Y(n_646) );
INVx1_ASAP7_75t_L g930 ( .A(n_83), .Y(n_930) );
OAI211xp5_ASAP7_75t_SL g942 ( .A1(n_83), .A2(n_424), .B(n_943), .C(n_945), .Y(n_942) );
INVx1_ASAP7_75t_L g776 ( .A(n_85), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_86), .A2(n_169), .B1(n_504), .B2(n_509), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_86), .A2(n_169), .B1(n_378), .B2(n_599), .Y(n_831) );
INVxp67_ASAP7_75t_L g836 ( .A(n_87), .Y(n_836) );
INVx1_ASAP7_75t_L g954 ( .A(n_88), .Y(n_954) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_89), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_89), .A2(n_219), .B1(n_616), .B2(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g515 ( .A(n_90), .Y(n_515) );
INVx1_ASAP7_75t_L g982 ( .A(n_91), .Y(n_982) );
INVx1_ASAP7_75t_L g406 ( .A(n_92), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_92), .A2(n_200), .B1(n_323), .B2(n_361), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_94), .A2(n_119), .B1(n_541), .B2(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_94), .A2(n_119), .B1(n_565), .B2(n_567), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_95), .A2(n_185), .B1(n_367), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_95), .A2(n_185), .B1(n_460), .B2(n_461), .Y(n_459) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_96), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_96), .A2(n_168), .B1(n_463), .B2(n_799), .Y(n_924) );
INVx1_ASAP7_75t_L g1062 ( .A(n_97), .Y(n_1062) );
INVxp33_ASAP7_75t_L g388 ( .A(n_98), .Y(n_388) );
AO221x2_ASAP7_75t_L g1014 ( .A1(n_99), .A2(n_157), .B1(n_1015), .B2(n_1020), .C(n_1021), .Y(n_1014) );
INVx1_ASAP7_75t_L g964 ( .A(n_101), .Y(n_964) );
OAI22xp33_ASAP7_75t_SL g994 ( .A1(n_101), .A2(n_131), .B1(n_247), .B2(n_807), .Y(n_994) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_102), .A2(n_260), .B1(n_399), .B2(n_400), .Y(n_259) );
INVx1_ASAP7_75t_L g399 ( .A(n_102), .Y(n_399) );
INVx1_ASAP7_75t_L g518 ( .A(n_103), .Y(n_518) );
INVx1_ASAP7_75t_L g238 ( .A(n_104), .Y(n_238) );
INVx1_ASAP7_75t_L g873 ( .A(n_105), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_105), .A2(n_186), .B1(n_325), .B2(n_461), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_106), .A2(n_187), .B1(n_553), .B2(n_774), .C(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_106), .A2(n_187), .B1(n_323), .B2(n_361), .Y(n_794) );
INVx1_ASAP7_75t_L g768 ( .A(n_107), .Y(n_768) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_108), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_109), .A2(n_152), .B1(n_1020), .B2(n_1035), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_110), .Y(n_422) );
INVx1_ASAP7_75t_L g302 ( .A(n_112), .Y(n_302) );
INVx1_ASAP7_75t_L g865 ( .A(n_113), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_114), .A2(n_142), .B1(n_565), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_114), .A2(n_142), .B1(n_539), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_115), .A2(n_121), .B1(n_322), .B2(n_323), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_115), .A2(n_121), .B1(n_329), .B2(n_334), .Y(n_365) );
INVx1_ASAP7_75t_L g689 ( .A(n_117), .Y(n_689) );
CKINVDCx14_ASAP7_75t_R g755 ( .A(n_118), .Y(n_755) );
XOR2xp5_ASAP7_75t_L g891 ( .A(n_120), .B(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g767 ( .A(n_122), .Y(n_767) );
INVxp33_ASAP7_75t_SL g273 ( .A(n_124), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_124), .A2(n_135), .B1(n_338), .B2(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g651 ( .A(n_125), .Y(n_651) );
INVxp33_ASAP7_75t_L g704 ( .A(n_126), .Y(n_704) );
INVxp33_ASAP7_75t_L g644 ( .A(n_128), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_128), .A2(n_136), .B1(n_675), .B2(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g957 ( .A(n_129), .Y(n_957) );
INVx1_ASAP7_75t_L g648 ( .A(n_130), .Y(n_648) );
INVx1_ASAP7_75t_L g967 ( .A(n_131), .Y(n_967) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_132), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_132), .A2(n_183), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_134), .A2(n_144), .B1(n_1029), .B2(n_1032), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_135), .Y(n_287) );
INVxp33_ASAP7_75t_L g643 ( .A(n_136), .Y(n_643) );
INVxp33_ASAP7_75t_SL g304 ( .A(n_137), .Y(n_304) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_137), .A2(n_155), .B1(n_329), .B2(n_334), .Y(n_328) );
INVxp33_ASAP7_75t_L g660 ( .A(n_138), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_139), .A2(n_198), .B1(n_411), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_139), .A2(n_198), .B1(n_327), .B2(n_468), .Y(n_673) );
INVx1_ASAP7_75t_L g902 ( .A(n_140), .Y(n_902) );
INVx1_ASAP7_75t_L g525 ( .A(n_141), .Y(n_525) );
INVx1_ASAP7_75t_L g978 ( .A(n_143), .Y(n_978) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_143), .A2(n_154), .B1(n_759), .B2(n_770), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_145), .A2(n_189), .B1(n_1015), .B2(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g693 ( .A(n_146), .Y(n_693) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_147), .B(n_238), .Y(n_1007) );
AND3x2_ASAP7_75t_L g1019 ( .A(n_147), .B(n_238), .C(n_1006), .Y(n_1019) );
INVxp33_ASAP7_75t_SL g591 ( .A(n_148), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_148), .A2(n_210), .B1(n_373), .B2(n_571), .Y(n_614) );
INVxp33_ASAP7_75t_L g661 ( .A(n_149), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_149), .A2(n_153), .B1(n_367), .B2(n_411), .Y(n_671) );
INVx1_ASAP7_75t_L g912 ( .A(n_150), .Y(n_912) );
INVx2_ASAP7_75t_L g251 ( .A(n_151), .Y(n_251) );
INVx1_ASAP7_75t_L g656 ( .A(n_153), .Y(n_656) );
INVx1_ASAP7_75t_L g981 ( .A(n_154), .Y(n_981) );
INVxp33_ASAP7_75t_SL g282 ( .A(n_155), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_156), .A2(n_162), .B1(n_1020), .B2(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1006 ( .A(n_160), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_161), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_161), .A2(n_196), .B1(n_323), .B2(n_749), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g1058 ( .A(n_163), .Y(n_1058) );
INVx1_ASAP7_75t_L g1111 ( .A(n_164), .Y(n_1111) );
INVxp33_ASAP7_75t_SL g1233 ( .A(n_165), .Y(n_1233) );
INVx1_ASAP7_75t_L g438 ( .A(n_166), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_166), .A2(n_207), .B1(n_451), .B2(n_452), .Y(n_450) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_167), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_167), .A2(n_203), .B1(n_288), .B2(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_168), .Y(n_904) );
INVx1_ASAP7_75t_L g899 ( .A(n_170), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_171), .Y(n_860) );
INVx1_ASAP7_75t_L g796 ( .A(n_172), .Y(n_796) );
INVxp33_ASAP7_75t_SL g1248 ( .A(n_173), .Y(n_1248) );
INVx1_ASAP7_75t_L g823 ( .A(n_174), .Y(n_823) );
INVx1_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
INVx2_ASAP7_75t_L g349 ( .A(n_175), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g763 ( .A1(n_176), .A2(n_262), .B(n_764), .C(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g785 ( .A(n_176), .Y(n_785) );
INVx1_ASAP7_75t_L g830 ( .A(n_177), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_177), .A2(n_222), .B1(n_460), .B2(n_461), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_178), .A2(n_205), .B1(n_447), .B2(n_667), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_178), .A2(n_205), .B1(n_470), .B2(n_848), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g855 ( .A(n_179), .B(n_856), .Y(n_855) );
INVxp33_ASAP7_75t_SL g1234 ( .A(n_180), .Y(n_1234) );
INVxp33_ASAP7_75t_SL g602 ( .A(n_181), .Y(n_602) );
AO22x2_ASAP7_75t_L g580 ( .A1(n_182), .A2(n_581), .B1(n_636), .B2(n_637), .Y(n_580) );
CKINVDCx14_ASAP7_75t_R g636 ( .A(n_182), .Y(n_636) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_183), .Y(n_707) );
INVx1_ASAP7_75t_L g410 ( .A(n_184), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_184), .A2(n_229), .B1(n_468), .B2(n_470), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_184), .A2(n_424), .B(n_478), .C(n_483), .Y(n_477) );
INVx1_ASAP7_75t_L g870 ( .A(n_186), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_188), .A2(n_209), .B1(n_1029), .B2(n_1032), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_190), .Y(n_696) );
INVx1_ASAP7_75t_L g778 ( .A(n_191), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_193), .Y(n_514) );
INVx1_ASAP7_75t_L g434 ( .A(n_194), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g490 ( .A1(n_194), .A2(n_262), .B(n_491), .C(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g927 ( .A(n_195), .Y(n_927) );
OAI22xp33_ASAP7_75t_SL g946 ( .A1(n_195), .A2(n_223), .B1(n_247), .B2(n_807), .Y(n_946) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_196), .Y(n_701) );
INVx1_ASAP7_75t_L g588 ( .A(n_197), .Y(n_588) );
INVx1_ASAP7_75t_L g1075 ( .A(n_199), .Y(n_1075) );
INVx1_ASAP7_75t_L g407 ( .A(n_200), .Y(n_407) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_201), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_202), .B(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1018 ( .A(n_202), .Y(n_1018) );
INVxp33_ASAP7_75t_SL g595 ( .A(n_203), .Y(n_595) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_206), .Y(n_372) );
INVx1_ASAP7_75t_L g431 ( .A(n_207), .Y(n_431) );
INVx1_ASAP7_75t_L g952 ( .A(n_208), .Y(n_952) );
INVx1_ASAP7_75t_L g584 ( .A(n_210), .Y(n_584) );
INVx1_ASAP7_75t_L g1243 ( .A(n_212), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_213), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_214), .Y(n_937) );
INVx1_ASAP7_75t_L g863 ( .A(n_215), .Y(n_863) );
INVx2_ASAP7_75t_L g250 ( .A(n_217), .Y(n_250) );
INVx1_ASAP7_75t_L g969 ( .A(n_218), .Y(n_969) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_219), .Y(n_592) );
INVx1_ASAP7_75t_L g526 ( .A(n_220), .Y(n_526) );
INVxp33_ASAP7_75t_SL g1253 ( .A(n_221), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_221), .A2(n_233), .B1(n_1277), .B2(n_1279), .Y(n_1276) );
INVxp33_ASAP7_75t_L g833 ( .A(n_222), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_224), .A2(n_1287), .B1(n_1288), .B2(n_1289), .Y(n_1286) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_224), .Y(n_1288) );
BUFx3_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
INVx1_ASAP7_75t_L g308 ( .A(n_227), .Y(n_308) );
BUFx3_ASAP7_75t_L g271 ( .A(n_228), .Y(n_271) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
INVx1_ASAP7_75t_L g421 ( .A(n_229), .Y(n_421) );
INVx1_ASAP7_75t_L g797 ( .A(n_231), .Y(n_797) );
INVx1_ASAP7_75t_L g916 ( .A(n_232), .Y(n_916) );
INVx1_ASAP7_75t_L g1250 ( .A(n_233), .Y(n_1250) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_254), .B(n_997), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_241), .Y(n_235) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_236), .B(n_242), .Y(n_1285) );
NOR2xp33_ASAP7_75t_SL g236 ( .A(n_237), .B(n_239), .Y(n_236) );
INVx1_ASAP7_75t_SL g1293 ( .A(n_237), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_237), .B(n_239), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_239), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g398 ( .A(n_244), .B(n_353), .Y(n_398) );
OR2x6_ASAP7_75t_L g426 ( .A(n_244), .B(n_353), .Y(n_426) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g369 ( .A(n_245), .B(n_253), .Y(n_369) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g896 ( .A(n_246), .B(n_387), .Y(n_896) );
INVx8_ASAP7_75t_L g394 ( .A(n_247), .Y(n_394) );
OR2x6_ASAP7_75t_L g247 ( .A(n_248), .B(n_252), .Y(n_247) );
OR2x6_ASAP7_75t_L g397 ( .A(n_248), .B(n_386), .Y(n_397) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_248), .Y(n_777) );
INVx2_ASAP7_75t_SL g784 ( .A(n_248), .Y(n_784) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_248), .Y(n_898) );
INVx2_ASAP7_75t_SL g974 ( .A(n_248), .Y(n_974) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g331 ( .A(n_250), .Y(n_331) );
AND2x4_ASAP7_75t_L g335 ( .A(n_250), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g341 ( .A(n_250), .B(n_251), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_250), .Y(n_344) );
INVx1_ASAP7_75t_L g383 ( .A(n_250), .Y(n_383) );
INVx1_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
INVx2_ASAP7_75t_L g336 ( .A(n_251), .Y(n_336) );
INVx1_ASAP7_75t_L g380 ( .A(n_251), .Y(n_380) );
INVx1_ASAP7_75t_L g482 ( .A(n_251), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_251), .B(n_331), .Y(n_810) );
AND2x4_ASAP7_75t_L g379 ( .A(n_252), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g381 ( .A(n_253), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g599 ( .A(n_253), .B(n_382), .Y(n_599) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_685), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B1(n_578), .B2(n_684), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
XNOR2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_401), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g400 ( .A(n_260), .Y(n_400) );
AOI211x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_309), .B(n_314), .C(n_370), .Y(n_260) );
NAND4xp25_ASAP7_75t_L g261 ( .A(n_262), .B(n_272), .C(n_286), .D(n_301), .Y(n_261) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_262), .B(n_583), .C(n_587), .D(n_590), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g934 ( .A(n_262), .B(n_935), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g986 ( .A(n_262), .B(n_987), .Y(n_986) );
CKINVDCx8_ASAP7_75t_R g262 ( .A(n_263), .Y(n_262) );
INVx5_ASAP7_75t_L g439 ( .A(n_263), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_263), .B(n_503), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_263), .A2(n_303), .B1(n_305), .B2(n_651), .C(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x6_ASAP7_75t_L g283 ( .A(n_265), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g760 ( .A(n_265), .Y(n_760) );
AND2x2_ASAP7_75t_L g765 ( .A(n_265), .B(n_327), .Y(n_765) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x6_ASAP7_75t_L g299 ( .A(n_266), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_311), .Y(n_320) );
INVx2_ASAP7_75t_L g355 ( .A(n_267), .Y(n_355) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_268), .Y(n_327) );
INVx2_ASAP7_75t_L g359 ( .A(n_268), .Y(n_359) );
INVx1_ASAP7_75t_L g471 ( .A(n_268), .Y(n_471) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_268), .Y(n_655) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g280 ( .A(n_270), .Y(n_280) );
AND2x4_ASAP7_75t_L g284 ( .A(n_270), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g281 ( .A(n_271), .Y(n_281) );
AND2x4_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_282), .B2(n_283), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_274), .A2(n_283), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_274), .A2(n_283), .B1(n_704), .B2(n_705), .Y(n_703) );
AOI22xp5_ASAP7_75t_SL g819 ( .A1(n_274), .A2(n_303), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_274), .A2(n_283), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
AND2x6_ASAP7_75t_L g305 ( .A(n_275), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g430 ( .A(n_275), .B(n_277), .Y(n_430) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g505 ( .A(n_276), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_278), .Y(n_469) );
INVx2_ASAP7_75t_L g535 ( .A(n_278), .Y(n_535) );
INVx2_ASAP7_75t_SL g630 ( .A(n_278), .Y(n_630) );
INVx2_ASAP7_75t_L g738 ( .A(n_278), .Y(n_738) );
INVx1_ASAP7_75t_L g848 ( .A(n_278), .Y(n_848) );
HB1xp67_ASAP7_75t_L g1278 ( .A(n_278), .Y(n_1278) );
INVx6_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g303 ( .A(n_279), .B(n_293), .Y(n_303) );
INVx2_ASAP7_75t_L g326 ( .A(n_279), .Y(n_326) );
BUFx2_ASAP7_75t_L g460 ( .A(n_279), .Y(n_460) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
INVx1_ASAP7_75t_L g297 ( .A(n_281), .Y(n_297) );
AOI22xp5_ASAP7_75t_SL g428 ( .A1(n_283), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_283), .A2(n_430), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_283), .A2(n_430), .B1(n_660), .B2(n_661), .Y(n_659) );
CKINVDCx6p67_ASAP7_75t_R g770 ( .A(n_283), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_283), .A2(n_305), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_283), .A2(n_305), .B1(n_862), .B2(n_863), .Y(n_861) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
BUFx3_ASAP7_75t_L g361 ( .A(n_284), .Y(n_361) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_284), .Y(n_463) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_284), .Y(n_540) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_284), .Y(n_546) );
INVx2_ASAP7_75t_SL g633 ( .A(n_284), .Y(n_633) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_284), .Y(n_675) );
INVx1_ASAP7_75t_L g495 ( .A(n_285), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_291), .B2(n_292), .C1(n_298), .C2(n_299), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_290), .Y(n_461) );
INVx2_ASAP7_75t_SL g537 ( .A(n_290), .Y(n_537) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_290), .Y(n_678) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_290), .Y(n_1279) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_292), .A2(n_299), .B1(n_647), .B2(n_648), .C1(n_654), .C2(n_656), .Y(n_653) );
AND2x2_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AND2x4_ASAP7_75t_L g436 ( .A(n_293), .B(n_295), .Y(n_436) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g506 ( .A(n_296), .Y(n_506) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_299), .A2(n_413), .B1(n_416), .B2(n_433), .C1(n_434), .C2(n_435), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_299), .A2(n_413), .B1(n_416), .B2(n_436), .Y(n_496) );
INVx3_ASAP7_75t_L g509 ( .A(n_299), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g583 ( .A1(n_299), .A2(n_436), .B1(n_470), .B2(n_584), .C1(n_585), .C2(n_586), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g708 ( .A1(n_299), .A2(n_435), .B1(n_696), .B2(n_698), .C1(n_709), .C2(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_299), .A2(n_436), .B1(n_767), .B2(n_768), .Y(n_766) );
AOI222xp33_ASAP7_75t_L g935 ( .A1(n_299), .A2(n_505), .B1(n_916), .B2(n_936), .C1(n_937), .C2(n_938), .Y(n_935) );
AOI222xp33_ASAP7_75t_L g987 ( .A1(n_299), .A2(n_505), .B1(n_544), .B2(n_982), .C1(n_988), .C2(n_989), .Y(n_987) );
AOI222xp33_ASAP7_75t_L g1238 ( .A1(n_299), .A2(n_435), .B1(n_1239), .B2(n_1240), .C1(n_1242), .C2(n_1243), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_304), .B2(n_305), .Y(n_301) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_302), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_303), .A2(n_305), .B1(n_422), .B2(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_303), .A2(n_305), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_303), .A2(n_305), .B1(n_588), .B2(n_589), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_303), .A2(n_305), .B1(n_693), .B2(n_707), .Y(n_706) );
INVx4_ASAP7_75t_L g762 ( .A(n_303), .Y(n_762) );
AOI22xp5_ASAP7_75t_SL g858 ( .A1(n_303), .A2(n_430), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_303), .A2(n_305), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
INVx4_ASAP7_75t_L g771 ( .A(n_305), .Y(n_771) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
INVx1_ASAP7_75t_L g625 ( .A(n_306), .Y(n_625) );
INVx1_ASAP7_75t_L g635 ( .A(n_306), .Y(n_635) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_306), .Y(n_680) );
INVx2_ASAP7_75t_L g968 ( .A(n_306), .Y(n_968) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
INVx1_ASAP7_75t_L g465 ( .A(n_307), .Y(n_465) );
INVx1_ASAP7_75t_L g743 ( .A(n_307), .Y(n_743) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_307), .Y(n_799) );
INVx1_ASAP7_75t_L g494 ( .A(n_308), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g757 ( .A1(n_309), .A2(n_758), .A3(n_763), .B(n_769), .Y(n_757) );
AOI211xp5_ASAP7_75t_L g817 ( .A1(n_309), .A2(n_818), .B(n_828), .C(n_837), .Y(n_817) );
AOI211xp5_ASAP7_75t_L g856 ( .A1(n_309), .A2(n_857), .B(n_868), .C(n_877), .Y(n_856) );
OAI31xp33_ASAP7_75t_SL g932 ( .A1(n_309), .A2(n_933), .A3(n_934), .B(n_939), .Y(n_932) );
OAI31xp33_ASAP7_75t_L g983 ( .A1(n_309), .A2(n_984), .A3(n_985), .B(n_986), .Y(n_983) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
AND2x4_ASAP7_75t_L g441 ( .A(n_310), .B(n_312), .Y(n_441) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g354 ( .A(n_311), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g318 ( .A(n_313), .Y(n_318) );
OR2x6_ASAP7_75t_L g895 ( .A(n_313), .B(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_351), .Y(n_314) );
AOI33xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_321), .A3(n_324), .B1(n_328), .B2(n_337), .B3(n_345), .Y(n_315) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_316), .B(n_459), .C(n_462), .Y(n_458) );
AOI33xp33_ASAP7_75t_L g530 ( .A1(n_316), .A2(n_531), .A3(n_533), .B1(n_538), .B2(n_543), .B3(n_545), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_316), .B(n_673), .C(n_674), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_316), .B(n_847), .C(n_849), .Y(n_846) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_316), .B(n_885), .C(n_886), .Y(n_884) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI22xp5_ASAP7_75t_SL g918 ( .A1(n_317), .A2(n_747), .B1(n_919), .B2(n_925), .Y(n_918) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_318), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g368 ( .A(n_318), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g606 ( .A(n_318), .B(n_369), .Y(n_606) );
OR2x6_ASAP7_75t_L g621 ( .A(n_318), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g788 ( .A(n_318), .B(n_622), .Y(n_788) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g622 ( .A(n_320), .Y(n_622) );
INVx1_ASAP7_75t_L g741 ( .A(n_322), .Y(n_741) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_SL g357 ( .A(n_326), .Y(n_357) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_327), .Y(n_433) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g385 ( .A(n_330), .B(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_330), .Y(n_451) );
BUFx2_ASAP7_75t_L g553 ( .A(n_330), .Y(n_553) );
INVx1_ASAP7_75t_L g566 ( .A(n_330), .Y(n_566) );
INVx1_ASAP7_75t_L g617 ( .A(n_330), .Y(n_617) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_330), .Y(n_718) );
BUFx2_ASAP7_75t_L g729 ( .A(n_330), .Y(n_729) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_SL g731 ( .A(n_334), .Y(n_731) );
BUFx3_ASAP7_75t_L g774 ( .A(n_334), .Y(n_774) );
INVx2_ASAP7_75t_SL g1258 ( .A(n_334), .Y(n_1258) );
INVx4_ASAP7_75t_L g1264 ( .A(n_334), .Y(n_1264) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g391 ( .A(n_335), .Y(n_391) );
INVx3_ASAP7_75t_L g454 ( .A(n_335), .Y(n_454) );
INVx1_ASAP7_75t_L g557 ( .A(n_335), .Y(n_557) );
AND2x4_ASAP7_75t_L g343 ( .A(n_336), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_SL g367 ( .A(n_339), .Y(n_367) );
INVx2_ASAP7_75t_L g667 ( .A(n_339), .Y(n_667) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g456 ( .A(n_340), .Y(n_456) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g561 ( .A(n_341), .Y(n_561) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_342), .Y(n_373) );
INVx2_ASAP7_75t_SL g734 ( .A(n_342), .Y(n_734) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g374 ( .A(n_343), .B(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g412 ( .A(n_343), .Y(n_412) );
INVx1_ASAP7_75t_L g448 ( .A(n_343), .Y(n_448) );
BUFx3_ASAP7_75t_L g457 ( .A(n_343), .Y(n_457) );
BUFx2_ASAP7_75t_L g524 ( .A(n_343), .Y(n_524) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_343), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_345), .B(n_450), .C(n_455), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_345), .B(n_669), .C(n_671), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_345), .B(n_842), .C(n_845), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_345), .B(n_882), .C(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g917 ( .A(n_345), .Y(n_917) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x6_ASAP7_75t_L g549 ( .A(n_347), .B(n_550), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
AOI33xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .A3(n_360), .B1(n_365), .B2(n_366), .B3(n_368), .Y(n_351) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_352), .B(n_467), .C(n_472), .Y(n_466) );
AOI33xp33_ASAP7_75t_L g619 ( .A1(n_352), .A2(n_620), .A3(n_623), .B1(n_626), .B2(n_627), .B3(n_631), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_352), .B(n_677), .C(n_679), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_352), .B(n_852), .C(n_853), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_352), .B(n_888), .C(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g970 ( .A(n_352), .Y(n_970) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x4_ASAP7_75t_L g532 ( .A(n_353), .B(n_354), .Y(n_532) );
INVx1_ASAP7_75t_L g1241 ( .A(n_358), .Y(n_1241) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g544 ( .A(n_359), .Y(n_544) );
INVx2_ASAP7_75t_SL g750 ( .A(n_361), .Y(n_750) );
BUFx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g542 ( .A(n_363), .Y(n_542) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_368), .B(n_445), .C(n_446), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g547 ( .A1(n_368), .A2(n_548), .A3(n_552), .B1(n_558), .B2(n_564), .B3(n_570), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_368), .B(n_664), .C(n_666), .Y(n_663) );
INVx2_ASAP7_75t_L g726 ( .A(n_368), .Y(n_726) );
BUFx3_ASAP7_75t_L g779 ( .A(n_368), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_368), .B(n_839), .C(n_840), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g878 ( .A(n_368), .B(n_879), .C(n_880), .Y(n_878) );
AOI31xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_384), .A3(n_393), .B(n_398), .Y(n_370) );
AOI211xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_374), .C(n_377), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_373), .A2(n_414), .B1(n_486), .B2(n_696), .C1(n_697), .C2(n_698), .Y(n_695) );
CKINVDCx11_ASAP7_75t_R g424 ( .A(n_374), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_374), .A2(n_447), .B(n_597), .C(n_598), .Y(n_596) );
AOI211xp5_ASAP7_75t_L g829 ( .A1(n_374), .A2(n_803), .B(n_830), .C(n_831), .Y(n_829) );
AOI211xp5_ASAP7_75t_L g869 ( .A1(n_374), .A2(n_608), .B(n_870), .C(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
INVx2_ASAP7_75t_L g485 ( .A(n_379), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g802 ( .A1(n_379), .A2(n_486), .B1(n_767), .B2(n_768), .C1(n_797), .C2(n_803), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_379), .A2(n_486), .B1(n_937), .B2(n_938), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_379), .A2(n_486), .B1(n_988), .B2(n_989), .Y(n_993) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g481 ( .A(n_383), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_383), .B(n_482), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_388), .B1(n_389), .B2(n_392), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_385), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_385), .A2(n_408), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_385), .A2(n_408), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_385), .A2(n_389), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_385), .A2(n_423), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_385), .A2(n_394), .B1(n_833), .B2(n_834), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_385), .A2(n_394), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_385), .A2(n_389), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AND2x4_ASAP7_75t_L g389 ( .A(n_386), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g408 ( .A(n_386), .B(n_390), .Y(n_408) );
INVx1_ASAP7_75t_L g808 ( .A(n_386), .Y(n_808) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_389), .A2(n_394), .B1(n_700), .B2(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_391), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_394), .A2(n_423), .B1(n_514), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_394), .A2(n_396), .B1(n_588), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_394), .A2(n_396), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_394), .A2(n_423), .B1(n_796), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_394), .A2(n_396), .B1(n_1236), .B2(n_1253), .Y(n_1252) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_396), .A2(n_408), .B1(n_821), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_396), .A2(n_408), .B1(n_860), .B2(n_876), .Y(n_875) );
INVx5_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
AOI31xp33_ASAP7_75t_L g593 ( .A1(n_398), .A2(n_594), .A3(n_596), .B(n_600), .Y(n_593) );
AOI31xp33_ASAP7_75t_L g828 ( .A1(n_398), .A2(n_829), .A3(n_832), .B(n_835), .Y(n_828) );
AOI31xp33_ASAP7_75t_L g868 ( .A1(n_398), .A2(n_869), .A3(n_872), .B(n_875), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_498), .B1(n_576), .B2(n_577), .Y(n_401) );
INVx1_ASAP7_75t_L g576 ( .A(n_402), .Y(n_576) );
AOI221x1_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_425), .B1(n_427), .B2(n_440), .C(n_442), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .C(n_420), .D(n_424), .Y(n_404) );
INVx1_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
INVx5_ASAP7_75t_SL g811 ( .A(n_408), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_413), .B2(n_414), .C1(n_416), .C2(n_417), .Y(n_409) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g574 ( .A(n_412), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_413), .A2(n_416), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_414), .A2(n_417), .B1(n_521), .B2(n_522), .C1(n_525), .C2(n_526), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g1249 ( .A1(n_414), .A2(n_486), .B1(n_1242), .B2(n_1243), .C1(n_1250), .C2(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_417), .A2(n_484), .B1(n_524), .B2(n_646), .C1(n_647), .C2(n_648), .Y(n_645) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x4_ASAP7_75t_L g486 ( .A(n_418), .B(n_419), .Y(n_486) );
INVx1_ASAP7_75t_L g476 ( .A(n_420), .Y(n_476) );
NAND4xp25_ASAP7_75t_SL g516 ( .A(n_424), .B(n_517), .C(n_520), .D(n_527), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_424), .B(n_642), .C(n_645), .D(n_649), .Y(n_641) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_424), .B(n_692), .C(n_695), .D(n_699), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_424), .B(n_802), .C(n_804), .Y(n_801) );
NAND4xp25_ASAP7_75t_SL g1245 ( .A(n_424), .B(n_1246), .C(n_1249), .D(n_1252), .Y(n_1245) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_425), .A2(n_476), .A3(n_477), .B(n_487), .Y(n_475) );
AOI221x1_ASAP7_75t_L g500 ( .A1(n_425), .A2(n_440), .B1(n_501), .B2(n_516), .C(n_529), .Y(n_500) );
AOI221x1_ASAP7_75t_L g640 ( .A1(n_425), .A2(n_441), .B1(n_641), .B2(n_652), .C(n_662), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_425), .A2(n_691), .B1(n_702), .B2(n_711), .C(n_713), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_425), .A2(n_801), .B(n_806), .Y(n_800) );
OAI31xp33_ASAP7_75t_SL g940 ( .A1(n_425), .A2(n_941), .A3(n_942), .B(n_946), .Y(n_940) );
OAI31xp33_ASAP7_75t_SL g990 ( .A1(n_425), .A2(n_991), .A3(n_992), .B(n_994), .Y(n_990) );
AOI221x1_ASAP7_75t_L g1230 ( .A1(n_425), .A2(n_440), .B1(n_1231), .B2(n_1245), .C(n_1254), .Y(n_1230) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .C(n_437), .D(n_439), .Y(n_427) );
INVxp67_ASAP7_75t_L g489 ( .A(n_428), .Y(n_489) );
BUFx4f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_439), .B(n_703), .C(n_706), .D(n_708), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g818 ( .A(n_439), .B(n_819), .C(n_822), .D(n_825), .Y(n_818) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_439), .B(n_858), .C(n_861), .D(n_864), .Y(n_857) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_439), .Y(n_1244) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_440), .A2(n_489), .A3(n_490), .B(n_497), .Y(n_488) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI211x1_ASAP7_75t_SL g581 ( .A1(n_441), .A2(n_582), .B(n_593), .C(n_603), .Y(n_581) );
INVx1_ASAP7_75t_L g712 ( .A(n_441), .Y(n_712) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_443), .B(n_475), .C(n_488), .Y(n_474) );
AND4x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_449), .C(n_458), .D(n_466), .Y(n_443) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g665 ( .A(n_453), .Y(n_665) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g613 ( .A(n_454), .Y(n_613) );
INVx3_ASAP7_75t_L g721 ( .A(n_454), .Y(n_721) );
BUFx2_ASAP7_75t_L g803 ( .A(n_457), .Y(n_803) );
INVx1_ASAP7_75t_L g753 ( .A(n_461), .Y(n_753) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g1270 ( .A(n_469), .Y(n_1270) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_480), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_775) );
OAI22xp33_ASAP7_75t_SL g781 ( .A1(n_480), .A2(n_782), .B1(n_783), .B2(n_785), .Y(n_781) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_480), .A2(n_973), .B1(n_981), .B2(n_982), .Y(n_980) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g915 ( .A(n_481), .Y(n_915) );
BUFx2_ASAP7_75t_L g944 ( .A(n_481), .Y(n_944) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g508 ( .A(n_492), .Y(n_508) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g793 ( .A(n_493), .Y(n_793) );
INVx1_ASAP7_75t_L g923 ( .A(n_493), .Y(n_923) );
BUFx2_ASAP7_75t_L g929 ( .A(n_493), .Y(n_929) );
BUFx4f_ASAP7_75t_L g962 ( .A(n_493), .Y(n_962) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OR2x2_ASAP7_75t_L g761 ( .A(n_494), .B(n_495), .Y(n_761) );
INVx2_ASAP7_75t_L g577 ( .A(n_498), .Y(n_577) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .C(n_513), .Y(n_501) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g867 ( .A(n_505), .Y(n_867) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g1251 ( .A(n_523), .Y(n_1251) );
INVx1_ASAP7_75t_L g1260 ( .A(n_523), .Y(n_1260) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_547), .Y(n_529) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g747 ( .A(n_532), .Y(n_747) );
BUFx4f_ASAP7_75t_L g1282 ( .A(n_532), .Y(n_1282) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g936 ( .A(n_537), .Y(n_936) );
BUFx4f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g953 ( .A(n_540), .Y(n_953) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI33xp33_ASAP7_75t_L g604 ( .A1(n_548), .A2(n_605), .A3(n_607), .B1(n_610), .B2(n_614), .B3(n_615), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_548), .B(n_728), .C(n_732), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g1261 ( .A(n_548), .B(n_1262), .C(n_1265), .Y(n_1261) );
INVx5_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx6_ASAP7_75t_L g786 ( .A(n_549), .Y(n_786) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g569 ( .A(n_557), .Y(n_569) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g572 ( .A(n_561), .Y(n_572) );
INVx2_ASAP7_75t_L g724 ( .A(n_561), .Y(n_724) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g609 ( .A(n_563), .Y(n_609) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g1267 ( .A(n_572), .Y(n_1267) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g684 ( .A(n_578), .Y(n_684) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_638), .B1(n_639), .B2(n_683), .Y(n_579) );
INVx1_ASAP7_75t_L g683 ( .A(n_580), .Y(n_683) );
INVx1_ASAP7_75t_L g637 ( .A(n_581), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_619), .Y(n_603) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g618 ( .A(n_612), .Y(n_618) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g908 ( .A(n_613), .Y(n_908) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g670 ( .A(n_617), .Y(n_670) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_621), .Y(n_744) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g850 ( .A(n_633), .Y(n_850) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g682 ( .A(n_640), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .C(n_659), .Y(n_652) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_668), .C(n_672), .D(n_676), .Y(n_662) );
INVx2_ASAP7_75t_L g1273 ( .A(n_675), .Y(n_1273) );
BUFx2_ASAP7_75t_L g710 ( .A(n_678), .Y(n_710) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_812), .Y(n_686) );
XNOR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_754), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_689), .A2(n_1003), .B1(n_1024), .B2(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_727), .C(n_735), .D(n_745), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_722), .C(n_725), .Y(n_714) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g911 ( .A(n_721), .Y(n_911) );
BUFx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_725), .B(n_1256), .C(n_1259), .Y(n_1255) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .C(n_744), .Y(n_735) );
BUFx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_741), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_744), .B(n_1269), .C(n_1271), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .C(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g787 ( .A1(n_747), .A2(n_788), .B1(n_789), .B2(n_795), .Y(n_787) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
XNOR2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND3x1_ASAP7_75t_SL g756 ( .A(n_757), .B(n_772), .C(n_800), .Y(n_756) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx2_ASAP7_75t_L g791 ( .A(n_761), .Y(n_791) );
INVx1_ASAP7_75t_L g959 ( .A(n_761), .Y(n_959) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_765), .A2(n_823), .B(n_824), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_765), .A2(n_865), .B(n_866), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_779), .B1(n_780), .B2(n_786), .C(n_787), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_776), .A2(n_778), .B1(n_790), .B2(n_792), .C(n_794), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_777), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_913) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_788), .A2(n_951), .A3(n_956), .B1(n_963), .B2(n_966), .B3(n_970), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g795 ( .A1(n_790), .A2(n_792), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_795) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g920 ( .A(n_791), .Y(n_920) );
INVx2_ASAP7_75t_L g926 ( .A(n_791), .Y(n_926) );
BUFx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g955 ( .A(n_799), .Y(n_955) );
OR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g906 ( .A(n_810), .Y(n_906) );
XOR2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_890), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_854), .B2(n_855), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g837 ( .A(n_838), .B(n_841), .C(n_846), .D(n_851), .Y(n_837) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_881), .C(n_884), .D(n_887), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_947), .B1(n_995), .B2(n_996), .Y(n_890) );
INVx1_ASAP7_75t_L g995 ( .A(n_891), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_932), .C(n_940), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_918), .Y(n_893) );
OAI33xp33_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_897), .A3(n_903), .B1(n_909), .B2(n_913), .B3(n_917), .Y(n_894) );
OAI33xp33_ASAP7_75t_L g971 ( .A1(n_895), .A2(n_917), .A3(n_972), .B1(n_975), .B2(n_976), .B3(n_980), .Y(n_971) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_899), .B1(n_900), .B2(n_902), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g919 ( .A1(n_899), .A2(n_902), .B1(n_920), .B2(n_921), .C(n_924), .Y(n_919) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_900), .A2(n_957), .B1(n_960), .B2(n_973), .Y(n_972) );
BUFx6f_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp33_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_905), .B1(n_907), .B2(n_908), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_905), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_905), .A2(n_911), .B1(n_952), .B2(n_954), .Y(n_975) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g977 ( .A(n_906), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_911), .A2(n_977), .B1(n_978), .B2(n_979), .Y(n_976) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_928), .B2(n_930), .C(n_931), .Y(n_925) );
INVx2_ASAP7_75t_SL g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g996 ( .A(n_947), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_983), .C(n_990), .Y(n_948) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_971), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B1(n_960), .B2(n_961), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_958), .A2(n_961), .B1(n_964), .B2(n_965), .Y(n_963) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g1274 ( .A(n_968), .Y(n_1274) );
INVx1_ASAP7_75t_L g1281 ( .A(n_968), .Y(n_1281) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1008), .B(n_1225), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
BUFx2_ASAP7_75t_SL g999 ( .A(n_1000), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_1000), .A2(n_1113), .B1(n_1114), .B2(n_1115), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_1001), .A2(n_1023), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1021 ( .A1(n_1003), .A2(n_1022), .B1(n_1023), .B2(n_1026), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_1003), .A2(n_1023), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1004), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1005), .B(n_1018), .Y(n_1025) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_1007), .B(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1007), .Y(n_1031) );
NOR2x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1162), .Y(n_1008) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1100), .C(n_1123), .Y(n_1009) );
AOI211xp5_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1036), .B(n_1064), .C(n_1092), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1011), .B(n_1083), .Y(n_1165) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_1012), .A2(n_1027), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1027), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_1013), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1013), .B(n_1049), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1013), .B(n_1027), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1013 ( .A(n_1014), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_1014), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1014), .B(n_1027), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1014), .B(n_1027), .Y(n_1144) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1015), .Y(n_1078) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1015), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1019), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1016), .B(n_1019), .Y(n_1035) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_1017), .B(n_1019), .Y(n_1020) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1020), .Y(n_1053) );
INVx1_ASAP7_75t_SL g1059 ( .A(n_1020), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_1023), .Y(n_1114) );
BUFx6f_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1025), .Y(n_1030) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1027), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1027), .B(n_1071), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1027), .B(n_1071), .Y(n_1120) );
OAI21xp33_ASAP7_75t_L g1124 ( .A1(n_1027), .A2(n_1125), .B(n_1127), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1027), .B(n_1072), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1034), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_1031), .B(n_1033), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1295 ( .A(n_1033), .Y(n_1295) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1035), .Y(n_1057) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1047), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1038), .B(n_1146), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_1038), .B(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1039), .B(n_1054), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1039), .B(n_1055), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1040), .B(n_1044), .Y(n_1067) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1040), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1040), .B(n_1055), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1040), .B(n_1044), .Y(n_1184) );
NOR2xp33_ASAP7_75t_SL g1214 ( .A(n_1040), .B(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_1043), .B(n_1054), .Y(n_1085) );
NOR3xp33_ASAP7_75t_L g1105 ( .A(n_1043), .B(n_1083), .C(n_1106), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1043), .B(n_1054), .Y(n_1135) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1044), .B(n_1054), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1044), .B(n_1098), .Y(n_1097) );
OAI322xp33_ASAP7_75t_L g1168 ( .A1(n_1044), .A2(n_1169), .A3(n_1172), .B1(n_1173), .B2(n_1175), .C1(n_1177), .C2(n_1179), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1178 ( .A(n_1044), .B(n_1054), .Y(n_1178) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1054), .Y(n_1048) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1049), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1049), .B(n_1054), .Y(n_1099) );
INVx4_ASAP7_75t_L g1104 ( .A(n_1049), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1049), .B(n_1134), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1049), .B(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1049), .B(n_1174), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1049), .B(n_1072), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1049), .B(n_1088), .Y(n_1215) );
AND2x6_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_1053), .A2(n_1109), .B1(n_1110), .B2(n_1111), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1054), .B(n_1067), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1054), .B(n_1103), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1054), .B(n_1097), .Y(n_1158) );
CKINVDCx6p67_ASAP7_75t_R g1054 ( .A(n_1055), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1055), .B(n_1103), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1055), .B(n_1097), .Y(n_1138) );
AOI32xp33_ASAP7_75t_L g1140 ( .A1(n_1055), .A2(n_1119), .A3(n_1141), .B1(n_1145), .B2(n_1147), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1055), .B(n_1067), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1055), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1055), .B(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1055), .B(n_1219), .Y(n_1218) );
OR2x6_ASAP7_75t_SL g1055 ( .A(n_1056), .B(n_1061), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1059), .A2(n_1077), .B1(n_1078), .B2(n_1079), .Y(n_1076) );
OAI221xp5_ASAP7_75t_L g1064 ( .A1(n_1065), .A2(n_1068), .B1(n_1081), .B2(n_1086), .C(n_1089), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1067), .B(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1067), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1069), .Y(n_1197) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1069), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1070), .B(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1080), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1071), .B(n_1088), .Y(n_1087) );
INVx3_ASAP7_75t_L g1132 ( .A(n_1071), .Y(n_1132) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1071), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1071), .B(n_1116), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1071), .B(n_1107), .Y(n_1172) );
INVx3_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1072), .B(n_1144), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1076), .Y(n_1072) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NOR2x1_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1085), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1083), .B(n_1138), .Y(n_1137) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1083), .B(n_1190), .Y(n_1189) );
NOR2x1_ASAP7_75t_R g1205 ( .A(n_1083), .B(n_1146), .Y(n_1205) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1084), .B(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1084), .B(n_1134), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1084), .B(n_1150), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1084), .B(n_1138), .Y(n_1223) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1085), .Y(n_1152) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
AOI322xp5_ASAP7_75t_L g1151 ( .A1(n_1087), .A2(n_1132), .A3(n_1152), .B1(n_1153), .B2(n_1155), .C1(n_1156), .C2(n_1158), .Y(n_1151) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1088), .Y(n_1094) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1088), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1088), .B(n_1155), .Y(n_1176) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1088), .Y(n_1192) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1096), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1095), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1099), .Y(n_1096) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1097), .Y(n_1146) );
AOI211xp5_ASAP7_75t_L g1200 ( .A1(n_1098), .A2(n_1201), .B(n_1202), .C(n_1205), .Y(n_1200) );
O2A1O1Ixp33_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1105), .B(n_1116), .C(n_1117), .Y(n_1100) );
INVxp67_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1104), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1104), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1104), .B(n_1184), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1104), .B(n_1143), .Y(n_1221) );
OAI31xp33_ASAP7_75t_L g1123 ( .A1(n_1106), .A2(n_1124), .A3(n_1136), .B(n_1139), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_1106), .A2(n_1144), .B1(n_1211), .B2(n_1216), .C(n_1220), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_1107), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1107), .A2(n_1186), .B1(n_1195), .B2(n_1196), .Y(n_1185) );
OR2x6_ASAP7_75t_SL g1107 ( .A(n_1108), .B(n_1112), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1116), .B(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1121), .Y(n_1118) );
AOI322xp5_ASAP7_75t_L g1211 ( .A1(n_1119), .A2(n_1132), .A3(n_1135), .B1(n_1170), .B2(n_1171), .C1(n_1212), .C2(n_1214), .Y(n_1211) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1121), .B(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1122), .Y(n_1148) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
OAI21xp5_ASAP7_75t_SL g1127 ( .A1(n_1128), .A2(n_1130), .B(n_1135), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1129), .B(n_1150), .Y(n_1149) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1133), .Y(n_1130) );
INVx1_ASAP7_75t_SL g1131 ( .A(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1132), .B(n_1137), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1132), .B(n_1158), .Y(n_1194) );
AOI21xp5_ASAP7_75t_L g1193 ( .A1(n_1133), .A2(n_1146), .B(n_1187), .Y(n_1193) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1133), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1135), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1138), .Y(n_1167) );
NAND3xp33_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1151), .C(n_1159), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1143), .B(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1148), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1150), .Y(n_1187) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
A2O1A1Ixp33_ASAP7_75t_L g1207 ( .A1(n_1154), .A2(n_1167), .B(n_1183), .C(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1155), .Y(n_1190) );
AOI211xp5_ASAP7_75t_SL g1206 ( .A1(n_1155), .A2(n_1207), .B(n_1210), .C(n_1222), .Y(n_1206) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1157), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1158), .B(n_1178), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1158), .B(n_1192), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1158), .B(n_1209), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
AOI211xp5_ASAP7_75t_L g1188 ( .A1(n_1160), .A2(n_1189), .B(n_1191), .C(n_1193), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1185), .C(n_1206), .Y(n_1162) );
AOI211xp5_ASAP7_75t_SL g1163 ( .A1(n_1164), .A2(n_1166), .B(n_1168), .C(n_1181), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g1164 ( .A(n_1165), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1196 ( .A1(n_1167), .A2(n_1197), .B(n_1198), .C(n_1200), .Y(n_1196) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1172), .Y(n_1195) );
OAI211xp5_ASAP7_75t_L g1186 ( .A1(n_1175), .A2(n_1187), .B(n_1188), .C(n_1194), .Y(n_1186) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1184), .Y(n_1213) );
AOI21xp5_ASAP7_75t_L g1222 ( .A1(n_1216), .A2(n_1223), .B(n_1224), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1230), .Y(n_1283) );
NAND4xp25_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .C(n_1238), .D(n_1244), .Y(n_1231) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NAND4xp25_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1261), .C(n_1268), .D(n_1275), .Y(n_1254) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_1273), .Y(n_1272) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1280), .C(n_1282), .Y(n_1275) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
HB1xp67_ASAP7_75t_L g1287 ( .A(n_1283), .Y(n_1287) );
BUFx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1287), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_1292), .Y(n_1291) );
OAI21xp5_ASAP7_75t_L g1294 ( .A1(n_1293), .A2(n_1295), .B(n_1296), .Y(n_1294) );
endmodule