module fake_jpeg_26093_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_5),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_3),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_17),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_17),
.C(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_20),
.C(n_23),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_22),
.B(n_18),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_35),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_40),
.C(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_40),
.Y(n_43)
);


endmodule