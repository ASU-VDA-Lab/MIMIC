module real_aes_16774_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g848 ( .A(n_0), .B(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_1), .A2(n_3), .B1(n_172), .B2(n_499), .Y(n_498) );
OAI22x1_ASAP7_75t_R g108 ( .A1(n_2), .A2(n_46), .B1(n_109), .B2(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_4), .A2(n_44), .B1(n_129), .B2(n_152), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_5), .A2(n_27), .B1(n_152), .B2(n_228), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_6), .A2(n_16), .B1(n_171), .B2(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_7), .A2(n_62), .B1(n_189), .B2(n_230), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_8), .A2(n_17), .B1(n_128), .B2(n_129), .Y(n_515) );
INVx1_ASAP7_75t_L g849 ( .A(n_9), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_10), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_11), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_12), .A2(n_19), .B1(n_188), .B2(n_191), .Y(n_187) );
OR2x2_ASAP7_75t_L g803 ( .A(n_13), .B(n_41), .Y(n_803) );
BUFx2_ASAP7_75t_L g854 ( .A(n_13), .Y(n_854) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_14), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_15), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_18), .A2(n_829), .B(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g822 ( .A(n_20), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_21), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_22), .A2(n_102), .B1(n_171), .B2(n_172), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_23), .A2(n_40), .B1(n_137), .B2(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_24), .B(n_132), .Y(n_131) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_25), .A2(n_58), .B(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_26), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_26), .A2(n_80), .B1(n_478), .B2(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_28), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_29), .B(n_134), .Y(n_485) );
INVx4_ASAP7_75t_R g527 ( .A(n_30), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_31), .A2(n_49), .B1(n_157), .B2(n_158), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_32), .A2(n_55), .B1(n_158), .B2(n_171), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_33), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_34), .B(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_35), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_36), .B(n_152), .Y(n_492) );
INVx1_ASAP7_75t_L g501 ( .A(n_37), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_SL g567 ( .A1(n_38), .A2(n_129), .B(n_133), .C(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_39), .A2(n_56), .B1(n_129), .B2(n_158), .Y(n_474) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_41), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_42), .A2(n_90), .B1(n_129), .B2(n_227), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_43), .A2(n_48), .B1(n_128), .B2(n_129), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_45), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_47), .A2(n_61), .B1(n_171), .B2(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g489 ( .A(n_50), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_51), .B(n_129), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_52), .Y(n_548) );
INVx2_ASAP7_75t_L g798 ( .A(n_53), .Y(n_798) );
BUFx3_ASAP7_75t_L g801 ( .A(n_54), .Y(n_801) );
INVx1_ASAP7_75t_L g818 ( .A(n_54), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_57), .A2(n_91), .B1(n_129), .B2(n_158), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_59), .Y(n_528) );
AOI22x1_ASAP7_75t_SL g789 ( .A1(n_60), .A2(n_69), .B1(n_790), .B2(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_60), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_63), .A2(n_78), .B1(n_157), .B2(n_175), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_64), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_65), .A2(n_81), .B1(n_128), .B2(n_129), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_66), .A2(n_100), .B1(n_171), .B2(n_191), .Y(n_217) );
INVx1_ASAP7_75t_L g124 ( .A(n_67), .Y(n_124) );
AND2x4_ASAP7_75t_L g143 ( .A(n_68), .B(n_144), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_69), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_70), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_70), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_71), .A2(n_93), .B1(n_157), .B2(n_158), .Y(n_497) );
AO22x1_ASAP7_75t_L g506 ( .A1(n_72), .A2(n_79), .B1(n_204), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g144 ( .A(n_73), .Y(n_144) );
AND2x2_ASAP7_75t_L g570 ( .A(n_74), .B(n_146), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_75), .B(n_230), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_76), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_77), .A2(n_105), .B1(n_840), .B2(n_855), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g811 ( .A(n_80), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_82), .B(n_152), .Y(n_549) );
INVx2_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_84), .B(n_146), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_85), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_86), .A2(n_101), .B1(n_158), .B2(n_230), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_87), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_88), .B(n_179), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_89), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_92), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_94), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_95), .B(n_146), .Y(n_545) );
INVx1_ASAP7_75t_L g461 ( .A(n_96), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_96), .B(n_817), .Y(n_816) );
NAND2xp33_ASAP7_75t_L g139 ( .A(n_97), .B(n_132), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_98), .A2(n_194), .B(n_230), .C(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g529 ( .A(n_99), .B(n_530), .Y(n_529) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_103), .B(n_138), .Y(n_553) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_794), .B(n_804), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_789), .B1(n_792), .B2(n_793), .Y(n_106) );
INVx2_ASAP7_75t_L g792 ( .A(n_107), .Y(n_792) );
XNOR2x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_458), .B1(n_462), .B2(n_786), .Y(n_111) );
XNOR2x1_ASAP7_75t_SL g819 ( .A(n_112), .B(n_820), .Y(n_819) );
NAND2x1p5_ASAP7_75t_L g112 ( .A(n_113), .B(n_402), .Y(n_112) );
NOR3x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_320), .C(n_357), .Y(n_113) );
NAND4xp75_ASAP7_75t_L g114 ( .A(n_115), .B(n_240), .C(n_274), .D(n_304), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI32xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_162), .A3(n_212), .B1(n_221), .B2(n_235), .Y(n_116) );
OR2x2_ASAP7_75t_L g221 ( .A(n_117), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_118), .A2(n_432), .B(n_434), .Y(n_431) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_147), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_119), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g303 ( .A(n_119), .B(n_249), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_119), .B(n_214), .Y(n_398) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g247 ( .A(n_120), .Y(n_247) );
OAI21x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_145), .Y(n_120) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_121), .A2(n_125), .B(n_145), .Y(n_280) );
INVx2_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx4_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_122), .B(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g209 ( .A(n_122), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_122), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_122), .B(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g493 ( .A(n_122), .B(n_476), .Y(n_493) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g179 ( .A(n_123), .Y(n_179) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_135), .B(n_141), .Y(n_125) );
O2A1O1Ixp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_131), .C(n_133), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_128), .A2(n_548), .B(n_549), .C(n_550), .Y(n_547) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
INVx1_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_130), .Y(n_132) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_130), .Y(n_152) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
INVx1_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
INVx2_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
INVx1_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
INVx3_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_132), .Y(n_507) );
INVx6_ASAP7_75t_L g140 ( .A(n_133), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_133), .A2(n_506), .B(n_508), .C(n_511), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_133), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_133), .B(n_506), .Y(n_579) );
BUFx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
INVx1_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
INVx1_ASAP7_75t_L g488 ( .A(n_134), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_140), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_138), .A2(n_208), .B1(n_527), .B2(n_528), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_140), .A2(n_151), .B1(n_153), .B2(n_156), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_140), .A2(n_153), .B1(n_170), .B2(n_174), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_140), .A2(n_187), .B1(n_192), .B2(n_193), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_140), .A2(n_153), .B1(n_203), .B2(n_206), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_140), .A2(n_193), .B1(n_217), .B2(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_140), .A2(n_226), .B1(n_229), .B2(n_231), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_140), .A2(n_153), .B1(n_265), .B2(n_266), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_140), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_140), .A2(n_231), .B1(n_497), .B2(n_498), .Y(n_496) );
OAI22x1_ASAP7_75t_L g514 ( .A1(n_140), .A2(n_231), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_SL g232 ( .A(n_142), .Y(n_232) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx10_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
BUFx10_ASAP7_75t_L g476 ( .A(n_143), .Y(n_476) );
INVx1_ASAP7_75t_L g512 ( .A(n_143), .Y(n_512) );
INVx2_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_146), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g271 ( .A(n_147), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_147), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_148), .Y(n_258) );
INVx1_ASAP7_75t_L g302 ( .A(n_148), .Y(n_302) );
AND2x2_ASAP7_75t_L g346 ( .A(n_148), .B(n_280), .Y(n_346) );
OR2x2_ASAP7_75t_L g400 ( .A(n_148), .B(n_224), .Y(n_400) );
AO31x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .A3(n_159), .B(n_160), .Y(n_148) );
INVx2_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
AO31x2_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_186), .A3(n_195), .B(n_197), .Y(n_185) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_149), .A2(n_202), .A3(n_209), .B(n_210), .Y(n_201) );
AO31x2_ASAP7_75t_L g513 ( .A1(n_149), .A2(n_182), .A3(n_514), .B(n_517), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_152), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g475 ( .A(n_154), .Y(n_475) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g551 ( .A(n_155), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_158), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g499 ( .A(n_158), .Y(n_499) );
AO31x2_ASAP7_75t_L g471 ( .A1(n_159), .A2(n_472), .A3(n_476), .B(n_477), .Y(n_471) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_163), .A2(n_326), .B1(n_418), .B2(n_420), .Y(n_417) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_183), .Y(n_163) );
INVx4_ASAP7_75t_L g243 ( .A(n_164), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_164), .A2(n_223), .B1(n_255), .B2(n_257), .Y(n_254) );
OR2x2_ASAP7_75t_L g260 ( .A(n_164), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g379 ( .A(n_164), .B(n_278), .Y(n_379) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g299 ( .A(n_165), .B(n_184), .Y(n_299) );
AND2x2_ASAP7_75t_L g390 ( .A(n_165), .B(n_262), .Y(n_390) );
AND2x2_ASAP7_75t_L g445 ( .A(n_165), .B(n_201), .Y(n_445) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
AND2x4_ASAP7_75t_L g366 ( .A(n_166), .B(n_262), .Y(n_366) );
AO31x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .A3(n_176), .B(n_180), .Y(n_166) );
AO31x2_ASAP7_75t_L g215 ( .A1(n_167), .A2(n_195), .A3(n_216), .B(n_219), .Y(n_215) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_168), .A2(n_522), .B(n_525), .Y(n_521) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_173), .B(n_565), .Y(n_564) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_176), .A2(n_232), .A3(n_264), .B(n_267), .Y(n_263) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_176), .A2(n_521), .B(n_529), .Y(n_520) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_178), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_178), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g182 ( .A(n_179), .Y(n_182) );
INVx2_ASAP7_75t_L g196 ( .A(n_179), .Y(n_196) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_179), .A2(n_510), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_182), .B(n_268), .Y(n_267) );
NAND2x1_ASAP7_75t_L g242 ( .A(n_183), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_183), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
INVx2_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_184), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g285 ( .A(n_184), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_184), .B(n_287), .Y(n_312) );
AND2x2_ASAP7_75t_L g315 ( .A(n_184), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g375 ( .A(n_184), .Y(n_375) );
INVx4_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_185), .B(n_200), .Y(n_253) );
BUFx2_ASAP7_75t_L g291 ( .A(n_185), .Y(n_291) );
AND2x2_ASAP7_75t_L g340 ( .A(n_185), .B(n_201), .Y(n_340) );
AND2x2_ASAP7_75t_L g382 ( .A(n_185), .B(n_263), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_185), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_190), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
AO31x2_ASAP7_75t_L g495 ( .A1(n_195), .A2(n_232), .A3(n_496), .B(n_500), .Y(n_495) );
AOI21x1_ASAP7_75t_L g559 ( .A1(n_195), .A2(n_560), .B(n_570), .Y(n_559) );
BUFx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_196), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_196), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_196), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g530 ( .A(n_196), .Y(n_530) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_201), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g293 ( .A(n_201), .B(n_263), .Y(n_293) );
INVx1_ASAP7_75t_L g316 ( .A(n_201), .Y(n_316) );
INVx2_ASAP7_75t_L g336 ( .A(n_201), .Y(n_336) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_201), .Y(n_381) );
OAI21xp33_ASAP7_75t_SL g484 ( .A1(n_204), .A2(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_209), .A2(n_225), .A3(n_232), .B(n_233), .Y(n_224) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g300 ( .A(n_213), .B(n_301), .Y(n_300) );
NOR2x1p5_ASAP7_75t_L g406 ( .A(n_213), .B(n_400), .Y(n_406) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g223 ( .A(n_214), .B(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_214), .B(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g248 ( .A(n_215), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g306 ( .A(n_215), .B(n_224), .Y(n_306) );
BUFx2_ASAP7_75t_L g419 ( .A(n_215), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_221), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g457 ( .A(n_221), .Y(n_457) );
INVx2_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g393 ( .A(n_223), .Y(n_393) );
AND2x4_ASAP7_75t_L g416 ( .A(n_223), .B(n_346), .Y(n_416) );
AND2x2_ASAP7_75t_L g440 ( .A(n_223), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g249 ( .A(n_224), .Y(n_249) );
BUFx2_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
INVx1_ASAP7_75t_L g329 ( .A(n_224), .Y(n_329) );
OR2x2_ASAP7_75t_L g451 ( .A(n_224), .B(n_308), .Y(n_451) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_228), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_231), .B(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g297 ( .A(n_237), .Y(n_297) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_238), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_238), .Y(n_318) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g259 ( .A(n_239), .Y(n_259) );
OR2x2_ASAP7_75t_L g296 ( .A(n_239), .B(n_288), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B(n_250), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_245), .A2(n_339), .B1(n_341), .B2(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
OR2x2_ASAP7_75t_L g384 ( .A(n_247), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g392 ( .A(n_247), .Y(n_392) );
AND2x2_ASAP7_75t_L g405 ( .A(n_247), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g367 ( .A(n_248), .B(n_346), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_254), .B1(n_260), .B2(n_269), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g277 ( .A(n_256), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g345 ( .A(n_256), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g354 ( .A(n_256), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_256), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_257), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g342 ( .A(n_259), .B(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g356 ( .A(n_259), .Y(n_356) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
AND2x4_ASAP7_75t_L g335 ( .A(n_263), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_263), .Y(n_351) );
INVx1_ASAP7_75t_L g415 ( .A(n_263), .Y(n_415) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x4_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
INVx1_ASAP7_75t_L g282 ( .A(n_273), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_283), .B1(n_294), .B2(n_300), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_279), .Y(n_332) );
INVx1_ASAP7_75t_L g308 ( .A(n_280), .Y(n_308) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_289), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_285), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g437 ( .A(n_286), .Y(n_437) );
INVx1_ASAP7_75t_L g456 ( .A(n_286), .Y(n_456) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1_ASAP7_75t_L g433 ( .A(n_290), .B(n_356), .Y(n_433) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g449 ( .A(n_291), .Y(n_449) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx2_ASAP7_75t_L g387 ( .A(n_295), .Y(n_387) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g376 ( .A(n_296), .Y(n_376) );
AND2x4_ASAP7_75t_L g378 ( .A(n_297), .B(n_335), .Y(n_378) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_301), .A2(n_447), .B1(n_450), .B2(n_452), .Y(n_446) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g371 ( .A(n_302), .Y(n_371) );
INVx1_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
AND2x4_ASAP7_75t_L g418 ( .A(n_303), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g426 ( .A(n_303), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
AND2x4_ASAP7_75t_SL g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_SL g369 ( .A(n_306), .Y(n_369) );
INVx2_ASAP7_75t_L g385 ( .A(n_306), .Y(n_385) );
INVx1_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
AND2x2_ASAP7_75t_L g443 ( .A(n_307), .B(n_354), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .C(n_317), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_314), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g355 ( .A(n_315), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_315), .B(n_390), .Y(n_423) );
INVx1_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_318), .B(n_382), .Y(n_408) );
INVx1_ASAP7_75t_L g363 ( .A(n_319), .Y(n_363) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_337), .C(n_347), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_326), .B(n_333), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g441 ( .A(n_324), .Y(n_441) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI32xp33_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_378), .A3(n_379), .B1(n_380), .B2(n_383), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_328), .B(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_335), .B(n_356), .Y(n_396) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_340), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g401 ( .A(n_340), .B(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g429 ( .A(n_343), .Y(n_429) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_345), .A2(n_348), .B1(n_352), .B2(n_355), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_346), .B(n_354), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_348), .A2(n_406), .B1(n_443), .B2(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g444 ( .A(n_350), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_352), .A2(n_395), .B1(n_397), .B2(n_401), .Y(n_394) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g436 ( .A(n_356), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_377), .C(n_386), .D(n_394), .Y(n_357) );
O2A1O1Ixp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_364), .B(n_367), .C(n_368), .Y(n_358) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g422 ( .A(n_366), .B(n_381), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_366), .B(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_373), .A2(n_411), .B1(n_413), .B2(n_416), .Y(n_410) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_378), .A2(n_383), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_391), .Y(n_386) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_R g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_401), .A2(n_418), .B1(n_455), .B2(n_457), .Y(n_454) );
NOR3x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_424), .C(n_438), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_417), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
INVx1_ASAP7_75t_L g427 ( .A(n_419), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_421), .A2(n_425), .B1(n_428), .B2(n_430), .C(n_431), .Y(n_424) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
NAND4xp25_ASAP7_75t_SL g438 ( .A(n_439), .B(n_442), .C(n_446), .D(n_454), .Y(n_438) );
AND2x2_ASAP7_75t_L g452 ( .A(n_445), .B(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_460), .Y(n_788) );
AND2x2_ASAP7_75t_L g838 ( .A(n_460), .B(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g847 ( .A(n_461), .Y(n_847) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_663), .Y(n_463) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_611), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_502), .B(n_531), .C(n_596), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_468), .A2(n_532), .B(n_747), .Y(n_746) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
INVx2_ASAP7_75t_L g592 ( .A(n_469), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_469), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g703 ( .A(n_470), .B(n_481), .Y(n_703) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g571 ( .A(n_471), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_471), .B(n_495), .Y(n_608) );
AND2x2_ASAP7_75t_L g641 ( .A(n_471), .B(n_558), .Y(n_641) );
OR2x2_ASAP7_75t_L g646 ( .A(n_471), .B(n_495), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_475), .A2(n_491), .B(n_492), .Y(n_490) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_475), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g556 ( .A(n_476), .Y(n_556) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g785 ( .A(n_480), .Y(n_785) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_494), .Y(n_480) );
AND2x2_ASAP7_75t_L g586 ( .A(n_481), .B(n_495), .Y(n_586) );
INVx3_ASAP7_75t_L g594 ( .A(n_481), .Y(n_594) );
NAND2x1p5_ASAP7_75t_SL g626 ( .A(n_481), .B(n_610), .Y(n_626) );
INVx1_ASAP7_75t_L g644 ( .A(n_481), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_481), .B(n_589), .Y(n_669) );
BUFx2_ASAP7_75t_L g755 ( .A(n_481), .Y(n_755) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_490), .B(n_493), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
BUFx4f_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g539 ( .A(n_495), .Y(n_539) );
INVx1_ASAP7_75t_L g595 ( .A(n_495), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_495), .B(n_571), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_495), .B(n_558), .Y(n_704) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_519), .Y(n_502) );
INVx1_ASAP7_75t_L g762 ( .A(n_503), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
OR2x2_ASAP7_75t_L g534 ( .A(n_504), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g599 ( .A(n_504), .Y(n_599) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_512), .A2(n_561), .B(n_567), .Y(n_560) );
INVx2_ASAP7_75t_L g535 ( .A(n_513), .Y(n_535) );
OR2x2_ASAP7_75t_L g600 ( .A(n_513), .B(n_520), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_513), .B(n_520), .Y(n_605) );
INVx2_ASAP7_75t_L g650 ( .A(n_513), .Y(n_650) );
AND2x2_ASAP7_75t_L g691 ( .A(n_513), .B(n_544), .Y(n_691) );
AND2x2_ASAP7_75t_L g725 ( .A(n_513), .B(n_622), .Y(n_725) );
INVx1_ASAP7_75t_L g536 ( .A(n_519), .Y(n_536) );
INVx1_ASAP7_75t_L g655 ( .A(n_519), .Y(n_655) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g575 ( .A(n_520), .B(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g616 ( .A(n_520), .B(n_577), .Y(n_616) );
INVx2_ASAP7_75t_L g622 ( .A(n_520), .Y(n_622) );
AND2x2_ASAP7_75t_L g677 ( .A(n_520), .B(n_544), .Y(n_677) );
AND2x2_ASAP7_75t_L g734 ( .A(n_520), .B(n_543), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_537), .B1(n_572), .B2(n_583), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_534), .B(n_713), .C(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g631 ( .A(n_535), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_535), .B(n_543), .Y(n_681) );
INVx1_ASAP7_75t_L g781 ( .A(n_536), .Y(n_781) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_538), .B(n_736), .Y(n_772) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g627 ( .A(n_539), .Y(n_627) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_557), .Y(n_541) );
INVx1_ASAP7_75t_L g615 ( .A(n_542), .Y(n_615) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g695 ( .A(n_543), .B(n_576), .Y(n_695) );
AND2x2_ASAP7_75t_L g714 ( .A(n_543), .B(n_621), .Y(n_714) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
BUFx3_ASAP7_75t_L g620 ( .A(n_544), .Y(n_620) );
AND2x2_ASAP7_75t_L g649 ( .A(n_544), .B(n_650), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_552), .B(n_555), .Y(n_546) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g742 ( .A(n_557), .Y(n_742) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
INVx2_ASAP7_75t_L g610 ( .A(n_558), .Y(n_610) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g589 ( .A(n_559), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B(n_566), .Y(n_561) );
INVx1_ASAP7_75t_L g590 ( .A(n_571), .Y(n_590) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_574), .B(n_581), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g629 ( .A(n_575), .B(n_630), .Y(n_629) );
BUFx2_ASAP7_75t_L g759 ( .A(n_575), .Y(n_759) );
INVx1_ASAP7_75t_L g604 ( .A(n_576), .Y(n_604) );
AND2x2_ASAP7_75t_L g684 ( .A(n_576), .B(n_622), .Y(n_684) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g621 ( .A(n_577), .B(n_622), .Y(n_621) );
AOI21x1_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_582), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g717 ( .A(n_582), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_591), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_584), .A2(n_625), .B1(n_628), .B2(n_632), .Y(n_624) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_585), .A2(n_605), .B1(n_637), .B2(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
BUFx2_ASAP7_75t_SL g623 ( .A(n_586), .Y(n_623) );
AND2x4_ASAP7_75t_L g741 ( .A(n_586), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g750 ( .A(n_586), .Y(n_750) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g662 ( .A(n_588), .Y(n_662) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_589), .B(n_594), .Y(n_720) );
INVxp67_ASAP7_75t_L g749 ( .A(n_589), .Y(n_749) );
AND2x2_ASAP7_75t_L g754 ( .A(n_589), .B(n_620), .Y(n_754) );
OR2x2_ASAP7_75t_L g736 ( .A(n_590), .B(n_610), .Y(n_736) );
INVx1_ASAP7_75t_L g617 ( .A(n_591), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_592), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g656 ( .A(n_593), .B(n_641), .Y(n_656) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_594), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
OR2x2_ASAP7_75t_L g735 ( .A(n_594), .B(n_736), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B(n_606), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g659 ( .A(n_598), .Y(n_659) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g653 ( .A(n_599), .B(n_650), .Y(n_653) );
INVx2_ASAP7_75t_L g777 ( .A(n_599), .Y(n_777) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
AND2x2_ASAP7_75t_L g706 ( .A(n_603), .B(n_649), .Y(n_706) );
AND2x2_ASAP7_75t_L g731 ( .A(n_603), .B(n_677), .Y(n_731) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g634 ( .A(n_604), .Y(n_634) );
AND2x2_ASAP7_75t_L g661 ( .A(n_605), .B(n_615), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_605), .B(n_660), .Y(n_673) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g758 ( .A(n_608), .Y(n_758) );
OR2x2_ASAP7_75t_L g774 ( .A(n_608), .B(n_669), .Y(n_774) );
INVx1_ASAP7_75t_L g698 ( .A(n_610), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_635), .C(n_657), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_617), .B1(n_618), .B2(n_623), .C(n_624), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g637 ( .A(n_616), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_616), .B(n_681), .Y(n_765) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g660 ( .A(n_620), .Y(n_660) );
AND3x1_ASAP7_75t_L g756 ( .A(n_620), .B(n_757), .C(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g743 ( .A(n_621), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g753 ( .A(n_621), .Y(n_753) );
INVxp67_ASAP7_75t_L g767 ( .A(n_623), .Y(n_767) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
OR2x2_ASAP7_75t_L g722 ( .A(n_626), .B(n_646), .Y(n_722) );
INVx2_ASAP7_75t_L g757 ( .A(n_626), .Y(n_757) );
INVx1_ASAP7_75t_L g675 ( .A(n_627), .Y(n_675) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_629), .A2(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_630), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g638 ( .A(n_631), .Y(n_638) );
OR2x2_ASAP7_75t_L g732 ( .A(n_631), .B(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g692 ( .A(n_634), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_634), .B(n_691), .Y(n_771) );
AND3x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_642), .C(n_647), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x2_ASAP7_75t_L g686 ( .A(n_638), .B(n_677), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_639), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_705) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OAI321xp33_ASAP7_75t_L g728 ( .A1(n_640), .A2(n_729), .A3(n_730), .B1(n_732), .B2(n_735), .C(n_737), .Y(n_728) );
AND2x2_ASAP7_75t_L g780 ( .A(n_640), .B(n_645), .Y(n_780) );
AND2x2_ASAP7_75t_L g678 ( .A(n_641), .B(n_644), .Y(n_678) );
INVx2_ASAP7_75t_L g687 ( .A(n_643), .Y(n_687) );
AND2x2_ASAP7_75t_L g696 ( .A(n_643), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g708 ( .A(n_646), .B(n_698), .Y(n_708) );
INVx2_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_656), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g744 ( .A(n_650), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_653), .B(n_660), .Y(n_670) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_662), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_660), .B(n_684), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_660), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g761 ( .A(n_660), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g729 ( .A(n_662), .Y(n_729) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_664), .B(n_726), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_688), .C(n_711), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_679), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B1(n_671), .B2(n_674), .C(n_676), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OR2x2_ASAP7_75t_L g719 ( .A(n_668), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI21xp33_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_685), .B(n_687), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g716 ( .A(n_684), .B(n_717), .Y(n_716) );
OAI21xp33_ASAP7_75t_SL g699 ( .A1(n_685), .A2(n_700), .B(n_705), .Y(n_699) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_693), .B(n_696), .C(n_699), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_690), .B(n_765), .Y(n_764) );
NAND2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_698), .B(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_701), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_718), .B1(n_721), .B2(n_723), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_720), .Y(n_783) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_763), .C(n_778), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_745), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_741), .B(n_743), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_751), .C(n_760), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
AOI32xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .A3(n_755), .B1(n_756), .B2(n_759), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g779 ( .A(n_754), .B(n_780), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_768), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI22x1_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B1(n_773), .B2(n_775), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g782 ( .A1(n_771), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx8_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx12f_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g793 ( .A(n_789), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx5_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x6_ASAP7_75t_SL g796 ( .A(n_797), .B(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx3_ASAP7_75t_L g808 ( .A(n_798), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_798), .B(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_801), .B(n_803), .Y(n_839) );
AND2x6_ASAP7_75t_SL g815 ( .A(n_802), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_809), .B(n_832), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B(n_824), .Y(n_809) );
OAI31xp33_ASAP7_75t_SL g824 ( .A1(n_810), .A2(n_819), .A3(n_825), .B(n_828), .Y(n_824) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_819), .Y(n_812) );
BUFx12f_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx4_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx5_ASAP7_75t_L g827 ( .A(n_815), .Y(n_827) );
INVx5_ASAP7_75t_L g831 ( .A(n_815), .Y(n_831) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_818), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
BUFx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx3_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx6_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx10_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
BUFx8_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_842), .Y(n_841) );
OR2x6_ASAP7_75t_L g842 ( .A(n_843), .B(n_850), .Y(n_842) );
OR2x6_ASAP7_75t_L g857 ( .A(n_843), .B(n_850), .Y(n_857) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NOR2x1p5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2x1p5_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx4_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx11_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
endmodule