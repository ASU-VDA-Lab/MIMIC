module fake_jpeg_7029_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_19),
.C(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_15),
.B1(n_20),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_12),
.B1(n_15),
.B2(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_12),
.C(n_18),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_28),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_76),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_9),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_75),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_49),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_87),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_59),
.C(n_42),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_89),
.C(n_90),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_91),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_65),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_41),
.C(n_47),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_48),
.B(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_66),
.B(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_79),
.A3(n_80),
.B1(n_87),
.B2(n_85),
.C1(n_9),
.C2(n_75),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_72),
.C(n_76),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_94),
.C(n_97),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_108),
.C(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_107),
.C(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_87),
.B1(n_71),
.B2(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_102),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_101),
.Y(n_107)
);

AOI211xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_50),
.B(n_69),
.C(n_71),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_93),
.C(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_108),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_104),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_78),
.B(n_84),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_115),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_117),
.B(n_118),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_122),
.Y(n_125)
);


endmodule