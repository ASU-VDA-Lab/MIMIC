module fake_jpeg_3734_n_120 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_9),
.Y(n_12)
);

BUFx3_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_14),
.B1(n_19),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_42),
.B1(n_16),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_30),
.B(n_13),
.C(n_26),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_34),
.B(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_48),
.B1(n_37),
.B2(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_63),
.B1(n_49),
.B2(n_38),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_46),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_36),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_65),
.C(n_50),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_33),
.C(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_42),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_60),
.C(n_59),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_77),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_43),
.B1(n_32),
.B2(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_40),
.B1(n_45),
.B2(n_58),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_12),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_76),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_47),
.C(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_45),
.B1(n_40),
.B2(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_35),
.B(n_45),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_21),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_86),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_68),
.B1(n_11),
.B2(n_54),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_35),
.C(n_30),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_54),
.C(n_22),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_87),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_99),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_82),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.Y(n_113)
);

AOI321xp33_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_94),
.A3(n_98),
.B1(n_101),
.B2(n_100),
.C(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_111),
.A3(n_109),
.B1(n_9),
.B2(n_21),
.C1(n_22),
.C2(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_116),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_21),
.A3(n_22),
.B1(n_4),
.B2(n_5),
.C1(n_1),
.C2(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_118),
.Y(n_120)
);


endmodule