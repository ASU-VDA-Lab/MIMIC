module real_jpeg_2120_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_4),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_33),
.B1(n_38),
.B2(n_86),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_86),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_77),
.B1(n_79),
.B2(n_86),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_33),
.B1(n_38),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_66),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_66),
.B1(n_77),
.B2(n_79),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_42),
.B1(n_61),
.B2(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_42),
.B1(n_77),
.B2(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_33),
.B1(n_38),
.B2(n_42),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_30),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_7),
.B(n_43),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_38),
.B(n_58),
.C(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_7),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_7),
.B(n_60),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_7),
.A2(n_33),
.B1(n_38),
.B2(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_7),
.B(n_74),
.C(n_77),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_7),
.B(n_106),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_95),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_8),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_8),
.A2(n_33),
.B1(n_38),
.B2(n_138),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_138),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_8),
.A2(n_77),
.B1(n_79),
.B2(n_138),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_9),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_33),
.B1(n_38),
.B2(n_116),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_116),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_9),
.A2(n_77),
.B1(n_79),
.B2(n_116),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_10),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_33),
.B1(n_38),
.B2(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_178),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_10),
.A2(n_77),
.B1(n_79),
.B2(n_178),
.Y(n_288)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_20),
.B(n_345),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_14),
.B(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_15),
.A2(n_26),
.B1(n_61),
.B2(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_26),
.B1(n_33),
.B2(n_38),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_15),
.A2(n_26),
.B1(n_77),
.B2(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_33),
.B1(n_38),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_16),
.A2(n_61),
.B1(n_62),
.B2(n_69),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_16),
.A2(n_27),
.B1(n_30),
.B2(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_16),
.A2(n_69),
.B1(n_77),
.B2(n_79),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_23),
.B(n_344),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_24),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_24),
.B(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_41),
.B2(n_43),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_25),
.A2(n_31),
.B1(n_43),
.B2(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g198 ( 
.A1(n_27),
.A2(n_36),
.A3(n_38),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_27),
.A2(n_87),
.B(n_228),
.C(n_237),
.Y(n_236)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_41),
.B(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_31),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_31),
.A2(n_43),
.B1(n_137),
.B2(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_32),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_85),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_32),
.B(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_32),
.A2(n_87),
.B1(n_88),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_32),
.A2(n_113),
.B(n_192),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_33),
.B(n_39),
.Y(n_200)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

OAI21x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_340),
.B(n_342),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_328),
.B(n_339),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_154),
.B(n_325),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_141),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_117),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_52),
.B(n_117),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_98),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_82),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_54),
.A2(n_55),
.B(n_70),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_54),
.B(n_82),
.C(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_70),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_56),
.A2(n_65),
.B1(n_67),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_56),
.A2(n_67),
.B1(n_92),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_56),
.A2(n_194),
.B(n_196),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_56),
.A2(n_196),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_57),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_57),
.A2(n_60),
.B1(n_195),
.B2(n_212),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_57),
.A2(n_60),
.B(n_332),
.Y(n_331)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_60),
.B(n_175),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_61),
.A2(n_64),
.B(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_62),
.B(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_67),
.A2(n_134),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_67),
.A2(n_174),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_76),
.B1(n_80),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_71),
.A2(n_76),
.B1(n_221),
.B2(n_255),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_71),
.A2(n_223),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_95),
.B1(n_111),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_72),
.A2(n_95),
.B1(n_132),
.B2(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_72),
.A2(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_72),
.B(n_224),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_76),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_76),
.A2(n_244),
.B(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_77),
.B(n_284),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_97),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_84),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g152 ( 
.A(n_84),
.B(n_90),
.C(n_94),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_84),
.B(n_145),
.C(n_152),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_136),
.B(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_94),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_94),
.B(n_146),
.C(n_150),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_95),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B(n_112),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_100),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_102),
.B1(n_112),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_101),
.A2(n_102),
.B1(n_109),
.B2(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_107),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_106),
.B1(n_129),
.B2(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_103),
.A2(n_228),
.B(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_104),
.A2(n_105),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_104),
.A2(n_105),
.B1(n_203),
.B2(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_104),
.B(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_104),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_104),
.A2(n_105),
.B1(n_259),
.B2(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_105),
.A2(n_218),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_105),
.B(n_232),
.Y(n_261)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_106),
.A2(n_231),
.B(n_288),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_124),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_135),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_135),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_140),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_141),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_153),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_142),
.B(n_153),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_147),
.Y(n_334)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_151),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_179),
.B(n_324),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_156),
.B(n_159),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.C(n_176),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_167),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_168),
.B(n_170),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_205),
.B(n_323),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_181),
.B(n_183),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_184),
.B(n_188),
.Y(n_308)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_190),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_197),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_191),
.B(n_193),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_197),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_198),
.A2(n_201),
.B1(n_202),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI31xp33_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_305),
.A3(n_315),
.B(n_320),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_249),
.B(n_304),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_233),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_208),
.B(n_233),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.C(n_225),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_209),
.B(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_214),
.C(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_219),
.B(n_225),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_229),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_245),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_234),
.B(n_246),
.C(n_248),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_235),
.B(n_240),
.C(n_241),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_299),
.B(n_303),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_268),
.B(n_298),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_262),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_258),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_280),
.B(n_297),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_291),
.B(n_296),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_286),
.B(n_290),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_319),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_338),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_338),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_333),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_335),
.C(n_337),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_341),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule