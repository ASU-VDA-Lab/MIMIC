module fake_jpeg_14864_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_33),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_51),
.CON(n_71),
.SN(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_48),
.B1(n_44),
.B2(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_1),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_40),
.C(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_42),
.B2(n_54),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_53),
.B1(n_47),
.B2(n_45),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_43),
.B1(n_51),
.B2(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_7),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_5),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

CKINVDCx11_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_96),
.B1(n_11),
.B2(n_13),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_9),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_20),
.Y(n_109)
);

AND2x4_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_83),
.B1(n_91),
.B2(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_80),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.C(n_103),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_101),
.C(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_97),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_120),
.B(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.C(n_99),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_107),
.A3(n_117),
.B1(n_114),
.B2(n_102),
.C(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_23),
.C(n_24),
.Y(n_132)
);

AOI321xp33_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_26),
.A3(n_27),
.B1(n_29),
.B2(n_31),
.C(n_32),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_39),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_34),
.Y(n_135)
);


endmodule