module fake_jpeg_18453_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_47)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_45),
.B1(n_27),
.B2(n_42),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_52),
.B1(n_61),
.B2(n_24),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_15),
.B1(n_19),
.B2(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_22),
.B(n_27),
.Y(n_56)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_45),
.C(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_44),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_43),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_34),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_98),
.Y(n_125)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_87),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_41),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_23),
.C(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_102),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_39),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_29),
.B(n_26),
.C(n_24),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_31),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_41),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_99),
.C(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_29),
.B1(n_26),
.B2(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_46),
.B1(n_18),
.B2(n_24),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_42),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_22),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_39),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_42),
.C(n_39),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_49),
.B(n_30),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_118),
.B1(n_121),
.B2(n_108),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_137),
.B1(n_68),
.B2(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_138),
.C(n_99),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_100),
.B(n_99),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_74),
.C(n_80),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_32),
.A3(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_141),
.Y(n_146)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_100),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_72),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_147),
.B1(n_155),
.B2(n_157),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_79),
.B1(n_76),
.B2(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_148),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_83),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_154),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_127),
.B1(n_132),
.B2(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_171),
.B(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_73),
.B1(n_71),
.B2(n_91),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_71),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_161),
.B(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_114),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_84),
.B1(n_96),
.B2(n_95),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_173),
.B1(n_175),
.B2(n_158),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_93),
.B(n_84),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_96),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_175),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_108),
.A2(n_86),
.B1(n_102),
.B2(n_85),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_31),
.B(n_25),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_86),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_144),
.C(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_157),
.C(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_199),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_R g181 ( 
.A(n_171),
.B(n_122),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_195),
.B(n_159),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_141),
.B1(n_142),
.B2(n_126),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_183),
.A2(n_201),
.B1(n_2),
.B2(n_4),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_192),
.B1(n_205),
.B2(n_0),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_122),
.B1(n_139),
.B2(n_142),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_139),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_119),
.B(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_126),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_150),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_172),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_131),
.B1(n_129),
.B2(n_23),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_152),
.A2(n_131),
.B1(n_66),
.B2(n_17),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_0),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_147),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_176),
.B1(n_191),
.B2(n_196),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_208),
.B(n_210),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_170),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_211),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_174),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_215),
.B1(n_184),
.B2(n_195),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_232),
.C(n_223),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_154),
.B(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_177),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_160),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_9),
.B1(n_8),
.B2(n_3),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_9),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_233),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_234),
.B1(n_205),
.B2(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_8),
.C(n_3),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_2),
.C(n_4),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_187),
.C(n_200),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_187),
.C(n_196),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_211),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_207),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_223),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_268),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_218),
.B1(n_224),
.B2(n_176),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_244),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_228),
.C(n_213),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_260),
.B(n_265),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_215),
.B(n_216),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_257),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_218),
.B(n_227),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_179),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_232),
.C(n_198),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_270),
.C(n_274),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_203),
.C(n_185),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_189),
.C(n_233),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_185),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_284),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_239),
.B1(n_255),
.B2(n_252),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_277),
.B1(n_283),
.B2(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_241),
.C(n_246),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_240),
.B1(n_241),
.B2(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_240),
.C(n_186),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_186),
.C(n_197),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_268),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_267),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_263),
.B(n_199),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_264),
.B1(n_259),
.B2(n_7),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_281),
.B1(n_286),
.B2(n_5),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_5),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_296),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_290),
.B1(n_281),
.B2(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_5),
.C(n_6),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_311),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_306),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_302),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_309),
.C(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_305),
.C(n_308),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_304),
.B(n_303),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_311),
.Y(n_320)
);


endmodule