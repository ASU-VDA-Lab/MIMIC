module fake_jpeg_27301_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_49),
.Y(n_96)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_36),
.B1(n_32),
.B2(n_19),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_40),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_36),
.B1(n_19),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_67),
.B1(n_61),
.B2(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_36),
.B1(n_42),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_90),
.B1(n_92),
.B2(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_44),
.B1(n_45),
.B2(n_27),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_45),
.B1(n_18),
.B2(n_35),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_105),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_52),
.B1(n_66),
.B2(n_58),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_91),
.B1(n_97),
.B2(n_93),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_107),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_25),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_48),
.B1(n_22),
.B2(n_26),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_80),
.B1(n_72),
.B2(n_77),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_120),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_85),
.C(n_43),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_40),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_40),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_86),
.Y(n_148)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_89),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_20),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_43),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_43),
.CI(n_48),
.CON(n_134),
.SN(n_134)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_152),
.Y(n_173)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_141),
.Y(n_165)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_54),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_100),
.B(n_102),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_156),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_43),
.CI(n_16),
.CON(n_152),
.SN(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_103),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_95),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_109),
.B(n_122),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_160),
.B(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_97),
.B1(n_108),
.B2(n_111),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_164),
.B1(n_183),
.B2(n_142),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_132),
.B(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_111),
.B1(n_108),
.B2(n_93),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_43),
.B(n_81),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_168),
.B(n_170),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_23),
.B(n_127),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_178),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_119),
.B(n_123),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_38),
.B(n_86),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_166),
.B(n_160),
.C(n_172),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_28),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_190),
.C(n_145),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_117),
.B1(n_112),
.B2(n_99),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_117),
.B1(n_112),
.B2(n_99),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_144),
.B1(n_131),
.B2(n_147),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_65),
.C(n_64),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_192),
.B(n_196),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_213),
.B(n_200),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_140),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_215),
.B1(n_162),
.B2(n_179),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_189),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_134),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_172),
.B(n_168),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_147),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_157),
.C(n_134),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_173),
.C(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_212),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_216),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_220),
.B1(n_176),
.B2(n_182),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_152),
.B1(n_142),
.B2(n_35),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_0),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_18),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_10),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_241),
.B1(n_202),
.B2(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_165),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_222),
.A2(n_224),
.B(n_246),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_163),
.B(n_165),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_211),
.B1(n_193),
.B2(n_202),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_233),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_190),
.B1(n_180),
.B2(n_173),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_236),
.B1(n_240),
.B2(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_30),
.B1(n_29),
.B2(n_4),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_242),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_8),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_214),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_192),
.B1(n_213),
.B2(n_207),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_195),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_191),
.A2(n_8),
.B(n_14),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_1),
.B(n_3),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_244),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

HAxp5_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_3),
.CON(n_246),
.SN(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_252),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_228),
.C(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_261),
.C(n_266),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_206),
.C(n_204),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.Y(n_272)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_204),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_245),
.B1(n_234),
.B2(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_9),
.C(n_11),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_224),
.A2(n_12),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_247),
.B(n_244),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_12),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_269),
.B(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_227),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_279),
.B(n_284),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_244),
.B(n_225),
.Y(n_279)
);

XOR2x1_ASAP7_75t_SL g281 ( 
.A(n_255),
.B(n_222),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_285),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_229),
.B(n_243),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_279),
.Y(n_306)
);

BUFx12_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_253),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_287),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_249),
.C(n_248),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

BUFx12_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_301),
.C(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_265),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_262),
.C(n_252),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_277),
.B1(n_300),
.B2(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_289),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_295),
.C(n_280),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_309),
.Y(n_316)
);

OAI22x1_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_259),
.B1(n_283),
.B2(n_246),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_290),
.B(n_247),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_312),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_283),
.C(n_282),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_260),
.B1(n_243),
.B2(n_263),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_289),
.Y(n_320)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_320),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_292),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_295),
.C(n_291),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_247),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_316),
.A2(n_314),
.B(n_307),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_326),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_311),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_315),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_325),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.A3(n_334),
.B1(n_325),
.B2(n_317),
.C1(n_323),
.C2(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_329),
.B(n_267),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_280),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_268),
.B(n_257),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_15),
.Y(n_341)
);


endmodule