module fake_jpeg_18083_n_274 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_14),
.B1(n_11),
.B2(n_19),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_14),
.B2(n_32),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_52),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_32),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_39),
.B1(n_42),
.B2(n_14),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_25),
.B(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_39),
.B1(n_42),
.B2(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_42),
.B1(n_35),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_36),
.B1(n_40),
.B2(n_29),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_53),
.B1(n_54),
.B2(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_49),
.B1(n_38),
.B2(n_58),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_94),
.B(n_79),
.Y(n_102)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_59),
.B1(n_46),
.B2(n_48),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_90),
.B1(n_73),
.B2(n_67),
.Y(n_118)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_87),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_38),
.B1(n_40),
.B2(n_14),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_93),
.B1(n_79),
.B2(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_43),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_43),
.CI(n_44),
.CON(n_107),
.SN(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_11),
.B1(n_19),
.B2(n_33),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_72),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_17),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_73),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_23),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_65),
.Y(n_101)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_17),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_107),
.B(n_23),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_104),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_105),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_80),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_111),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_78),
.A3(n_67),
.B1(n_70),
.B2(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_113),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_22),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_78),
.C(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_91),
.C(n_83),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_25),
.B1(n_28),
.B2(n_12),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_57),
.B1(n_69),
.B2(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_71),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_126),
.C(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_91),
.C(n_83),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_85),
.B(n_10),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_20),
.B1(n_7),
.B2(n_2),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_141),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_133),
.B1(n_139),
.B2(n_149),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_28),
.B1(n_12),
.B2(n_57),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_7),
.B1(n_10),
.B2(n_2),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_56),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_144),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_12),
.B1(n_23),
.B2(n_18),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_16),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_18),
.B(n_16),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_30),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_30),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_30),
.C(n_21),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_104),
.C(n_99),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_12),
.B1(n_18),
.B2(n_1),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_151),
.B(n_153),
.Y(n_190)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_170),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_131),
.C(n_138),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_119),
.B1(n_107),
.B2(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_107),
.B1(n_105),
.B2(n_21),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_165),
.B1(n_169),
.B2(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_172),
.B(n_20),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_21),
.B1(n_15),
.B2(n_2),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_169),
.B(n_166),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_128),
.B1(n_129),
.B2(n_148),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_195),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_131),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_164),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_9),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_134),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_144),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_5),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_15),
.C(n_20),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_152),
.C(n_156),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_15),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_9),
.C(n_3),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_208),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_168),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_207),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_154),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_156),
.B1(n_154),
.B2(n_171),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_20),
.C(n_1),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_215),
.C(n_193),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_5),
.B(n_8),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_5),
.B(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_198),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_187),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_179),
.B1(n_183),
.B2(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_182),
.C(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_237),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_199),
.B(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_205),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_227),
.C(n_209),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.C(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_208),
.B1(n_201),
.B2(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_225),
.C(n_6),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_249),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_3),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_3),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_6),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_234),
.B(n_231),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_256),
.B(n_8),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_257),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_232),
.B(n_4),
.Y(n_256)
);

NOR3x1_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_4),
.C(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_0),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_6),
.C(n_8),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_257),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_9),
.B(n_0),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_0),
.C(n_1),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_261),
.B(n_260),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_270),
.B(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_0),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);


endmodule