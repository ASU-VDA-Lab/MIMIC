module fake_jpeg_2505_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_1),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_63),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_75),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_55),
.B(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_52),
.B(n_48),
.C(n_59),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_60),
.B1(n_47),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_51),
.B1(n_53),
.B2(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_59),
.B1(n_67),
.B2(n_48),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_43),
.B1(n_53),
.B2(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_49),
.B1(n_67),
.B2(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_1),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_6),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_28),
.C(n_40),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_27),
.B(n_39),
.C(n_12),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

OAI221xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.C(n_15),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_26),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_29),
.C(n_38),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_23),
.C(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_16),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_122),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_118),
.B(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_124),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_120),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_137),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_136),
.A3(n_135),
.B1(n_132),
.B2(n_139),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_155),
.C(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_157),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_146),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_145),
.B(n_18),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_17),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_20),
.B(n_30),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_32),
.Y(n_164)
);


endmodule