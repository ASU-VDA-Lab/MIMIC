module fake_netlist_6_3660_n_87 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_87);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_87;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_0),
.B1(n_8),
.B2(n_3),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_12),
.B(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_8),
.A2(n_4),
.B1(n_9),
.B2(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AND2x6_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_1),
.B(n_27),
.C(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_1),
.B1(n_34),
.B2(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

OAI21x1_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_22),
.B(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_31),
.B(n_26),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_25),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_39),
.B(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_22),
.B1(n_30),
.B2(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OR2x6_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_44),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_53),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_52),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

OAI211xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_47),
.B(n_24),
.C(n_23),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_20),
.A3(n_23),
.B1(n_59),
.B2(n_54),
.C(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR4xp25_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_20),
.C(n_55),
.D(n_59),
.Y(n_73)
);

AOI211xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_66),
.B(n_28),
.C(n_62),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_51),
.B1(n_62),
.B2(n_60),
.C(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_51),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_51),
.B1(n_22),
.B2(n_60),
.C(n_49),
.Y(n_77)
);

NAND3x1_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_60),
.C(n_30),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_51),
.C(n_57),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_48),
.Y(n_80)
);

NAND4xp25_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_48),
.C(n_30),
.D(n_67),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_77),
.B1(n_67),
.B2(n_79),
.C(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

AOI221x1_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_81),
.B1(n_30),
.B2(n_78),
.C(n_48),
.Y(n_85)
);

OAI21x1_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_30),
.B(n_84),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_30),
.B(n_85),
.Y(n_87)
);


endmodule