module fake_jpeg_8944_n_278 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_52),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_14),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_29),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_37),
.B(n_34),
.C(n_31),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_72),
.B1(n_48),
.B2(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_33),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_74),
.B1(n_53),
.B2(n_46),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_37),
.B(n_34),
.C(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_29),
.B1(n_38),
.B2(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_72),
.B1(n_61),
.B2(n_83),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_69),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_56),
.B1(n_71),
.B2(n_74),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_89),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_90),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_87),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_26),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_95),
.C(n_62),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_22),
.B1(n_63),
.B2(n_16),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_22),
.B1(n_56),
.B2(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_32),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_107),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_115),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_57),
.CI(n_62),
.CON(n_100),
.SN(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_82),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_113),
.C(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_106),
.B1(n_117),
.B2(n_40),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_62),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_77),
.B(n_82),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_69),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_68),
.B1(n_18),
.B2(n_25),
.C(n_20),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_68),
.C(n_70),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_76),
.C(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_28),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_94),
.B1(n_93),
.B2(n_71),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_40),
.B1(n_47),
.B2(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_123),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_129),
.C(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_131),
.B(n_137),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_25),
.B(n_18),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_90),
.B(n_13),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_118),
.B(n_107),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_70),
.C(n_49),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_126),
.C(n_113),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_112),
.B1(n_100),
.B2(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_137),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_125),
.B(n_109),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_148),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_151),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

XNOR2x2_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_114),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_156),
.Y(n_179)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_102),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_100),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_136),
.B1(n_139),
.B2(n_124),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_139),
.B1(n_109),
.B2(n_140),
.Y(n_170)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_174),
.B1(n_164),
.B2(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_108),
.B1(n_105),
.B2(n_131),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_186),
.C(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_178),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_104),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_183),
.B(n_13),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_24),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_171),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_141),
.B1(n_149),
.B2(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_203),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_162),
.B1(n_144),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_205),
.B1(n_167),
.B2(n_173),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_84),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_156),
.B1(n_160),
.B2(n_110),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_179),
.B1(n_168),
.B2(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_7),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_17),
.B(n_20),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_66),
.B1(n_16),
.B2(n_23),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_175),
.C(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_210),
.C(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_185),
.C(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_84),
.C(n_75),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_65),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_9),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_17),
.B(n_10),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_205),
.B1(n_204),
.B2(n_23),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_27),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_10),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_44),
.C(n_41),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_27),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_27),
.CI(n_21),
.CON(n_229),
.SN(n_229)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_9),
.B(n_12),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_44),
.B1(n_41),
.B2(n_24),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_32),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_24),
.B1(n_21),
.B2(n_6),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_6),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_207),
.B1(n_213),
.B2(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_245),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_221),
.B1(n_217),
.B2(n_24),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_217),
.B(n_6),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_247),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_32),
.C(n_21),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_0),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_5),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_5),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_233),
.C(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_229),
.C(n_32),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_242),
.B(n_8),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_229),
.B(n_8),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_11),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_246),
.B(n_238),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_265),
.A3(n_11),
.B1(n_12),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_247),
.B(n_249),
.C(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_258),
.B(n_250),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_250),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_261),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_271),
.B(n_270),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_272),
.B(n_2),
.C(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_1),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_1),
.C(n_2),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_2),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_4),
.Y(n_278)
);


endmodule