module fake_jpeg_17387_n_49 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_49);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_37;
wire n_29;
wire n_43;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_10),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B(n_34),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_15),
.A2(n_0),
.B1(n_30),
.B2(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_26),
.C(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_30),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_25),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_36),
.B(n_32),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.C(n_18),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_16),
.B(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_45),
.B1(n_22),
.B2(n_19),
.Y(n_48)
);

INVxp33_ASAP7_75t_SL g49 ( 
.A(n_48),
.Y(n_49)
);


endmodule