module fake_jpeg_19678_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_23),
.B1(n_1),
.B2(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_18),
.B1(n_23),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_39),
.B1(n_26),
.B2(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_22),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_28),
.C(n_22),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_29),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_49),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_22),
.B1(n_16),
.B2(n_17),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_0),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_1),
.B1(n_4),
.B2(n_11),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_6),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_9),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_49),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_50),
.B1(n_64),
.B2(n_60),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_50),
.B(n_54),
.Y(n_78)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_46),
.B(n_55),
.C(n_52),
.D(n_44),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_65),
.Y(n_84)
);

AOI211xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_48),
.B(n_59),
.C(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_71),
.B1(n_69),
.B2(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_72),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_85),
.C(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_65),
.C(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_90),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_87),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_81),
.B(n_79),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_69),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_37),
.C(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_86),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_87),
.C(n_83),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_83),
.B(n_94),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_98),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_10),
.Y(n_103)
);


endmodule