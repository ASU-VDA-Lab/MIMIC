module real_jpeg_22588_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_139;
wire n_33;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_8),
.B1(n_45),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_7),
.B1(n_48),
.B2(n_54),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_6),
.B1(n_37),
.B2(n_48),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_6),
.B(n_72),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_1),
.A2(n_5),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_5),
.B1(n_24),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_6),
.B1(n_37),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_37),
.B(n_45),
.C(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_9),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_5),
.A2(n_6),
.B1(n_24),
.B2(n_37),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_6),
.B(n_9),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_10),
.B1(n_35),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_6),
.B(n_53),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_7),
.B(n_48),
.C(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_6),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_10),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_10),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_32),
.B(n_37),
.C(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_87),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_86),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_78),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_67),
.B2(n_77),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_29),
.B2(n_38),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_21),
.A2(n_23),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_24),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_26),
.B(n_37),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_29),
.A2(n_38),
.B1(n_61),
.B2(n_82),
.Y(n_81)
);

AOI211xp5_ASAP7_75t_SL g84 ( 
.A1(n_29),
.A2(n_58),
.B(n_76),
.C(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_29),
.A2(n_38),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_29),
.A2(n_38),
.B1(n_96),
.B2(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_73),
.C(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_29),
.A2(n_38),
.B1(n_51),
.B2(n_59),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_29),
.A2(n_38),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_29),
.B(n_130),
.C(n_139),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_31),
.B(n_37),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_35),
.A2(n_37),
.B(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_38),
.B(n_96),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_38),
.A2(n_59),
.B(n_124),
.C(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_60),
.B2(n_64),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_41),
.B1(n_68),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_59),
.B(n_68),
.C(n_75),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_42),
.A2(n_58),
.B1(n_122),
.B2(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_51),
.A2(n_59),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_73),
.C(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_74),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_102),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_73),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_102),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_73),
.A2(n_102),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

NAND2x1_ASAP7_75t_SL g140 ( 
.A(n_73),
.B(n_119),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_81),
.Y(n_158)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_159),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_154),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_142),
.B(n_153),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_126),
.B(n_141),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_115),
.B(n_125),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_104),
.B(n_114),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_144),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);


endmodule