module fake_ariane_974_n_2231 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2231);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2231;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_967;
wire n_274;
wire n_437;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g238 ( 
.A(n_24),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_109),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_29),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_190),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_29),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_150),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_25),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_100),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_138),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_145),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_152),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_68),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_62),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_47),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_162),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_128),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_112),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_61),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_158),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_147),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_55),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_125),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_97),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_199),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_68),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_139),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_228),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_61),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_182),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_41),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_122),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_79),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_168),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_23),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_70),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_204),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_133),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_73),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_75),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_114),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_95),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_186),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_16),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_45),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_16),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_79),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_132),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_135),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_20),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_92),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_77),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_197),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_72),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_35),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_126),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_90),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_175),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_165),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_116),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_73),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_88),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_36),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_196),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_81),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_55),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_1),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_185),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_69),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_57),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_172),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_96),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_176),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_32),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_149),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_167),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_177),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_82),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_194),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_4),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_36),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_66),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_39),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_27),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_235),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_32),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_66),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_217),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_198),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_17),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_123),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_208),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_30),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_205),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_206),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_74),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_118),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_161),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_74),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_39),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_45),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_153),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_160),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_127),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_101),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_108),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_18),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_200),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_230),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_58),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_44),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_12),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_131),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_98),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_203),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_195),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_54),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_21),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_102),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_51),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_232),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_85),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_40),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_91),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_28),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_11),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_0),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_12),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_10),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_13),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_78),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_43),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_104),
.Y(n_412)
);

BUFx8_ASAP7_75t_SL g413 ( 
.A(n_183),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_226),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_44),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_3),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_136),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_120),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_51),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_184),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_22),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_163),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_60),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_134),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_221),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_47),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_144),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_87),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_170),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_99),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_25),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_94),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_42),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_58),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_236),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_223),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_137),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_72),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_67),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_124),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_84),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_148),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_0),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_65),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_59),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_201),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_130),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_42),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_115),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_225),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_54),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_141),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_78),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_20),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_49),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_2),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_15),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_34),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_19),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_18),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_50),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_10),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_37),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_121),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_106),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_159),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_297),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_322),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_322),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_324),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_359),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_250),
.B(n_80),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_341),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_239),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_318),
.B(n_4),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_252),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_326),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_404),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_329),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_372),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_241),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_258),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_287),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_238),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_302),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_337),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_241),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_302),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_241),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_246),
.B(n_5),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_360),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_292),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_360),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_357),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_239),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_337),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_317),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_467),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_317),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_249),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_242),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_378),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_255),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_317),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_373),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_263),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_254),
.B(n_6),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_266),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_334),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_323),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_275),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_279),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_323),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_425),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_447),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_281),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_256),
.B(n_6),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_343),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_323),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_344),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_367),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_298),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_423),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_313),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_240),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_240),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_325),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_358),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_361),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_363),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_377),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_379),
.B(n_7),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_243),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_390),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_399),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_379),
.B(n_8),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_451),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_406),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_243),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_272),
.B(n_9),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_411),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_334),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_433),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_438),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_244),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_453),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_244),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_456),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_247),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_247),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_454),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_464),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_458),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_245),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_337),
.B(n_9),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_257),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_459),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_245),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_301),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_L g579 ( 
.A(n_407),
.B(n_13),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_248),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_248),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_251),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_251),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_257),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_413),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_273),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_285),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_249),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_259),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_276),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_259),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_265),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_261),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_267),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_291),
.B(n_14),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_586),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_522),
.B(n_285),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_586),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_531),
.B(n_267),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_533),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_587),
.B(n_261),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_534),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_568),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_R g605 ( 
.A(n_585),
.B(n_283),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_569),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_489),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_569),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_575),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_592),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_491),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_536),
.B(n_268),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_584),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_584),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_501),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_488),
.B(n_496),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_538),
.B(n_310),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_552),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_538),
.B(n_539),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_590),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_497),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_594),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_505),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_500),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_503),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_511),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_503),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_511),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_518),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_504),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_488),
.B(n_262),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_527),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_507),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_509),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_528),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_468),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_506),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_509),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_565),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_574),
.B(n_260),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_506),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_496),
.B(n_262),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_539),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_565),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_556),
.Y(n_652)
);

NAND2x1_ASAP7_75t_L g653 ( 
.A(n_574),
.B(n_310),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_567),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_339),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_356),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_471),
.B(n_375),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_494),
.B(n_268),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_560),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_546),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_570),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_546),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_493),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_469),
.B(n_294),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_468),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_555),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_555),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_571),
.Y(n_673)
);

OA21x2_ASAP7_75t_L g674 ( 
.A1(n_557),
.A2(n_319),
.B(n_314),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_563),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_514),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_513),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_502),
.B(n_269),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_480),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_498),
.B(n_510),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_495),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_519),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_480),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_521),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_588),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_R g687 ( 
.A(n_485),
.B(n_269),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_561),
.B(n_271),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_563),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_524),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_498),
.B(n_321),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_525),
.Y(n_692)
);

INVx4_ASAP7_75t_SL g693 ( 
.A(n_647),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_663),
.B(n_667),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_477),
.B1(n_573),
.B2(n_566),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_647),
.A2(n_595),
.B1(n_545),
.B2(n_576),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_663),
.B(n_566),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_667),
.B(n_573),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_670),
.B(n_260),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_621),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_670),
.B(n_510),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_598),
.B(n_278),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_691),
.B(n_577),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_647),
.A2(n_572),
.B1(n_564),
.B2(n_529),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_597),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_661),
.B(n_512),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_642),
.B(n_476),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_658),
.B(n_508),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_650),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_630),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_681),
.B(n_577),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_630),
.Y(n_714)
);

INVx6_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_679),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_601),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_648),
.A2(n_580),
.B1(n_582),
.B2(n_581),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_660),
.B(n_580),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_661),
.B(n_512),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_660),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_662),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_598),
.B(n_486),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_661),
.B(n_517),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_679),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_597),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_597),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_647),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_647),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_647),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_688),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_597),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_655),
.B(n_581),
.Y(n_733)
);

XNOR2xp5_ASAP7_75t_L g734 ( 
.A(n_603),
.B(n_478),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_643),
.B(n_473),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_683),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_683),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_598),
.B(n_656),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_666),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_666),
.Y(n_741)
);

AND2x2_ASAP7_75t_SL g742 ( 
.A(n_674),
.B(n_278),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_666),
.Y(n_743)
);

INVx6_ASAP7_75t_L g744 ( 
.A(n_598),
.Y(n_744)
);

BUFx4f_ASAP7_75t_L g745 ( 
.A(n_655),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_685),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_627),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_665),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_596),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_684),
.B(n_485),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_630),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_627),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_677),
.B(n_487),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_685),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_686),
.B(n_487),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_656),
.B(n_362),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_630),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_656),
.B(n_647),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_632),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_632),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_685),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_632),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_656),
.B(n_622),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_596),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_692),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_655),
.B(n_582),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_517),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_636),
.B(n_583),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_632),
.B(n_523),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_692),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_671),
.B(n_583),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_659),
.B(n_362),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_606),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_687),
.A2(n_515),
.B1(n_277),
.B2(n_280),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_692),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_602),
.A2(n_589),
.B1(n_593),
.B2(n_591),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_669),
.B(n_589),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_645),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_676),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_672),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_690),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_659),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_627),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_690),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_523),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_652),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_645),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_620),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_627),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_653),
.B(n_526),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_675),
.B(n_591),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_596),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_627),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_689),
.B(n_593),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_678),
.B(n_430),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_652),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_604),
.Y(n_800)
);

BUFx6f_ASAP7_75t_SL g801 ( 
.A(n_642),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_SL g802 ( 
.A(n_649),
.B(n_277),
.C(n_271),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_678),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_604),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_627),
.Y(n_805)
);

AND3x2_ASAP7_75t_L g806 ( 
.A(n_669),
.B(n_578),
.C(n_537),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_607),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_680),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_628),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_607),
.B(n_430),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_596),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_680),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_618),
.B(n_526),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_664),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_599),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_668),
.B(n_532),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_628),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_599),
.Y(n_819)
);

BUFx4f_ASAP7_75t_L g820 ( 
.A(n_674),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_628),
.B(n_532),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_628),
.B(n_330),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_653),
.B(n_470),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_SL g824 ( 
.A(n_605),
.B(n_475),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_674),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_609),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_610),
.B(n_441),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_674),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_610),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_616),
.B(n_472),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_628),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_616),
.B(n_264),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_628),
.B(n_332),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_673),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_599),
.B(n_474),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_615),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_623),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_599),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_481),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_615),
.B(n_333),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_624),
.B(n_482),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_629),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_608),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_624),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_629),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_631),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_629),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_613),
.B(n_280),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_625),
.B(n_483),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_625),
.B(n_484),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_617),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_799),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_694),
.B(n_631),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_808),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_728),
.B(n_264),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_728),
.B(n_274),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_713),
.A2(n_579),
.B1(n_431),
.B2(n_434),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_779),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_749),
.B(n_764),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_808),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_749),
.B(n_633),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_782),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_R g863 ( 
.A(n_773),
.B(n_626),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_813),
.B(n_612),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_772),
.A2(n_376),
.B1(n_401),
.B2(n_356),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_764),
.B(n_811),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_713),
.B(n_633),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_729),
.B(n_274),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_729),
.B(n_353),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_697),
.A2(n_638),
.B(n_644),
.C(n_635),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_847),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_785),
.A2(n_431),
.B1(n_434),
.B2(n_421),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_702),
.B(n_439),
.C(n_421),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_811),
.B(n_635),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_772),
.A2(n_376),
.B1(n_401),
.B2(n_353),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_731),
.B(n_638),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_784),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_819),
.B(n_705),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_SL g879 ( 
.A1(n_709),
.A2(n_634),
.B1(n_641),
.B2(n_637),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_759),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_819),
.B(n_644),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_787),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_835),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_717),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_705),
.B(n_646),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_750),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_843),
.B(n_646),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_736),
.B(n_614),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_780),
.B(n_651),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_731),
.A2(n_657),
.B(n_651),
.C(n_640),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_806),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_697),
.B(n_657),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_803),
.B(n_682),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_719),
.B(n_639),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_800),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_804),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_759),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_769),
.A2(n_640),
.B(n_639),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_742),
.A2(n_478),
.B1(n_640),
.B2(n_639),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_730),
.B(n_422),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_717),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_721),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_806),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_726),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_698),
.A2(n_540),
.B(n_541),
.C(n_535),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_719),
.B(n_654),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_739),
.B(n_654),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_807),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_772),
.A2(n_422),
.B1(n_424),
.B2(n_428),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_772),
.B(n_654),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_742),
.A2(n_772),
.B1(n_798),
.B2(n_820),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_812),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_775),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_798),
.A2(n_543),
.B1(n_542),
.B2(n_562),
.Y(n_914)
);

OAI22xp33_ASAP7_75t_L g915 ( 
.A1(n_774),
.A2(n_439),
.B1(n_443),
.B2(n_444),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_798),
.B(n_424),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_798),
.B(n_763),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_698),
.B(n_284),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_715),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_851),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_817),
.B(n_288),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_715),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_730),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_798),
.B(n_763),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_745),
.B(n_428),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_763),
.B(n_429),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_826),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_763),
.B(n_429),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_775),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_763),
.B(n_432),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_696),
.B(n_432),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_745),
.B(n_435),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_696),
.B(n_435),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_721),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_715),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_795),
.B(n_436),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_817),
.B(n_290),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_829),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_718),
.B(n_444),
.C(n_443),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_837),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_795),
.B(n_436),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_816),
.B(n_440),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_816),
.B(n_440),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_726),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_820),
.B(n_449),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_699),
.B(n_449),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_699),
.B(n_767),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_695),
.B(n_490),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_699),
.B(n_450),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_704),
.B(n_293),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_704),
.A2(n_550),
.B(n_559),
.C(n_558),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_753),
.B(n_614),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_699),
.B(n_450),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_699),
.B(n_452),
.Y(n_954)
);

OAI22xp33_ASAP7_75t_L g955 ( 
.A1(n_774),
.A2(n_445),
.B1(n_448),
.B2(n_455),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_755),
.B(n_492),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_712),
.B(n_295),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_771),
.B(n_448),
.C(n_445),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_768),
.B(n_452),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_SL g960 ( 
.A(n_771),
.B(n_455),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_768),
.B(n_466),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_844),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_733),
.A2(n_466),
.B1(n_366),
.B2(n_369),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_825),
.B(n_338),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_846),
.B(n_296),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_825),
.A2(n_547),
.B(n_554),
.C(n_553),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_740),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_708),
.B(n_544),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_828),
.B(n_342),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_791),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_744),
.A2(n_457),
.B1(n_460),
.B2(n_462),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_708),
.B(n_548),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_850),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_741),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_712),
.B(n_300),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_707),
.B(n_304),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_733),
.B(n_306),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_828),
.A2(n_549),
.B(n_457),
.C(n_460),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_794),
.B(n_345),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_743),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_788),
.A2(n_352),
.B(n_348),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_815),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_849),
.B(n_600),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_746),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_726),
.Y(n_985)
);

NAND2x1_ASAP7_75t_L g986 ( 
.A(n_838),
.B(n_253),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_708),
.B(n_600),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_766),
.B(n_307),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_720),
.B(n_311),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_754),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_724),
.B(n_312),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_761),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_744),
.B(n_327),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_726),
.B(n_365),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_710),
.B(n_462),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_744),
.B(n_328),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_747),
.B(n_371),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_710),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_747),
.B(n_380),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_722),
.B(n_463),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_716),
.B(n_335),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_747),
.B(n_382),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_725),
.B(n_340),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_747),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_842),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_SL g1006 ( 
.A(n_722),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_834),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_752),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_693),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_737),
.B(n_349),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_734),
.B(n_463),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_766),
.B(n_355),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_738),
.B(n_364),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_794),
.B(n_370),
.C(n_374),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_752),
.B(n_786),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_752),
.B(n_386),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_830),
.B(n_389),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_884),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_867),
.B(n_700),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_854),
.B(n_700),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_860),
.B(n_748),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_911),
.A2(n_777),
.B1(n_797),
.B2(n_830),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_913),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_982),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_858),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_1009),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_923),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_867),
.B(n_723),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_859),
.A2(n_866),
.B(n_894),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_863),
.Y(n_1030)
);

CKINVDCx10_ASAP7_75t_R g1031 ( 
.A(n_1006),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_915),
.A2(n_955),
.B(n_872),
.C(n_978),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_876),
.B(n_723),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_862),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_853),
.A2(n_838),
.B1(n_758),
.B2(n_790),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_973),
.B(n_952),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_876),
.B(n_839),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_957),
.A2(n_824),
.B1(n_802),
.B2(n_821),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_970),
.B(n_793),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_892),
.B(n_839),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_892),
.B(n_703),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_918),
.A2(n_824),
.B(n_802),
.C(n_821),
.Y(n_1042)
);

CKINVDCx8_ASAP7_75t_R g1043 ( 
.A(n_920),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_906),
.A2(n_790),
.B(n_832),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_902),
.A2(n_934),
.B(n_874),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_888),
.B(n_748),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_919),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_945),
.A2(n_814),
.B(n_735),
.C(n_776),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_861),
.A2(n_735),
.B(n_706),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_959),
.B(n_703),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_881),
.A2(n_706),
.B(n_701),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_983),
.A2(n_801),
.B1(n_756),
.B2(n_703),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_945),
.A2(n_727),
.B(n_701),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_889),
.B(n_783),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_947),
.A2(n_732),
.B(n_727),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_890),
.A2(n_966),
.B(n_964),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_961),
.B(n_703),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_911),
.A2(n_814),
.B1(n_765),
.B2(n_770),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1015),
.A2(n_732),
.B(n_796),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_964),
.A2(n_833),
.B(n_822),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1015),
.A2(n_831),
.B(n_818),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_863),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_864),
.B(n_783),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_855),
.A2(n_845),
.B(n_823),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_915),
.A2(n_841),
.B(n_711),
.C(n_781),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_855),
.A2(n_845),
.B(n_751),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_956),
.B(n_752),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_878),
.A2(n_848),
.B1(n_714),
.B2(n_757),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1017),
.B(n_703),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_883),
.B(n_756),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_886),
.B(n_801),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_1009),
.B(n_809),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_929),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_909),
.B(n_786),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_1007),
.Y(n_1075)
);

AO221x2_ASAP7_75t_L g1076 ( 
.A1(n_955),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.C(n_21),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1011),
.B(n_836),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_890),
.A2(n_762),
.B(n_760),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_966),
.A2(n_778),
.B(n_833),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_856),
.A2(n_786),
.B(n_805),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_995),
.B(n_840),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_979),
.B(n_786),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_856),
.A2(n_792),
.B(n_805),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_914),
.A2(n_416),
.B1(n_397),
.B2(n_408),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_950),
.B(n_918),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_998),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_868),
.A2(n_792),
.B(n_805),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_957),
.A2(n_756),
.B1(n_827),
.B2(n_810),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_868),
.A2(n_792),
.B(n_805),
.Y(n_1089)
);

AO21x1_ASAP7_75t_L g1090 ( 
.A1(n_969),
.A2(n_822),
.B(n_840),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_901),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_877),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_898),
.A2(n_789),
.B(n_810),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_950),
.A2(n_392),
.B(n_393),
.C(n_395),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_969),
.A2(n_446),
.B(n_418),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_921),
.B(n_937),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_869),
.A2(n_792),
.B(n_809),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_869),
.A2(n_809),
.B(n_286),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_887),
.B(n_693),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_923),
.B(n_693),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_921),
.B(n_756),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_919),
.B(n_809),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_914),
.A2(n_405),
.B1(n_402),
.B2(n_400),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_900),
.A2(n_368),
.B(n_289),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_900),
.A2(n_442),
.B(n_420),
.C(n_398),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_922),
.B(n_299),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_895),
.A2(n_465),
.B1(n_441),
.B2(n_387),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_975),
.B(n_977),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_907),
.A2(n_351),
.B(n_303),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_937),
.B(n_756),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_975),
.A2(n_354),
.B(n_305),
.C(n_308),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_968),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_977),
.B(n_810),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_968),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_968),
.B(n_810),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_978),
.A2(n_870),
.B(n_967),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_L g1117 ( 
.A(n_939),
.B(n_309),
.C(n_315),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1000),
.B(n_810),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_988),
.B(n_383),
.C(n_316),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_972),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_910),
.A2(n_827),
.B(n_331),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_R g1122 ( 
.A(n_998),
.B(n_320),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_880),
.A2(n_384),
.B(n_336),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_882),
.B(n_827),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_981),
.A2(n_827),
.B(n_26),
.C(n_27),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_896),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_988),
.A2(n_388),
.B(n_346),
.C(n_347),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_917),
.A2(n_827),
.B(n_331),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_872),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_922),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_897),
.A2(n_394),
.B(n_350),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_972),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_908),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_857),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_912),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_944),
.A2(n_403),
.B(n_381),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1004),
.A2(n_412),
.B(n_414),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_927),
.B(n_417),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_891),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1008),
.A2(n_437),
.B(n_427),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_972),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1012),
.B(n_37),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1012),
.A2(n_437),
.B(n_427),
.C(n_282),
.Y(n_1143)
);

AO221x2_ASAP7_75t_L g1144 ( 
.A1(n_971),
.A2(n_958),
.B1(n_1014),
.B2(n_873),
.C(n_933),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_974),
.A2(n_331),
.B(n_40),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_931),
.A2(n_38),
.B(n_41),
.C(n_43),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_948),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_871),
.A2(n_991),
.B(n_989),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_935),
.B(n_331),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_924),
.A2(n_331),
.B(n_437),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_976),
.A2(n_437),
.B(n_427),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_938),
.B(n_940),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_903),
.B(n_38),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_962),
.A2(n_427),
.B1(n_282),
.B2(n_270),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_899),
.B(n_46),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_936),
.A2(n_282),
.B(n_270),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_986),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1005),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_925),
.B(n_932),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_965),
.A2(n_941),
.B(n_943),
.C(n_942),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_926),
.A2(n_282),
.B(n_270),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_935),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_928),
.A2(n_282),
.B(n_270),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_963),
.A2(n_331),
.B1(n_270),
.B2(n_253),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_994),
.A2(n_331),
.B(n_253),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_904),
.B(n_253),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_930),
.A2(n_253),
.B(n_331),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_980),
.A2(n_990),
.B(n_992),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_899),
.A2(n_885),
.B1(n_852),
.B2(n_984),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_925),
.B(n_48),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_932),
.B(n_50),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_960),
.B(n_52),
.C(n_53),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_879),
.B(n_52),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_951),
.A2(n_53),
.B(n_56),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_987),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1001),
.A2(n_56),
.B(n_59),
.C(n_62),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_904),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_993),
.B(n_63),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_904),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1003),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_905),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_875),
.B(n_64),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_904),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_996),
.A2(n_67),
.B(n_69),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1010),
.A2(n_151),
.B(n_231),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_987),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1013),
.B(n_70),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_985),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_865),
.A2(n_71),
.B(n_75),
.C(n_76),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_985),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1016),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_994),
.A2(n_83),
.B(n_86),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_893),
.B(n_237),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_916),
.B(n_93),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_985),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_985),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_997),
.A2(n_117),
.B(n_119),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_946),
.A2(n_129),
.B(n_140),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_949),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_953),
.A2(n_142),
.B(n_143),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_997),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_954),
.A2(n_1016),
.B1(n_1002),
.B2(n_999),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1108),
.A2(n_1002),
.B(n_999),
.C(n_987),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1090),
.A2(n_146),
.A3(n_155),
.B(n_157),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1028),
.B(n_169),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1037),
.A2(n_1040),
.B1(n_1085),
.B2(n_1096),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1033),
.B(n_179),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1060),
.A2(n_187),
.A3(n_191),
.B(n_192),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1113),
.A2(n_207),
.B(n_211),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_216),
.B(n_219),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1029),
.A2(n_220),
.B(n_224),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1025),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1047),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1142),
.A2(n_1032),
.B(n_1038),
.C(n_1187),
.Y(n_1214)
);

AO21x1_ASAP7_75t_L g1215 ( 
.A1(n_1145),
.A2(n_1022),
.B(n_1058),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1145),
.A2(n_1174),
.B(n_1116),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1034),
.Y(n_1217)
);

AOI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1022),
.A2(n_1155),
.B(n_1174),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1169),
.B(n_1019),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1092),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1023),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1152),
.B(n_1126),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1018),
.B(n_1024),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1053),
.A2(n_1059),
.B(n_1078),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1116),
.A2(n_1051),
.B(n_1078),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1061),
.A2(n_1083),
.B(n_1080),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1114),
.B(n_1120),
.Y(n_1227)
);

AOI21xp33_ASAP7_75t_L g1228 ( 
.A1(n_1184),
.A2(n_1058),
.B(n_1042),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_1066),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1045),
.A2(n_1148),
.B(n_1044),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1165),
.A2(n_1095),
.A3(n_1202),
.B(n_1143),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1018),
.B(n_1075),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1133),
.B(n_1135),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1043),
.B(n_1062),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1159),
.A2(n_1088),
.B1(n_1170),
.B2(n_1094),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1128),
.A2(n_1121),
.B(n_1093),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1046),
.B(n_1036),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1202),
.A2(n_1101),
.B(n_1110),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1093),
.A2(n_1161),
.B(n_1163),
.Y(n_1239)
);

OAI22x1_ASAP7_75t_L g1240 ( 
.A1(n_1173),
.A2(n_1153),
.B1(n_1175),
.B2(n_1186),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1160),
.A2(n_1041),
.B(n_1193),
.C(n_1069),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1073),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1091),
.A2(n_1084),
.B1(n_1030),
.B2(n_1107),
.Y(n_1243)
);

AOI221x1_ASAP7_75t_L g1244 ( 
.A1(n_1172),
.A2(n_1068),
.B1(n_1154),
.B2(n_1190),
.C(n_1178),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1049),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1107),
.A2(n_1084),
.B1(n_1103),
.B2(n_1129),
.C(n_1134),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_SL g1247 ( 
.A1(n_1138),
.A2(n_1057),
.B(n_1050),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1168),
.B(n_1181),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1026),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1070),
.A2(n_1147),
.B(n_1182),
.C(n_1119),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1064),
.A2(n_1079),
.B(n_1156),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1132),
.B(n_1112),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1074),
.A2(n_1154),
.B(n_1196),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1132),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1027),
.A2(n_1035),
.B(n_1194),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1141),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1127),
.A2(n_1125),
.B(n_1111),
.C(n_1065),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1048),
.A2(n_1109),
.B(n_1124),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1026),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1068),
.A2(n_1151),
.A3(n_1191),
.B(n_1201),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_L g1261 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1077),
.B(n_1081),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1166),
.B(n_1192),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1132),
.B(n_1153),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1056),
.A2(n_1105),
.B(n_1185),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1115),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1047),
.B(n_1183),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1166),
.A2(n_1197),
.B(n_1198),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1067),
.A2(n_1100),
.B(n_1098),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1086),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1139),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1200),
.A2(n_1199),
.B(n_1140),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1054),
.A2(n_1144),
.B(n_1102),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1047),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1118),
.B(n_1144),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1071),
.B(n_1039),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1082),
.A2(n_1020),
.B(n_1099),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1171),
.A2(n_1076),
.B1(n_1164),
.B2(n_1021),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1130),
.B(n_1162),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1056),
.A2(n_1149),
.B(n_1196),
.Y(n_1281)
);

OAI22x1_ASAP7_75t_L g1282 ( 
.A1(n_1076),
.A2(n_1106),
.B1(n_1130),
.B2(n_1162),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1189),
.A2(n_1146),
.B(n_1104),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1177),
.A2(n_1195),
.B(n_1188),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1176),
.A2(n_1180),
.B(n_1131),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1115),
.A2(n_1072),
.B(n_1177),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1115),
.B(n_1122),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1190),
.A2(n_1117),
.B1(n_1052),
.B2(n_1103),
.Y(n_1288)
);

AOI21xp33_ASAP7_75t_L g1289 ( 
.A1(n_1183),
.A2(n_1195),
.B(n_1188),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1195),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1179),
.A2(n_1188),
.B(n_1123),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1072),
.A2(n_1136),
.B(n_1137),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1139),
.B(n_1157),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1031),
.A2(n_1108),
.B(n_1029),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1108),
.A2(n_1029),
.B(n_1142),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1031),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1108),
.A2(n_1037),
.B1(n_1040),
.B2(n_1085),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1063),
.B(n_952),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1150),
.A2(n_1167),
.B(n_1083),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1018),
.B(n_791),
.Y(n_1302)
);

AOI211xp5_ASAP7_75t_L g1303 ( 
.A1(n_1108),
.A2(n_915),
.B(n_955),
.C(n_774),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.C(n_1142),
.Y(n_1305)
);

AOI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1150),
.A2(n_1167),
.B(n_1083),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.C(n_1142),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1025),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1108),
.A2(n_1029),
.B(n_1142),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1024),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.C(n_1142),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1063),
.B(n_952),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1026),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1108),
.A2(n_1142),
.B(n_1085),
.C(n_1096),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1031),
.Y(n_1320)
);

AO21x1_ASAP7_75t_L g1321 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1028),
.B(n_1033),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1150),
.A2(n_1167),
.B(n_1083),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1108),
.B(n_808),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1062),
.B(n_854),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1047),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1108),
.A2(n_1037),
.B1(n_1040),
.B2(n_1085),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1108),
.A2(n_1142),
.B(n_1096),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1047),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1024),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1338)
);

INVx5_ASAP7_75t_L g1339 ( 
.A(n_1115),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1028),
.B(n_1033),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1030),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1028),
.B(n_1033),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1108),
.A2(n_1029),
.B(n_1142),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1108),
.A2(n_600),
.B1(n_1173),
.B2(n_614),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1028),
.B(n_1033),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.C(n_1142),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1145),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1024),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1108),
.A2(n_1029),
.B(n_1142),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1025),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1150),
.A2(n_1055),
.B(n_1053),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1096),
.C(n_1142),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1023),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1108),
.A2(n_1029),
.B(n_1142),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1025),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1023),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1029),
.A2(n_1040),
.B(n_1037),
.Y(n_1361)
);

AOI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_1108),
.A2(n_1142),
.B(n_1096),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1298),
.B(n_1312),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1223),
.B(n_1262),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1329),
.A2(n_1362),
.B(n_1214),
.C(n_1356),
.Y(n_1365)
);

AND2x6_ASAP7_75t_L g1366 ( 
.A(n_1264),
.B(n_1287),
.Y(n_1366)
);

AOI221x1_ASAP7_75t_L g1367 ( 
.A1(n_1329),
.A2(n_1362),
.B1(n_1307),
.B2(n_1311),
.C(n_1348),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1295),
.A2(n_1344),
.B(n_1309),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1297),
.A2(n_1328),
.B1(n_1305),
.B2(n_1335),
.Y(n_1369)
);

AOI222xp33_ASAP7_75t_L g1370 ( 
.A1(n_1345),
.A2(n_1243),
.B1(n_1246),
.B2(n_1297),
.C1(n_1328),
.C2(n_1288),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1294),
.B(n_1323),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1213),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1310),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1296),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1232),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1236),
.A2(n_1322),
.B(n_1317),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1295),
.A2(n_1344),
.B(n_1309),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1342),
.Y(n_1379)
);

OAI21xp33_ASAP7_75t_L g1380 ( 
.A1(n_1351),
.A2(n_1358),
.B(n_1206),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1381)
);

AOI22x1_ASAP7_75t_L g1382 ( 
.A1(n_1351),
.A2(n_1358),
.B1(n_1349),
.B2(n_1361),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1320),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1300),
.A2(n_1304),
.B(n_1301),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1303),
.B(n_1337),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1350),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1285),
.A2(n_1283),
.B(n_1294),
.C(n_1340),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1256),
.B(n_1237),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1266),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1270),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_SL g1391 ( 
.A(n_1318),
.B(n_1335),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1221),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1302),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1336),
.B(n_1206),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1254),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1397)
);

OAI31xp33_ASAP7_75t_L g1398 ( 
.A1(n_1288),
.A2(n_1218),
.A3(n_1228),
.B(n_1235),
.Y(n_1398)
);

AO21x1_ASAP7_75t_L g1399 ( 
.A1(n_1218),
.A2(n_1235),
.B(n_1228),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1346),
.B(n_1222),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1215),
.A2(n_1240),
.B1(n_1279),
.B2(n_1276),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1222),
.B(n_1325),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1212),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1271),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1217),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1252),
.B(n_1220),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1308),
.B(n_1354),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1314),
.A2(n_1338),
.B(n_1319),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1359),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1272),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1225),
.A2(n_1241),
.B(n_1257),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1219),
.A2(n_1203),
.B(n_1283),
.C(n_1250),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1219),
.B(n_1321),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1227),
.B(n_1277),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1276),
.A2(n_1216),
.B1(n_1282),
.B2(n_1357),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1339),
.B(n_1227),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1213),
.B(n_1327),
.Y(n_1419)
);

AND2x6_ASAP7_75t_L g1420 ( 
.A(n_1248),
.B(n_1213),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1242),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1327),
.B(n_1334),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1234),
.B(n_1275),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1280),
.C(n_1293),
.Y(n_1424)
);

AND2x2_ASAP7_75t_SL g1425 ( 
.A(n_1261),
.B(n_1334),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1267),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1290),
.Y(n_1427)
);

OR2x2_ASAP7_75t_SL g1428 ( 
.A(n_1280),
.B(n_1326),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1225),
.A2(n_1265),
.B(n_1244),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1255),
.A2(n_1230),
.B(n_1258),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1360),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1267),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1249),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1285),
.A2(n_1265),
.B1(n_1274),
.B2(n_1281),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1211),
.A2(n_1245),
.B(n_1238),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1226),
.A2(n_1229),
.B(n_1269),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1249),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1278),
.B(n_1209),
.C(n_1291),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1259),
.B(n_1313),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1259),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1313),
.B(n_1284),
.Y(n_1441)
);

INVx8_ASAP7_75t_L g1442 ( 
.A(n_1286),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1289),
.B(n_1253),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1260),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1208),
.A2(n_1204),
.B1(n_1247),
.B2(n_1231),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1208),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1292),
.B(n_1263),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1330),
.A2(n_1355),
.B(n_1353),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1204),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1204),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1273),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1331),
.A2(n_1352),
.B(n_1333),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1251),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1332),
.A2(n_1347),
.B(n_1239),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1210),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1224),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1268),
.B(n_1324),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1299),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1306),
.B(n_1298),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1305),
.A2(n_1108),
.B1(n_1311),
.B2(n_1307),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1223),
.B(n_1262),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1342),
.Y(n_1463)
);

NAND2x1_ASAP7_75t_L g1464 ( 
.A(n_1286),
.B(n_1183),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1266),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1230),
.A2(n_1225),
.B(n_1229),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1342),
.B(n_1062),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1345),
.A2(n_1108),
.B1(n_983),
.B2(n_625),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1342),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1337),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1266),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1233),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1223),
.B(n_1262),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1298),
.B(n_1312),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1296),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1221),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1305),
.B(n_1108),
.C(n_1307),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1337),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1329),
.A2(n_1108),
.B(n_1096),
.C(n_1085),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1213),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1233),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1345),
.A2(n_1108),
.B1(n_983),
.B2(n_625),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1296),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1342),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1213),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1233),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1295),
.A2(n_1358),
.B(n_1351),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1223),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1223),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1214),
.A2(n_1307),
.B(n_1305),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1295),
.A2(n_1358),
.B(n_1351),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1337),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1295),
.A2(n_1358),
.B(n_1351),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1221),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1233),
.Y(n_1503)
);

BUFx4_ASAP7_75t_SL g1504 ( 
.A(n_1296),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1298),
.B(n_1312),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1233),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_SL g1507 ( 
.A1(n_1285),
.A2(n_1142),
.B(n_1108),
.C(n_1295),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1337),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1305),
.A2(n_1108),
.B1(n_1311),
.B2(n_1307),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1337),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1305),
.B(n_1108),
.C(n_1307),
.Y(n_1511)
);

O2A1O1Ixp5_ASAP7_75t_SL g1512 ( 
.A1(n_1329),
.A2(n_1362),
.B(n_1228),
.C(n_1218),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1223),
.B(n_1262),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1213),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1288),
.A2(n_489),
.B1(n_491),
.B2(n_479),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1213),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1266),
.B(n_1339),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1389),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1516),
.A2(n_1370),
.B1(n_1469),
.B2(n_1487),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1479),
.A2(n_1511),
.B1(n_1369),
.B2(n_1460),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1405),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1370),
.A2(n_1371),
.B1(n_1398),
.B2(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1407),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1459),
.B(n_1380),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1377),
.A2(n_1452),
.B(n_1448),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1394),
.A2(n_1369),
.B1(n_1511),
.B2(n_1397),
.Y(n_1528)
);

CKINVDCx6p67_ASAP7_75t_R g1529 ( 
.A(n_1383),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1411),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1412),
.A2(n_1401),
.B1(n_1498),
.B2(n_1428),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1454),
.A2(n_1436),
.B(n_1430),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1421),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1444),
.Y(n_1534)
);

AOI222xp33_ASAP7_75t_L g1535 ( 
.A1(n_1380),
.A2(n_1498),
.B1(n_1385),
.B2(n_1363),
.C1(n_1505),
.C2(n_1476),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1420),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1398),
.A2(n_1509),
.B1(n_1399),
.B2(n_1391),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1449),
.A2(n_1478),
.B1(n_1392),
.B2(n_1406),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1420),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1366),
.A2(n_1400),
.B1(n_1413),
.B2(n_1443),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1477),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1431),
.Y(n_1542)
);

BUFx2_ASAP7_75t_R g1543 ( 
.A(n_1463),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1365),
.A2(n_1482),
.B1(n_1499),
.B2(n_1501),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1507),
.A2(n_1378),
.B(n_1368),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1502),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1420),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1389),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1389),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1504),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1429),
.Y(n_1551)
);

BUFx2_ASAP7_75t_SL g1552 ( 
.A(n_1470),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1415),
.A2(n_1435),
.B(n_1450),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1465),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1366),
.A2(n_1496),
.B1(n_1376),
.B2(n_1497),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1474),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1429),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1386),
.Y(n_1558)
);

INVx4_ASAP7_75t_SL g1559 ( 
.A(n_1366),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1374),
.B(n_1381),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1472),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1441),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1480),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1468),
.Y(n_1564)
);

AOI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1410),
.A2(n_1384),
.B(n_1457),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1395),
.B(n_1402),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1496),
.A2(n_1376),
.B1(n_1471),
.B2(n_1513),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1441),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1375),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1488),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1486),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1495),
.A2(n_1492),
.B1(n_1414),
.B2(n_1404),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1456),
.Y(n_1573)
);

CKINVDCx11_ASAP7_75t_R g1574 ( 
.A(n_1379),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1364),
.B(n_1462),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1393),
.A2(n_1416),
.B1(n_1417),
.B2(n_1514),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1494),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1503),
.Y(n_1578)
);

CKINVDCx9p33_ASAP7_75t_R g1579 ( 
.A(n_1490),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1506),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1475),
.B(n_1373),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1458),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1427),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1408),
.B(n_1512),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1423),
.Y(n_1585)
);

CKINVDCx6p67_ASAP7_75t_R g1586 ( 
.A(n_1437),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1388),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1458),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1372),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1372),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_1500),
.Y(n_1591)
);

INVx4_ASAP7_75t_SL g1592 ( 
.A(n_1402),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1439),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1517),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1446),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1508),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1372),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1467),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1465),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1396),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1510),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1434),
.A2(n_1382),
.B1(n_1437),
.B2(n_1390),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1517),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1425),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1485),
.B(n_1515),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1485),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1367),
.A2(n_1438),
.B(n_1387),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1396),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1485),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1418),
.B(n_1432),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1493),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1403),
.B(n_1461),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1493),
.Y(n_1613)
);

BUFx2_ASAP7_75t_R g1614 ( 
.A(n_1419),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1491),
.A2(n_1473),
.B1(n_1437),
.B2(n_1440),
.Y(n_1615)
);

CKINVDCx11_ASAP7_75t_R g1616 ( 
.A(n_1493),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1403),
.B(n_1461),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1515),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1515),
.Y(n_1619)
);

OAI21xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1455),
.A2(n_1491),
.B(n_1447),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1473),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1466),
.B(n_1519),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1467),
.A2(n_1438),
.B(n_1453),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1426),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1426),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1426),
.B(n_1440),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1433),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1424),
.A2(n_1445),
.B(n_1489),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1447),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1433),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1447),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1433),
.Y(n_1632)
);

AOI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1451),
.A2(n_1464),
.B(n_1518),
.Y(n_1633)
);

AO21x1_ASAP7_75t_L g1634 ( 
.A1(n_1455),
.A2(n_1445),
.B(n_1484),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1440),
.A2(n_1466),
.B(n_1481),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1442),
.A2(n_1483),
.B(n_1489),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1442),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1483),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1363),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1479),
.A2(n_1108),
.B1(n_1303),
.B2(n_1511),
.Y(n_1640)
);

CKINVDCx11_ASAP7_75t_R g1641 ( 
.A(n_1383),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1425),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1430),
.A2(n_1384),
.B(n_1410),
.Y(n_1643)
);

BUFx8_ASAP7_75t_SL g1644 ( 
.A(n_1383),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1479),
.A2(n_1108),
.B1(n_1303),
.B2(n_1511),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1420),
.Y(n_1646)
);

AOI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1371),
.A2(n_1452),
.B(n_1448),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1425),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1377),
.A2(n_1452),
.B(n_1448),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1389),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1386),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_SL g1652 ( 
.A(n_1477),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1420),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1425),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1409),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1409),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1409),
.Y(n_1657)
);

AOI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1371),
.A2(n_1452),
.B(n_1448),
.Y(n_1658)
);

AO21x1_ASAP7_75t_L g1659 ( 
.A1(n_1398),
.A2(n_1309),
.B(n_1295),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1377),
.A2(n_1452),
.B(n_1448),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1420),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1409),
.Y(n_1662)
);

CKINVDCx11_ASAP7_75t_R g1663 ( 
.A(n_1383),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1409),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1425),
.Y(n_1665)
);

BUFx4f_ASAP7_75t_SL g1666 ( 
.A(n_1375),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1409),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1442),
.B(n_1491),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1420),
.Y(n_1669)
);

AOI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1371),
.A2(n_1452),
.B(n_1448),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1373),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1516),
.A2(n_1345),
.B1(n_1370),
.B2(n_1108),
.Y(n_1672)
);

INVx3_ASAP7_75t_SL g1673 ( 
.A(n_1477),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1412),
.Y(n_1674)
);

AO21x1_ASAP7_75t_SL g1675 ( 
.A1(n_1498),
.A2(n_1218),
.B(n_1228),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1386),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1363),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1516),
.A2(n_1345),
.B1(n_1370),
.B2(n_1108),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1422),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1523),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1631),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1536),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1526),
.B(n_1551),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1559),
.B(n_1562),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1631),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1671),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1532),
.A2(n_1607),
.B(n_1545),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1561),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1563),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1548),
.Y(n_1690)
);

AOI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1647),
.A2(n_1670),
.B(n_1658),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1525),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1659),
.A2(n_1553),
.B(n_1584),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1659),
.A2(n_1553),
.B(n_1584),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1527),
.A2(n_1660),
.B(n_1649),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1537),
.A2(n_1524),
.B(n_1640),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1676),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1560),
.B(n_1528),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1557),
.B(n_1581),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1616),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1644),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1558),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1532),
.A2(n_1565),
.B(n_1623),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1556),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1539),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1571),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1577),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1582),
.B(n_1588),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1578),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1596),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1672),
.A2(n_1678),
.B1(n_1521),
.B2(n_1535),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1580),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1530),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1598),
.A2(n_1595),
.B(n_1544),
.Y(n_1717)
);

AOI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1522),
.A2(n_1602),
.B(n_1645),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1533),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1601),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1616),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1657),
.B(n_1662),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1664),
.B(n_1667),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1542),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1583),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1593),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1727)
);

AO21x2_ASAP7_75t_L g1728 ( 
.A1(n_1634),
.A2(n_1534),
.B(n_1633),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1562),
.B(n_1568),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1573),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1568),
.B(n_1587),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1589),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1573),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1568),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1628),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1628),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1559),
.B(n_1547),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1628),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1675),
.B(n_1585),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1643),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1639),
.B(n_1677),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1646),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1643),
.Y(n_1743)
);

BUFx8_ASAP7_75t_L g1744 ( 
.A(n_1569),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1643),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1546),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1540),
.B(n_1605),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1605),
.B(n_1591),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1653),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1653),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1567),
.B(n_1608),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1626),
.B(n_1661),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1661),
.Y(n_1753)
);

AO21x1_ASAP7_75t_SL g1754 ( 
.A1(n_1627),
.A2(n_1630),
.B(n_1603),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1669),
.B(n_1594),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1586),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1600),
.B(n_1576),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1620),
.Y(n_1758)
);

OR2x6_ASAP7_75t_L g1759 ( 
.A(n_1668),
.B(n_1636),
.Y(n_1759)
);

AOI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1606),
.A2(n_1619),
.B(n_1609),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1624),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1625),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1600),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1638),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1613),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1586),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1520),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1618),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1589),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1531),
.B(n_1665),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1590),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1590),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1674),
.B(n_1673),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1590),
.B(n_1611),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1597),
.B(n_1611),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1597),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1604),
.B(n_1642),
.Y(n_1778)
);

AO21x2_ASAP7_75t_L g1779 ( 
.A1(n_1615),
.A2(n_1610),
.B(n_1635),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1642),
.B(n_1654),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1599),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1538),
.A2(n_1555),
.B(n_1612),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1768),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1716),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1716),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1701),
.B(n_1552),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1705),
.A2(n_1612),
.B(n_1622),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1719),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1719),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1683),
.B(n_1679),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1713),
.A2(n_1648),
.B1(n_1654),
.B2(n_1665),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1705),
.A2(n_1612),
.B(n_1622),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1681),
.Y(n_1794)
);

INVxp67_ASAP7_75t_SL g1795 ( 
.A(n_1686),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1774),
.B(n_1529),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_L g1797 ( 
.A(n_1758),
.B(n_1520),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1701),
.B(n_1648),
.Y(n_1798)
);

NOR2xp67_ASAP7_75t_L g1799 ( 
.A(n_1758),
.B(n_1554),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1700),
.A2(n_1637),
.B1(n_1674),
.B2(n_1564),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1717),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1729),
.B(n_1731),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1717),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1731),
.B(n_1622),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1732),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1694),
.B(n_1696),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1727),
.B(n_1554),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1694),
.B(n_1617),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1694),
.B(n_1617),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1688),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1696),
.B(n_1617),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1730),
.B(n_1529),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1685),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1726),
.B(n_1549),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1685),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1730),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1739),
.B(n_1566),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1689),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1767),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1706),
.B(n_1549),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1733),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1739),
.B(n_1566),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1687),
.B(n_1566),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1695),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1767),
.Y(n_1825)
);

AOI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1698),
.A2(n_1650),
.B(n_1548),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1708),
.B(n_1621),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1687),
.B(n_1574),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1687),
.B(n_1574),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1709),
.B(n_1711),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1759),
.B(n_1592),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1769),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1687),
.B(n_1734),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1718),
.A2(n_1637),
.B1(n_1564),
.B2(n_1543),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1699),
.Y(n_1835)
);

AOI222xp33_ASAP7_75t_L g1836 ( 
.A1(n_1757),
.A2(n_1570),
.B1(n_1569),
.B2(n_1666),
.C1(n_1663),
.C2(n_1641),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1733),
.B(n_1710),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1714),
.B(n_1621),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1712),
.B(n_1650),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1720),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1704),
.Y(n_1841)
);

AND2x2_ASAP7_75t_SL g1842 ( 
.A(n_1684),
.B(n_1737),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_SL g1843 ( 
.A(n_1754),
.B(n_1759),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1749),
.Y(n_1844)
);

NAND4xp25_ASAP7_75t_L g1845 ( 
.A(n_1836),
.B(n_1741),
.C(n_1702),
.D(n_1721),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1830),
.Y(n_1846)
);

NAND4xp25_ASAP7_75t_L g1847 ( 
.A(n_1836),
.B(n_1741),
.C(n_1702),
.D(n_1721),
.Y(n_1847)
);

OAI21xp33_ASAP7_75t_L g1848 ( 
.A1(n_1806),
.A2(n_1718),
.B(n_1766),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1795),
.B(n_1725),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1795),
.B(n_1680),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1821),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1840),
.B(n_1693),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1810),
.B(n_1715),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1802),
.B(n_1748),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1802),
.B(n_1748),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1818),
.B(n_1722),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1801),
.A2(n_1743),
.B(n_1745),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1823),
.B(n_1747),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1797),
.B(n_1690),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1824),
.B(n_1723),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1834),
.B(n_1763),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1841),
.B(n_1766),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1783),
.B(n_1744),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1724),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1823),
.B(n_1747),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1835),
.B(n_1770),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1832),
.B(n_1761),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1834),
.A2(n_1771),
.B(n_1777),
.Y(n_1868)
);

NOR3xp33_ASAP7_75t_L g1869 ( 
.A(n_1800),
.B(n_1777),
.C(n_1749),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1828),
.B(n_1752),
.Y(n_1870)
);

NAND3xp33_ASAP7_75t_L g1871 ( 
.A(n_1806),
.B(n_1738),
.C(n_1736),
.Y(n_1871)
);

NAND3xp33_ASAP7_75t_L g1872 ( 
.A(n_1807),
.B(n_1814),
.C(n_1820),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1832),
.B(n_1761),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1807),
.B(n_1805),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_L g1875 ( 
.A(n_1814),
.B(n_1738),
.C(n_1736),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1828),
.A2(n_1771),
.B(n_1744),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1791),
.B(n_1754),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1829),
.A2(n_1744),
.B(n_1768),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1805),
.B(n_1762),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1829),
.B(n_1755),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1820),
.B(n_1735),
.C(n_1762),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_L g1882 ( 
.A(n_1812),
.B(n_1756),
.C(n_1740),
.D(n_1745),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1735),
.C(n_1753),
.Y(n_1883)
);

NAND3xp33_ASAP7_75t_L g1884 ( 
.A(n_1833),
.B(n_1750),
.C(n_1753),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1792),
.A2(n_1751),
.B1(n_1764),
.B2(n_1778),
.C(n_1780),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1843),
.A2(n_1782),
.B1(n_1779),
.B2(n_1751),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1797),
.B(n_1690),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1794),
.B(n_1772),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1830),
.Y(n_1889)
);

NAND3xp33_ASAP7_75t_L g1890 ( 
.A(n_1827),
.B(n_1773),
.C(n_1765),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1800),
.A2(n_1782),
.B1(n_1765),
.B2(n_1779),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1804),
.B(n_1808),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1815),
.B(n_1787),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1804),
.B(n_1728),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_L g1895 ( 
.A(n_1839),
.B(n_1756),
.C(n_1760),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1808),
.B(n_1728),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1815),
.B(n_1775),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1821),
.B(n_1776),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1812),
.A2(n_1756),
.B1(n_1614),
.B2(n_1682),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1837),
.B(n_1776),
.Y(n_1900)
);

OAI21xp33_ASAP7_75t_L g1901 ( 
.A1(n_1816),
.A2(n_1838),
.B(n_1813),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1803),
.A2(n_1743),
.B(n_1740),
.Y(n_1902)
);

OA21x2_ASAP7_75t_L g1903 ( 
.A1(n_1803),
.A2(n_1697),
.B(n_1691),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1826),
.A2(n_1782),
.B1(n_1779),
.B2(n_1746),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1799),
.B(n_1690),
.Y(n_1905)
);

NAND2xp33_ASAP7_75t_SL g1906 ( 
.A(n_1784),
.B(n_1550),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_R g1907 ( 
.A(n_1842),
.B(n_1550),
.Y(n_1907)
);

OA211x2_ASAP7_75t_L g1908 ( 
.A1(n_1796),
.A2(n_1579),
.B(n_1570),
.C(n_1663),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1809),
.B(n_1728),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1785),
.B(n_1786),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1809),
.B(n_1692),
.Y(n_1911)
);

AOI211xp5_ASAP7_75t_L g1912 ( 
.A1(n_1826),
.A2(n_1707),
.B(n_1742),
.C(n_1781),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1851),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1858),
.B(n_1788),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1858),
.B(n_1788),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1846),
.B(n_1816),
.Y(n_1916)
);

AND2x2_ASAP7_75t_SL g1917 ( 
.A(n_1891),
.B(n_1842),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1889),
.B(n_1816),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1848),
.B(n_1850),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1865),
.B(n_1892),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1888),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1907),
.Y(n_1922)
);

AND4x1_ASAP7_75t_L g1923 ( 
.A(n_1863),
.B(n_1839),
.C(n_1822),
.D(n_1817),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1865),
.B(n_1788),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1857),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1871),
.B(n_1831),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1910),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1857),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1870),
.B(n_1843),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1892),
.B(n_1788),
.Y(n_1930)
);

AND2x4_ASAP7_75t_SL g1931 ( 
.A(n_1877),
.B(n_1831),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1849),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1883),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1854),
.B(n_1793),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1857),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1854),
.B(n_1855),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1855),
.B(n_1793),
.Y(n_1937)
);

OR2x6_ASAP7_75t_L g1938 ( 
.A(n_1896),
.B(n_1831),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1852),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1902),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1902),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1845),
.B(n_1819),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1870),
.B(n_1793),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1894),
.B(n_1793),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1880),
.B(n_1811),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1903),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1903),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1862),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1907),
.B(n_1912),
.Y(n_1949)
);

NAND2x1p5_ASAP7_75t_L g1950 ( 
.A(n_1859),
.B(n_1831),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1884),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1872),
.B(n_1798),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1909),
.B(n_1844),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1853),
.B(n_1798),
.Y(n_1954)
);

NAND2x1p5_ASAP7_75t_L g1955 ( 
.A(n_1887),
.B(n_1905),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1903),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1867),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1856),
.B(n_1860),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1895),
.B(n_1785),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1881),
.B(n_1786),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1911),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1906),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1873),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1951),
.B(n_1869),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1916),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1920),
.B(n_1893),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1925),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1951),
.B(n_1900),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1920),
.B(n_1874),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_1864),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1920),
.B(n_1819),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1916),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1918),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1918),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1938),
.B(n_1875),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1936),
.B(n_1825),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1936),
.B(n_1825),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1931),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1960),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1960),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1945),
.B(n_1825),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1942),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1913),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1925),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1931),
.Y(n_1985)
);

OAI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1933),
.A2(n_1861),
.B(n_1868),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1948),
.B(n_1879),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_1959),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1945),
.B(n_1861),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1942),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1959),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1919),
.B(n_1866),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1927),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1932),
.B(n_1890),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1919),
.B(n_1898),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1958),
.B(n_1897),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1925),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1932),
.B(n_1901),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1939),
.B(n_1789),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1917),
.A2(n_1891),
.B(n_1886),
.C(n_1876),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1939),
.B(n_1789),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1945),
.B(n_1817),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1929),
.B(n_1822),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1927),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1957),
.B(n_1790),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1925),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1957),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1962),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1963),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1928),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1931),
.Y(n_2011)
);

OR2x6_ASAP7_75t_L g2012 ( 
.A(n_1938),
.B(n_1759),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1963),
.B(n_1790),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_L g2014 ( 
.A(n_1986),
.B(n_1933),
.C(n_1917),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1970),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1986),
.B(n_1847),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1996),
.B(n_1958),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1988),
.B(n_1958),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1989),
.B(n_1962),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1988),
.B(n_1952),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2000),
.A2(n_1917),
.B1(n_1949),
.B2(n_1904),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1999),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1996),
.B(n_1954),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1989),
.B(n_1962),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1978),
.B(n_1934),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1968),
.B(n_1954),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1978),
.B(n_1934),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1991),
.B(n_1952),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1991),
.B(n_1968),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2001),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1964),
.B(n_1923),
.Y(n_2031)
);

INVxp67_ASAP7_75t_SL g2032 ( 
.A(n_2008),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1979),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1979),
.B(n_1952),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1967),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1980),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1967),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1985),
.B(n_1934),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1980),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2005),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1967),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2013),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1969),
.B(n_1921),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1985),
.B(n_1937),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1995),
.B(n_1954),
.Y(n_2045)
);

AOI21xp33_ASAP7_75t_L g2046 ( 
.A1(n_1982),
.A2(n_1917),
.B(n_1926),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1984),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2011),
.B(n_1937),
.Y(n_2048)
);

CKINVDCx16_ASAP7_75t_R g2049 ( 
.A(n_2008),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1984),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1993),
.Y(n_2051)
);

INVx3_ASAP7_75t_SL g2052 ( 
.A(n_2011),
.Y(n_2052)
);

INVxp67_ASAP7_75t_L g2053 ( 
.A(n_1983),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1969),
.B(n_1921),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1994),
.B(n_1953),
.Y(n_2055)
);

NAND2x1_ASAP7_75t_L g2056 ( 
.A(n_1971),
.B(n_1929),
.Y(n_2056)
);

NAND2x1p5_ASAP7_75t_L g2057 ( 
.A(n_1975),
.B(n_1923),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1990),
.B(n_1913),
.C(n_1949),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1993),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2002),
.B(n_1937),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_1992),
.B(n_1961),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2004),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1965),
.B(n_1972),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_1998),
.Y(n_2064)
);

INVx1_ASAP7_75t_SL g2065 ( 
.A(n_2052),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_2057),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2045),
.B(n_1965),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2045),
.B(n_1972),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2019),
.B(n_2002),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2051),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_2032),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2017),
.B(n_1973),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2026),
.B(n_1973),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_2057),
.A2(n_1997),
.B(n_1984),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2023),
.B(n_1974),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2033),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2059),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2062),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2036),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2035),
.Y(n_2080)
);

INVxp67_ASAP7_75t_SL g2081 ( 
.A(n_2016),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2016),
.A2(n_1922),
.B1(n_1926),
.B2(n_1992),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2031),
.B(n_1644),
.Y(n_2083)
);

AOI31xp33_ASAP7_75t_L g2084 ( 
.A1(n_2014),
.A2(n_1955),
.A3(n_1950),
.B(n_1899),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2039),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2018),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2018),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_2049),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2029),
.B(n_1974),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2064),
.B(n_1966),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_2052),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2019),
.B(n_2003),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_2021),
.A2(n_1975),
.B1(n_1904),
.B2(n_1926),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2035),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2024),
.B(n_2003),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_2053),
.Y(n_2096)
);

AO21x2_ASAP7_75t_L g2097 ( 
.A1(n_2037),
.A2(n_2006),
.B(n_1997),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2024),
.B(n_1966),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2060),
.B(n_1981),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2015),
.B(n_2007),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2063),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_L g2102 ( 
.A(n_2058),
.B(n_1922),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2020),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2034),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2031),
.A2(n_1926),
.B1(n_1975),
.B2(n_1950),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2097),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2070),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2090),
.B(n_2029),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2081),
.B(n_2104),
.Y(n_2109)
);

AOI322xp5_ASAP7_75t_L g2110 ( 
.A1(n_2093),
.A2(n_2102),
.A3(n_2103),
.B1(n_2088),
.B2(n_2086),
.C1(n_2087),
.C2(n_2066),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2071),
.B(n_2022),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_2088),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2074),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2070),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2084),
.A2(n_2028),
.B(n_2020),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2071),
.B(n_2030),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2077),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2103),
.B(n_2043),
.Y(n_2118)
);

OAI321xp33_ASAP7_75t_L g2119 ( 
.A1(n_2082),
.A2(n_2028),
.A3(n_2055),
.B1(n_1926),
.B2(n_2054),
.C(n_2012),
.Y(n_2119)
);

OAI21xp33_ASAP7_75t_L g2120 ( 
.A1(n_2065),
.A2(n_2042),
.B(n_2040),
.Y(n_2120)
);

OAI31xp33_ASAP7_75t_L g2121 ( 
.A1(n_2066),
.A2(n_2046),
.A3(n_1975),
.B(n_1944),
.Y(n_2121)
);

AOI21xp5_ASAP7_75t_SL g2122 ( 
.A1(n_2083),
.A2(n_1926),
.B(n_2061),
.Y(n_2122)
);

OAI32xp33_ASAP7_75t_L g2123 ( 
.A1(n_2066),
.A2(n_1947),
.A3(n_1946),
.B1(n_1995),
.B2(n_2048),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2091),
.B(n_1641),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2086),
.B(n_2007),
.Y(n_2125)
);

OAI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2087),
.A2(n_1926),
.B1(n_1882),
.B2(n_1885),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2098),
.B(n_2009),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_2096),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2098),
.B(n_2060),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2077),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2074),
.A2(n_2105),
.B1(n_2080),
.B2(n_2094),
.Y(n_2131)
);

A2O1A1Ixp33_ASAP7_75t_L g2132 ( 
.A1(n_2096),
.A2(n_1944),
.B(n_1915),
.C(n_1924),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2069),
.Y(n_2133)
);

A2O1A1Ixp33_ASAP7_75t_L g2134 ( 
.A1(n_2101),
.A2(n_1944),
.B(n_1915),
.C(n_1924),
.Y(n_2134)
);

AOI221xp5_ASAP7_75t_L g2135 ( 
.A1(n_2101),
.A2(n_1946),
.B1(n_1947),
.B2(n_1956),
.C(n_2047),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_2076),
.B(n_2025),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2128),
.B(n_2069),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2107),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2109),
.Y(n_2139)
);

OAI221xp5_ASAP7_75t_L g2140 ( 
.A1(n_2115),
.A2(n_2089),
.B1(n_2100),
.B2(n_2068),
.C(n_2067),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2129),
.B(n_2092),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_2124),
.B(n_2112),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2106),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2124),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_2110),
.B(n_2089),
.Y(n_2145)
);

NAND2xp33_ASAP7_75t_L g2146 ( 
.A(n_2120),
.B(n_2067),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2133),
.B(n_2092),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2114),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2117),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2130),
.Y(n_2150)
);

AOI222xp33_ASAP7_75t_L g2151 ( 
.A1(n_2126),
.A2(n_2080),
.B1(n_2094),
.B2(n_2085),
.C1(n_2079),
.C2(n_1928),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2106),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2108),
.B(n_2095),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_2136),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2111),
.B(n_2095),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2125),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2136),
.B(n_2099),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_2116),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2118),
.Y(n_2159)
);

INVxp67_ASAP7_75t_SL g2160 ( 
.A(n_2113),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2122),
.B(n_2068),
.Y(n_2161)
);

OAI21xp5_ASAP7_75t_SL g2162 ( 
.A1(n_2145),
.A2(n_2126),
.B(n_2121),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_2144),
.B(n_2119),
.Y(n_2163)
);

AOI221x1_ASAP7_75t_SL g2164 ( 
.A1(n_2137),
.A2(n_2127),
.B1(n_2079),
.B2(n_2085),
.C(n_2078),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2141),
.Y(n_2165)
);

AOI221xp5_ASAP7_75t_L g2166 ( 
.A1(n_2145),
.A2(n_2140),
.B1(n_2160),
.B2(n_2146),
.C(n_2154),
.Y(n_2166)
);

AOI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_2146),
.A2(n_2154),
.B(n_2161),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2151),
.A2(n_2131),
.B(n_2135),
.Y(n_2168)
);

AOI322xp5_ASAP7_75t_L g2169 ( 
.A1(n_2139),
.A2(n_2132),
.A3(n_2134),
.B1(n_2037),
.B2(n_2050),
.C1(n_2041),
.C2(n_2047),
.Y(n_2169)
);

OAI221xp5_ASAP7_75t_SL g2170 ( 
.A1(n_2158),
.A2(n_2157),
.B1(n_2159),
.B2(n_2132),
.C(n_2144),
.Y(n_2170)
);

AOI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2156),
.A2(n_2123),
.B1(n_2134),
.B2(n_2078),
.C(n_2041),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_SL g2172 ( 
.A(n_2142),
.B(n_2072),
.C(n_2075),
.Y(n_2172)
);

OAI21xp33_ASAP7_75t_L g2173 ( 
.A1(n_2157),
.A2(n_2072),
.B(n_2073),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_2153),
.A2(n_2097),
.B1(n_2050),
.B2(n_2006),
.Y(n_2174)
);

NOR3xp33_ASAP7_75t_L g2175 ( 
.A(n_2155),
.B(n_2075),
.C(n_2073),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2141),
.B(n_2099),
.Y(n_2176)
);

NAND4xp25_ASAP7_75t_L g2177 ( 
.A(n_2166),
.B(n_2147),
.C(n_2148),
.D(n_2138),
.Y(n_2177)
);

NOR3xp33_ASAP7_75t_L g2178 ( 
.A(n_2163),
.B(n_2143),
.C(n_2152),
.Y(n_2178)
);

NAND3xp33_ASAP7_75t_L g2179 ( 
.A(n_2170),
.B(n_2150),
.C(n_2149),
.Y(n_2179)
);

NOR2x1_ASAP7_75t_L g2180 ( 
.A(n_2172),
.B(n_2143),
.Y(n_2180)
);

NOR2x1_ASAP7_75t_L g2181 ( 
.A(n_2167),
.B(n_2152),
.Y(n_2181)
);

NAND3xp33_ASAP7_75t_L g2182 ( 
.A(n_2162),
.B(n_2006),
.C(n_1997),
.Y(n_2182)
);

CKINVDCx6p67_ASAP7_75t_R g2183 ( 
.A(n_2176),
.Y(n_2183)
);

NAND4xp75_ASAP7_75t_L g2184 ( 
.A(n_2168),
.B(n_1908),
.C(n_2027),
.D(n_2025),
.Y(n_2184)
);

NOR2x1_ASAP7_75t_L g2185 ( 
.A(n_2165),
.B(n_2056),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2173),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2174),
.Y(n_2187)
);

NAND4xp75_ASAP7_75t_L g2188 ( 
.A(n_2171),
.B(n_2027),
.C(n_2044),
.D(n_2038),
.Y(n_2188)
);

NAND4xp75_ASAP7_75t_L g2189 ( 
.A(n_2164),
.B(n_2038),
.C(n_2048),
.D(n_2044),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2183),
.B(n_2175),
.Y(n_2190)
);

AND4x1_ASAP7_75t_L g2191 ( 
.A(n_2181),
.B(n_2179),
.C(n_2180),
.D(n_2178),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2177),
.B(n_1652),
.Y(n_2192)
);

NOR4xp25_ASAP7_75t_L g2193 ( 
.A(n_2186),
.B(n_2169),
.C(n_2010),
.D(n_2009),
.Y(n_2193)
);

AND4x1_ASAP7_75t_L g2194 ( 
.A(n_2185),
.B(n_1541),
.C(n_1981),
.D(n_1971),
.Y(n_2194)
);

NOR3x1_ASAP7_75t_L g2195 ( 
.A(n_2188),
.B(n_1878),
.C(n_1541),
.Y(n_2195)
);

A2O1A1Ixp33_ASAP7_75t_L g2196 ( 
.A1(n_2187),
.A2(n_2010),
.B(n_1947),
.C(n_1946),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2189),
.B(n_2004),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2190),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2191),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2195),
.B(n_2184),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2192),
.A2(n_2182),
.B1(n_2097),
.B2(n_2010),
.Y(n_2201)
);

NOR2xp67_ASAP7_75t_L g2202 ( 
.A(n_2197),
.B(n_2194),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2193),
.A2(n_1956),
.B1(n_1914),
.B2(n_1924),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2196),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2191),
.B(n_1987),
.Y(n_2205)
);

NOR2xp67_ASAP7_75t_SL g2206 ( 
.A(n_2199),
.B(n_1690),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_2202),
.B(n_2204),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2198),
.B(n_1946),
.Y(n_2208)
);

INVx1_ASAP7_75t_SL g2209 ( 
.A(n_2200),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2205),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2201),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2203),
.B(n_1946),
.Y(n_2212)
);

INVx1_ASAP7_75t_SL g2213 ( 
.A(n_2209),
.Y(n_2213)
);

XOR2x1_ASAP7_75t_L g2214 ( 
.A(n_2210),
.B(n_2211),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_2208),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2207),
.Y(n_2216)
);

INVxp67_ASAP7_75t_SL g2217 ( 
.A(n_2214),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2213),
.A2(n_2212),
.B1(n_2206),
.B2(n_1947),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_2217),
.B(n_2216),
.C(n_2215),
.Y(n_2219)
);

NOR2x1_ASAP7_75t_L g2220 ( 
.A(n_2218),
.B(n_2215),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_2219),
.A2(n_1956),
.B1(n_1947),
.B2(n_1935),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2220),
.Y(n_2222)
);

OAI22x1_ASAP7_75t_L g2223 ( 
.A1(n_2219),
.A2(n_1955),
.B1(n_1950),
.B2(n_1977),
.Y(n_2223)
);

OAI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2222),
.A2(n_1956),
.B(n_1915),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2221),
.B(n_1928),
.Y(n_2225)
);

OAI21xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2224),
.A2(n_2223),
.B(n_1976),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2225),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2227),
.B(n_1928),
.Y(n_2228)
);

AOI222xp33_ASAP7_75t_L g2229 ( 
.A1(n_2228),
.A2(n_2226),
.B1(n_1940),
.B2(n_1941),
.C1(n_1935),
.C2(n_1930),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2229),
.A2(n_1935),
.B1(n_1941),
.B2(n_1940),
.Y(n_2230)
);

AOI211xp5_ASAP7_75t_L g2231 ( 
.A1(n_2230),
.A2(n_1930),
.B(n_1943),
.C(n_1914),
.Y(n_2231)
);


endmodule