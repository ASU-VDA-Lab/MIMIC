module fake_jpeg_25867_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_29),
.C(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_20),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_36),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_40),
.C(n_38),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_16),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_38),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_11),
.C(n_4),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_72),
.B(n_12),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_20),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_14),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_57),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_62),
.C(n_54),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_15),
.C(n_11),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_82),
.B1(n_12),
.B2(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_14),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_74),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_85),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_68),
.B1(n_35),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_87),
.B1(n_84),
.B2(n_88),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_80),
.B1(n_52),
.B2(n_33),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_15),
.C(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_52),
.B1(n_18),
.B2(n_15),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_30),
.C(n_5),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_10),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_91),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_3),
.B(n_8),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_93),
.B(n_6),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_3),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_10),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule