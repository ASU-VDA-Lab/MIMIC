module real_aes_9803_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_102;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
wire n_91;
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_0), .A2(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g652 ( .A(n_0), .Y(n_652) );
INVx1_ASAP7_75t_L g138 ( .A(n_1), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_2), .B(n_61), .Y(n_509) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_2), .Y(n_597) );
INVx1_ASAP7_75t_L g635 ( .A(n_2), .Y(n_635) );
AND2x2_ASAP7_75t_L g651 ( .A(n_2), .B(n_634), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_3), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_4), .B(n_159), .Y(n_232) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_5), .A2(n_526), .B1(n_532), .B2(n_545), .C(n_556), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_5), .A2(n_54), .B1(n_604), .B2(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g518 ( .A(n_6), .Y(n_518) );
OR2x2_ASAP7_75t_L g531 ( .A(n_6), .B(n_516), .Y(n_531) );
OR2x2_ASAP7_75t_L g508 ( .A(n_7), .B(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g512 ( .A(n_7), .Y(n_512) );
BUFx2_ASAP7_75t_L g591 ( .A(n_7), .Y(n_591) );
INVx1_ASAP7_75t_L g650 ( .A(n_7), .Y(n_650) );
INVx1_ASAP7_75t_L g487 ( .A(n_8), .Y(n_487) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_9), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_10), .A2(n_43), .B1(n_542), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g655 ( .A(n_10), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_11), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_12), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_13), .B(n_198), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_14), .A2(n_54), .B1(n_584), .B2(n_585), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_14), .A2(n_73), .B1(n_610), .B2(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_15), .B(n_123), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_15), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_16), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_17), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_18), .B(n_116), .Y(n_202) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_20), .B(n_118), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_21), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_22), .B(n_123), .Y(n_231) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
OAI21xp33_ASAP7_75t_L g181 ( .A1(n_24), .A2(n_144), .B(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_25), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_26), .A2(n_498), .B1(n_499), .B2(n_682), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_26), .Y(n_682) );
INVx1_ASAP7_75t_L g516 ( .A(n_27), .Y(n_516) );
INVx1_ASAP7_75t_L g555 ( .A(n_27), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_28), .B(n_116), .Y(n_226) );
INVx1_ASAP7_75t_L g546 ( .A(n_29), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_29), .A2(n_50), .B1(n_600), .B2(n_604), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_30), .Y(n_168) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_31), .Y(n_490) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_32), .A2(n_55), .B(n_112), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_33), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_34), .B(n_116), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_35), .Y(n_246) );
AND2x6_ASAP7_75t_L g83 ( .A(n_36), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_36), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_36), .B(n_668), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_37), .A2(n_65), .B1(n_159), .B2(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_38), .B(n_172), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_39), .Y(n_161) );
INVx1_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_40), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_41), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_42), .B(n_184), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_43), .A2(n_72), .B1(n_657), .B2(n_659), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_44), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_45), .B(n_184), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_46), .B(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_47), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_48), .B(n_172), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_49), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g540 ( .A(n_50), .Y(n_540) );
INVx2_ASAP7_75t_L g150 ( .A(n_51), .Y(n_150) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_52), .A2(n_551), .B(n_553), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_52), .A2(n_71), .B1(n_610), .B2(n_616), .Y(n_609) );
INVx2_ASAP7_75t_L g507 ( .A(n_53), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_56), .B(n_124), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_57), .Y(n_564) );
INVx1_ASAP7_75t_L g142 ( .A(n_58), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_59), .Y(n_254) );
BUFx10_ASAP7_75t_L g677 ( .A(n_60), .Y(n_677) );
INVx1_ASAP7_75t_L g598 ( .A(n_61), .Y(n_598) );
INVx2_ASAP7_75t_L g634 ( .A(n_61), .Y(n_634) );
OR2x2_ASAP7_75t_L g501 ( .A(n_62), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g248 ( .A(n_63), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_64), .B(n_124), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_66), .B(n_172), .Y(n_204) );
INVx1_ASAP7_75t_L g153 ( .A(n_67), .Y(n_153) );
INVx2_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g178 ( .A(n_69), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g506 ( .A(n_70), .Y(n_506) );
INVx1_ASAP7_75t_L g544 ( .A(n_71), .Y(n_544) );
INVx1_ASAP7_75t_L g574 ( .A(n_72), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g559 ( .A1(n_73), .A2(n_560), .B(n_563), .C(n_573), .Y(n_559) );
BUFx3_ASAP7_75t_L g521 ( .A(n_74), .Y(n_521) );
INVx1_ASAP7_75t_L g537 ( .A(n_74), .Y(n_537) );
BUFx3_ASAP7_75t_L g523 ( .A(n_75), .Y(n_523) );
INVx1_ASAP7_75t_L g539 ( .A(n_75), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_76), .B(n_172), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_481), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_SL g127 ( .A(n_82), .Y(n_127) );
INVx8_ASAP7_75t_L g185 ( .A(n_82), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_82), .A2(n_129), .B(n_256), .Y(n_255) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AOI21xp33_ASAP7_75t_L g154 ( .A1(n_83), .A2(n_130), .B(n_152), .Y(n_154) );
INVx1_ASAP7_75t_L g165 ( .A(n_83), .Y(n_165) );
INVx1_ASAP7_75t_L g217 ( .A(n_83), .Y(n_217) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g695 ( .A1(n_86), .A2(n_696), .B(n_697), .Y(n_695) );
NAND2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
INVx2_ASAP7_75t_L g180 ( .A(n_90), .Y(n_180) );
INVx2_ASAP7_75t_L g182 ( .A(n_90), .Y(n_182) );
INVx2_ASAP7_75t_L g184 ( .A(n_90), .Y(n_184) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_91), .Y(n_116) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
INVx2_ASAP7_75t_L g160 ( .A(n_91), .Y(n_160) );
INVx1_ASAP7_75t_L g245 ( .A(n_91), .Y(n_245) );
OAI21xp33_ASAP7_75t_L g157 ( .A1(n_92), .A2(n_158), .B(n_164), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_92), .A2(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g233 ( .A(n_92), .Y(n_233) );
INVx5_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx5_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
BUFx12f_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx3_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
NAND4xp75_ASAP7_75t_L g99 ( .A(n_100), .B(n_340), .C(n_395), .D(n_442), .Y(n_99) );
NOR2x1_ASAP7_75t_L g100 ( .A(n_101), .B(n_290), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_102), .B(n_269), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_189), .B1(n_235), .B2(n_257), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_131), .Y(n_104) );
AND2x2_ASAP7_75t_L g275 ( .A(n_105), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g315 ( .A(n_105), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g329 ( .A(n_105), .B(n_262), .Y(n_329) );
INVx2_ASAP7_75t_L g346 ( .A(n_105), .Y(n_346) );
INVx2_ASAP7_75t_L g406 ( .A(n_105), .Y(n_406) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g260 ( .A(n_106), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g268 ( .A(n_106), .B(n_175), .Y(n_268) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g327 ( .A(n_107), .Y(n_327) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_113), .B(n_128), .Y(n_107) );
OAI21x1_ASAP7_75t_SL g223 ( .A1(n_108), .A2(n_224), .B(n_234), .Y(n_223) );
BUFx4f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_109), .B(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g194 ( .A(n_109), .Y(n_194) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g173 ( .A(n_111), .Y(n_173) );
OAI21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B(n_127), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_117), .B(n_120), .Y(n_114) );
INVx2_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx2_ASAP7_75t_L g228 ( .A(n_116), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_118), .B(n_142), .Y(n_141) );
INVxp67_ASAP7_75t_L g213 ( .A(n_118), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_118), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx2_ASAP7_75t_SL g126 ( .A(n_120), .Y(n_126) );
CKINVDCx6p67_ASAP7_75t_R g200 ( .A(n_120), .Y(n_200) );
INVx2_ASAP7_75t_SL g215 ( .A(n_120), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_126), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_123), .A2(n_147), .B1(n_149), .B2(n_150), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_123), .A2(n_159), .B1(n_209), .B2(n_210), .Y(n_208) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g250 ( .A(n_124), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_130), .B(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_130), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_155), .Y(n_131) );
INVx1_ASAP7_75t_L g277 ( .A(n_132), .Y(n_277) );
INVxp67_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g372 ( .A(n_133), .B(n_261), .Y(n_372) );
AND2x2_ASAP7_75t_L g386 ( .A(n_133), .B(n_156), .Y(n_386) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g263 ( .A(n_134), .B(n_156), .Y(n_263) );
AND2x2_ASAP7_75t_L g359 ( .A(n_134), .B(n_156), .Y(n_359) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g284 ( .A(n_135), .Y(n_284) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_145), .B(n_154), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_143), .Y(n_136) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_140), .A2(n_243), .B1(n_244), .B2(n_246), .Y(n_242) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_144), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_144), .B(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_144), .A2(n_178), .B1(n_181), .B2(n_183), .Y(n_177) );
INVx3_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_151), .B(n_152), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_149), .A2(n_498), .B1(n_499), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_149), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_150), .Y(n_693) );
AO21x1_ASAP7_75t_L g241 ( .A1(n_151), .A2(n_242), .B(n_247), .Y(n_241) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_151), .A2(n_250), .B(n_252), .Y(n_249) );
AND2x2_ASAP7_75t_L g276 ( .A(n_155), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g316 ( .A(n_155), .Y(n_316) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_174), .Y(n_155) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_156), .Y(n_266) );
INVx2_ASAP7_75t_SL g301 ( .A(n_156), .Y(n_301) );
INVx1_ASAP7_75t_L g310 ( .A(n_156), .Y(n_310) );
AND2x2_ASAP7_75t_L g471 ( .A(n_156), .B(n_327), .Y(n_471) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_166), .B(n_171), .Y(n_156) );
OAI22xp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B1(n_162), .B2(n_163), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
INVx2_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_162), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g176 ( .A(n_172), .Y(n_176) );
NOR2x1p5_ASAP7_75t_SL g216 ( .A(n_172), .B(n_217), .Y(n_216) );
BUFx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVx1_ASAP7_75t_L g344 ( .A(n_174), .Y(n_344) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g261 ( .A(n_175), .Y(n_261) );
AND2x2_ASAP7_75t_L g309 ( .A(n_175), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_175), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g399 ( .A(n_175), .Y(n_399) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .A3(n_185), .B(n_186), .Y(n_175) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_185), .A2(n_196), .B(n_201), .Y(n_195) );
OAI21x1_ASAP7_75t_SL g224 ( .A1(n_185), .A2(n_225), .B(n_230), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_218), .Y(n_189) );
OR2x2_ASAP7_75t_L g477 ( .A(n_190), .B(n_438), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_205), .Y(n_190) );
INVx2_ASAP7_75t_L g236 ( .A(n_191), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_191), .B(n_222), .Y(n_307) );
AND2x2_ASAP7_75t_L g331 ( .A(n_191), .B(n_274), .Y(n_331) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g272 ( .A(n_192), .Y(n_272) );
OAI21x1_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_195), .B(n_204), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_199), .B(n_200), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_200), .A2(n_208), .B(n_211), .C(n_216), .Y(n_207) );
INVx1_ASAP7_75t_L g221 ( .A(n_205), .Y(n_221) );
INVx1_ASAP7_75t_L g238 ( .A(n_205), .Y(n_238) );
INVx2_ASAP7_75t_L g296 ( .A(n_205), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_205), .B(n_239), .Y(n_305) );
AND2x2_ASAP7_75t_L g337 ( .A(n_205), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g349 ( .A(n_205), .B(n_222), .Y(n_349) );
INVx1_ASAP7_75t_L g427 ( .A(n_205), .Y(n_427) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .C(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g279 ( .A(n_220), .Y(n_279) );
AND2x2_ASAP7_75t_L g373 ( .A(n_220), .B(n_287), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_220), .B(n_354), .Y(n_375) );
AND2x4_ASAP7_75t_L g434 ( .A(n_220), .B(n_389), .Y(n_434) );
AND2x4_ASAP7_75t_L g449 ( .A(n_220), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g421 ( .A(n_222), .Y(n_421) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx3_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_229), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x2_ASAP7_75t_L g366 ( .A(n_236), .B(n_304), .Y(n_366) );
INVx1_ASAP7_75t_L g401 ( .A(n_236), .Y(n_401) );
INVx2_ASAP7_75t_L g450 ( .A(n_236), .Y(n_450) );
AND2x2_ASAP7_75t_L g468 ( .A(n_236), .B(n_349), .Y(n_468) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_237), .Y(n_352) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g364 ( .A(n_239), .Y(n_364) );
AND2x2_ASAP7_75t_L g392 ( .A(n_239), .B(n_274), .Y(n_392) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
INVx1_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_249), .B(n_255), .Y(n_240) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g256 ( .A(n_247), .Y(n_256) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_264), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_260), .B(n_300), .Y(n_367) );
AND2x4_ASAP7_75t_L g417 ( .A(n_262), .B(n_268), .Y(n_417) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g403 ( .A(n_263), .B(n_287), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_263), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g472 ( .A1(n_264), .A2(n_473), .B1(n_475), .B2(n_477), .C1(n_478), .C2(n_480), .Y(n_472) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g324 ( .A(n_266), .Y(n_324) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_268), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
AND2x2_ASAP7_75t_L g334 ( .A(n_268), .B(n_324), .Y(n_334) );
AND2x2_ASAP7_75t_L g385 ( .A(n_268), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g423 ( .A(n_268), .B(n_358), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_275), .B(n_278), .C(n_285), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
AND2x4_ASAP7_75t_L g322 ( .A(n_271), .B(n_274), .Y(n_322) );
BUFx2_ASAP7_75t_L g389 ( .A(n_271), .Y(n_389) );
AND2x2_ASAP7_75t_L g414 ( .A(n_271), .B(n_296), .Y(n_414) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g354 ( .A(n_272), .B(n_289), .Y(n_354) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g295 ( .A(n_274), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g413 ( .A(n_274), .Y(n_413) );
INVx2_ASAP7_75t_SL g441 ( .A(n_276), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_282), .B(n_326), .Y(n_452) );
AND2x2_ASAP7_75t_L g461 ( .A(n_282), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g343 ( .A(n_283), .B(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_283), .B(n_344), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_283), .B(n_327), .Y(n_458) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g466 ( .A(n_284), .B(n_327), .Y(n_466) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g294 ( .A(n_287), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g379 ( .A(n_287), .B(n_365), .Y(n_379) );
AND2x2_ASAP7_75t_L g433 ( .A(n_287), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g440 ( .A(n_287), .B(n_322), .Y(n_440) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_317), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_297), .B1(n_302), .B2(n_308), .C(n_311), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g312 ( .A(n_295), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g454 ( .A(n_295), .Y(n_454) );
INVx1_ASAP7_75t_L g390 ( .A(n_296), .Y(n_390) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_299), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_350) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g345 ( .A(n_300), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_327), .Y(n_371) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_304), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g465 ( .A(n_309), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g462 ( .A(n_310), .B(n_399), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_313), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_315), .A2(n_333), .B(n_335), .Y(n_332) );
OR2x2_ASAP7_75t_L g376 ( .A(n_316), .B(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_332), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B1(n_328), .B2(n_330), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g336 ( .A(n_322), .B(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_322), .A2(n_329), .B1(n_370), .B2(n_373), .C(n_374), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_322), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g408 ( .A(n_326), .B(n_359), .Y(n_408) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
INVx1_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_331), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g424 ( .A(n_331), .Y(n_424) );
AND2x2_ASAP7_75t_L g437 ( .A(n_331), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
INVx2_ASAP7_75t_L g438 ( .A(n_338), .Y(n_438) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_339), .Y(n_411) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_368), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_342), .B(n_360), .Y(n_341) );
O2A1O1Ixp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B(n_347), .C(n_350), .Y(n_342) );
AND2x2_ASAP7_75t_L g429 ( .A(n_346), .B(n_386), .Y(n_429) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_346), .Y(n_446) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g365 ( .A(n_349), .Y(n_365) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g432 ( .A(n_358), .Y(n_432) );
BUFx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_359), .B(n_377), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_366), .B(n_367), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_361), .A2(n_405), .B1(n_408), .B2(n_409), .Y(n_404) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g469 ( .A(n_363), .Y(n_469) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_364), .B(n_421), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_381), .Y(n_368) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_371), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_372), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g474 ( .A(n_372), .B(n_377), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_372), .B(n_471), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_379), .B2(n_380), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OA22x2_ASAP7_75t_L g451 ( .A1(n_379), .A2(n_452), .B1(n_453), .B2(n_456), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_387), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_391), .B(n_393), .Y(n_387) );
NAND2xp33_ASAP7_75t_SL g418 ( .A(n_388), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_396), .B(n_415), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B(n_404), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_403), .A2(n_445), .B(n_447), .Y(n_444) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AND2x2_ASAP7_75t_L g431 ( .A(n_406), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g447 ( .A(n_408), .Y(n_447) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g422 ( .A(n_410), .Y(n_422) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_430), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_423), .B2(n_424), .C1(n_425), .C2(n_429), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_426), .A2(n_460), .B1(n_463), .B2(n_464), .C(n_467), .Y(n_459) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_428), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_435), .Y(n_430) );
AOI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_439), .B(n_441), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g455 ( .A(n_438), .Y(n_455) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR3x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_459), .C(n_472), .Y(n_442) );
OAI21x1_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_448), .B(n_451), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g479 ( .A(n_454), .Y(n_479) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_663), .B1(n_681), .B2(n_683), .C(n_686), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_498), .B1(n_499), .B2(n_662), .Y(n_482) );
INVx1_ASAP7_75t_L g662 ( .A(n_483), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_492), .B2(n_493), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
XOR2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_496), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g500 ( .A(n_501), .B(n_524), .C(n_592), .D(n_647), .Y(n_500) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_508), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_L g603 ( .A(n_506), .B(n_507), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_506), .Y(n_607) );
INVx2_ASAP7_75t_L g613 ( .A(n_506), .Y(n_613) );
AND2x4_ASAP7_75t_L g620 ( .A(n_506), .B(n_608), .Y(n_620) );
INVx1_ASAP7_75t_L g644 ( .A(n_506), .Y(n_644) );
INVx2_ASAP7_75t_L g608 ( .A(n_507), .Y(n_608) );
INVx1_ASAP7_75t_L g615 ( .A(n_507), .Y(n_615) );
INVx1_ASAP7_75t_L g639 ( .A(n_507), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_508), .Y(n_640) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
BUFx2_ASAP7_75t_L g558 ( .A(n_514), .Y(n_558) );
AND2x4_ASAP7_75t_L g565 ( .A(n_514), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g570 ( .A(n_514), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g680 ( .A(n_514), .B(n_566), .Y(n_680) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g582 ( .A(n_517), .B(n_555), .Y(n_582) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g554 ( .A(n_518), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g580 ( .A(n_519), .Y(n_580) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g529 ( .A(n_521), .B(n_523), .Y(n_529) );
AND2x4_ASAP7_75t_L g552 ( .A(n_521), .B(n_539), .Y(n_552) );
INVx1_ASAP7_75t_L g568 ( .A(n_522), .Y(n_568) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g543 ( .A(n_523), .B(n_537), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_559), .A3(n_583), .B(n_587), .Y(n_524) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
AND2x4_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g561 ( .A(n_530), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g584 ( .A(n_531), .B(n_535), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_531), .B(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_540), .B1(n_541), .B2(n_544), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g549 ( .A(n_536), .B(n_538), .Y(n_549) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g586 ( .A(n_543), .Y(n_586) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_550), .Y(n_545) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g575 ( .A(n_548), .Y(n_575) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_552), .Y(n_562) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_552), .Y(n_577) );
BUFx2_ASAP7_75t_L g672 ( .A(n_553), .Y(n_672) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_569), .B2(n_570), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_564), .A2(n_569), .B1(n_637), .B2(n_641), .C(n_645), .Y(n_636) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g675 ( .A(n_567), .Y(n_675) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_576), .C(n_578), .Y(n_573) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g594 ( .A(n_590), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g630 ( .A(n_590), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_593), .B(n_636), .Y(n_592) );
AOI33xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_599), .A3(n_609), .B1(n_621), .B2(n_626), .B3(n_630), .Y(n_593) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g648 ( .A(n_601), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_603), .Y(n_629) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g646 ( .A(n_606), .Y(n_646) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_606), .Y(n_661) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_612), .Y(n_654) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g658 ( .A(n_618), .B(n_649), .Y(n_658) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g625 ( .A(n_620), .Y(n_625) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_L g641 ( .A(n_640), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g645 ( .A(n_640), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_652), .B1(n_653), .B2(n_655), .C(n_656), .Y(n_647) );
AND2x2_ASAP7_75t_L g653 ( .A(n_649), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g660 ( .A(n_649), .B(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x6_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
OR2x4_ASAP7_75t_L g690 ( .A(n_667), .B(n_671), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_668), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g696 ( .A(n_668), .Y(n_696) );
INVx1_ASAP7_75t_L g685 ( .A(n_669), .Y(n_685) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI31xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .A3(n_676), .B(n_678), .Y(n_671) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx6_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_691), .B1(n_693), .B2(n_694), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx8_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
endmodule