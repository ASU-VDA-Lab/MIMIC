module real_aes_6543_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g172 ( .A1(n_0), .A2(n_173), .B(n_174), .C(n_178), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_1), .B(n_167), .Y(n_180) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_3), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_4), .A2(n_161), .B(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_5), .A2(n_141), .B(n_158), .C(n_510), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_6), .A2(n_161), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_7), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_8), .B(n_167), .Y(n_472) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_9), .A2(n_133), .B(n_255), .Y(n_254) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_10), .A2(n_442), .B1(n_712), .B2(n_715), .C1(n_719), .C2(n_720), .Y(n_441) );
AND2x6_ASAP7_75t_L g158 ( .A(n_11), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_12), .A2(n_141), .B(n_158), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g563 ( .A(n_13), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_14), .B(n_41), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_15), .B(n_177), .Y(n_512) );
INVx1_ASAP7_75t_L g138 ( .A(n_16), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_17), .B(n_152), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_18), .A2(n_153), .B(n_521), .C(n_523), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_19), .B(n_167), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_20), .B(n_195), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_21), .A2(n_141), .B(n_187), .C(n_194), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_22), .A2(n_176), .B(n_229), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_23), .B(n_177), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_24), .B(n_177), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_25), .Y(n_490) );
INVx1_ASAP7_75t_L g460 ( .A(n_26), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_27), .A2(n_141), .B(n_194), .C(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_28), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_29), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_30), .A2(n_102), .B1(n_115), .B2(n_725), .Y(n_101) );
INVx1_ASAP7_75t_L g484 ( .A(n_31), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_32), .A2(n_161), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_34), .A2(n_156), .B(n_210), .C(n_211), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_35), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_36), .A2(n_176), .B(n_469), .C(n_471), .Y(n_468) );
INVxp67_ASAP7_75t_L g485 ( .A(n_37), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_38), .B(n_260), .Y(n_259) );
CKINVDCx14_ASAP7_75t_R g467 ( .A(n_39), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_40), .A2(n_141), .B(n_194), .C(n_459), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_42), .A2(n_178), .B(n_561), .C(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_43), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_44), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_45), .B(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_46), .B(n_161), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_47), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_48), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_49), .A2(n_156), .B(n_210), .C(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g175 ( .A(n_50), .Y(n_175) );
INVx1_ASAP7_75t_L g239 ( .A(n_51), .Y(n_239) );
INVx1_ASAP7_75t_L g528 ( .A(n_52), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_53), .B(n_161), .Y(n_236) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_54), .A2(n_71), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_54), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_55), .Y(n_199) );
CKINVDCx14_ASAP7_75t_R g559 ( .A(n_56), .Y(n_559) );
INVx1_ASAP7_75t_L g159 ( .A(n_57), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_58), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_59), .B(n_167), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_60), .A2(n_148), .B(n_193), .C(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_61), .A2(n_70), .B1(n_713), .B2(n_714), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_61), .Y(n_713) );
INVx1_ASAP7_75t_L g137 ( .A(n_62), .Y(n_137) );
INVx1_ASAP7_75t_SL g470 ( .A(n_63), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_65), .B(n_152), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_66), .B(n_167), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_67), .B(n_153), .Y(n_226) );
INVx1_ASAP7_75t_L g493 ( .A(n_68), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_69), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_70), .Y(n_714) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_72), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_73), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_74), .Y(n_248) );
INVx1_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_76), .A2(n_161), .B(n_558), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_77), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_78), .A2(n_161), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_79), .A2(n_185), .B(n_480), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_80), .Y(n_457) );
INVx1_ASAP7_75t_L g519 ( .A(n_81), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_82), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_83), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_84), .A2(n_161), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g522 ( .A(n_85), .Y(n_522) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g511 ( .A(n_87), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_88), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_89), .B(n_177), .Y(n_227) );
OR2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g446 ( .A(n_90), .B(n_112), .Y(n_446) );
INVx2_ASAP7_75t_L g711 ( .A(n_90), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_91), .A2(n_141), .B(n_156), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_92), .B(n_161), .Y(n_208) );
INVx1_ASAP7_75t_L g212 ( .A(n_93), .Y(n_212) );
INVxp67_ASAP7_75t_L g251 ( .A(n_94), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_95), .B(n_133), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
INVx1_ASAP7_75t_L g222 ( .A(n_98), .Y(n_222) );
INVx2_ASAP7_75t_L g531 ( .A(n_99), .Y(n_531) );
AND2x2_ASAP7_75t_L g241 ( .A(n_100), .B(n_197), .Y(n_241) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g726 ( .A(n_105), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g436 ( .A(n_110), .Y(n_436) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_110), .Y(n_439) );
NOR2x2_ASAP7_75t_L g722 ( .A(n_111), .B(n_711), .Y(n_722) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g710 ( .A(n_112), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_440), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g724 ( .A(n_119), .Y(n_724) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_436), .B(n_437), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_L g443 ( .A(n_126), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_126), .A2(n_448), .B1(n_716), .B2(n_717), .Y(n_715) );
OR3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_344), .C(n_393), .Y(n_126) );
NAND5xp2_ASAP7_75t_L g127 ( .A(n_128), .B(n_278), .C(n_307), .D(n_315), .E(n_330), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_201), .B(n_217), .C(n_262), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_181), .Y(n_129) );
AND2x2_ASAP7_75t_L g273 ( .A(n_130), .B(n_270), .Y(n_273) );
AND2x2_ASAP7_75t_L g306 ( .A(n_130), .B(n_182), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_130), .B(n_205), .Y(n_399) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
INVx2_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
BUFx2_ASAP7_75t_L g373 ( .A(n_131), .Y(n_373) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_164), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_132), .B(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_132), .B(n_216), .Y(n_215) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_132), .A2(n_221), .B(n_231), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_132), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_132), .A2(n_489), .B(n_496), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_132), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_133), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_133), .A2(n_256), .B(n_257), .Y(n_255) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g233 ( .A(n_134), .Y(n_233) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_135), .B(n_136), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_160), .Y(n_139) );
INVx5_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
BUFx3_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx1_ASAP7_75t_L g230 ( .A(n_143), .Y(n_230) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_145), .B(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
INVx1_ASAP7_75t_L g260 ( .A(n_145), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_149), .A2(n_152), .B1(n_484), .B2(n_485), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_149), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_149), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
INVx2_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_152), .B(n_251), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_152), .A2(n_192), .B(n_460), .C(n_461), .Y(n_459) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_153), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g471 ( .A(n_155), .Y(n_471) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_157), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_157), .A2(n_171), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_157), .A2(n_171), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_157), .A2(n_171), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_157), .A2(n_171), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_157), .A2(n_171), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g558 ( .A1(n_157), .A2(n_171), .B(n_559), .C(n_560), .Y(n_558) );
INVx4_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g161 ( .A(n_158), .B(n_162), .Y(n_161) );
BUFx3_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_158), .B(n_162), .Y(n_223) );
BUFx2_ASAP7_75t_L g185 ( .A(n_161), .Y(n_185) );
INVx1_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
AND2x2_ASAP7_75t_L g181 ( .A(n_166), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g271 ( .A(n_166), .Y(n_271) );
AND2x2_ASAP7_75t_L g357 ( .A(n_166), .B(n_270), .Y(n_357) );
AND2x2_ASAP7_75t_L g412 ( .A(n_166), .B(n_204), .Y(n_412) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_180), .Y(n_166) );
INVx2_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_176), .B(n_470), .Y(n_469) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g561 ( .A(n_177), .Y(n_561) );
INVx2_ASAP7_75t_L g495 ( .A(n_178), .Y(n_495) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_179), .Y(n_214) );
INVx1_ASAP7_75t_L g523 ( .A(n_179), .Y(n_523) );
INVx1_ASAP7_75t_L g329 ( .A(n_181), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_181), .B(n_205), .Y(n_376) );
INVx5_ASAP7_75t_L g270 ( .A(n_182), .Y(n_270) );
AND2x4_ASAP7_75t_L g291 ( .A(n_182), .B(n_271), .Y(n_291) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_182), .Y(n_313) );
AND2x2_ASAP7_75t_L g388 ( .A(n_182), .B(n_373), .Y(n_388) );
AND2x2_ASAP7_75t_L g391 ( .A(n_182), .B(n_206), .Y(n_391) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
AOI21xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_186), .B(n_195), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_192), .Y(n_187) );
INVx2_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_191), .A2(n_212), .B(n_213), .C(n_214), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_191), .A2(n_214), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_191), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_L g510 ( .A1(n_191), .A2(n_495), .B(n_511), .C(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_193), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_196), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g200 ( .A(n_197), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_197), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_236), .B(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_197), .A2(n_223), .B(n_457), .C(n_458), .Y(n_456) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_197), .A2(n_557), .B(n_564), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_200), .A2(n_507), .B(n_513), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_201), .B(n_271), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_201), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_205), .Y(n_202) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_271), .Y(n_296) );
AND2x2_ASAP7_75t_L g314 ( .A(n_203), .B(n_206), .Y(n_314) );
INVx1_ASAP7_75t_L g334 ( .A(n_203), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_203), .B(n_270), .Y(n_379) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_203), .Y(n_421) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_204), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_205), .B(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_205), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_205), .A2(n_266), .B(n_327), .C(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g333 ( .A(n_205), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g342 ( .A(n_205), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g346 ( .A(n_205), .B(n_270), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_205), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_205), .B(n_271), .Y(n_361) );
AND2x2_ASAP7_75t_L g411 ( .A(n_205), .B(n_412), .Y(n_411) );
INVx5_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
AND2x2_ASAP7_75t_L g316 ( .A(n_206), .B(n_269), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_206), .B(n_303), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_206), .B(n_357), .Y(n_375) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_242), .Y(n_217) );
INVx1_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_234), .Y(n_218) );
OR2x2_ASAP7_75t_L g266 ( .A(n_219), .B(n_234), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_219), .B(n_273), .C(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_219), .B(n_244), .Y(n_283) );
OR2x2_ASAP7_75t_L g298 ( .A(n_219), .B(n_286), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_219), .B(n_253), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_219), .B(n_435), .Y(n_434) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_220), .B(n_244), .Y(n_301) );
AND2x2_ASAP7_75t_L g340 ( .A(n_220), .B(n_254), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_220), .B(n_253), .Y(n_368) );
OR2x2_ASAP7_75t_L g371 ( .A(n_220), .B(n_253), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_223), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_223), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_259), .B(n_261), .Y(n_258) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g478 ( .A(n_233), .Y(n_478) );
INVx5_ASAP7_75t_SL g286 ( .A(n_234), .Y(n_286) );
OR2x2_ASAP7_75t_L g292 ( .A(n_234), .B(n_243), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_234), .B(n_309), .Y(n_308) );
AOI321xp33_ASAP7_75t_L g315 ( .A1(n_234), .A2(n_316), .A3(n_317), .B1(n_318), .B2(n_324), .C(n_326), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_234), .B(n_242), .Y(n_325) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_234), .Y(n_338) );
OR2x2_ASAP7_75t_L g385 ( .A(n_234), .B(n_283), .Y(n_385) );
AND2x2_ASAP7_75t_L g407 ( .A(n_234), .B(n_304), .Y(n_407) );
AND2x2_ASAP7_75t_L g426 ( .A(n_234), .B(n_244), .Y(n_426) );
OR2x6_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_244), .B(n_253), .Y(n_267) );
AND2x2_ASAP7_75t_L g276 ( .A(n_244), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g303 ( .A(n_244), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_244), .B(n_304), .Y(n_309) );
INVxp67_ASAP7_75t_L g339 ( .A(n_244), .Y(n_339) );
OR2x2_ASAP7_75t_L g381 ( .A(n_244), .B(n_286), .Y(n_381) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_252), .Y(n_244) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_245), .A2(n_465), .B(n_472), .Y(n_464) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_245), .A2(n_517), .B(n_524), .Y(n_516) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_245), .A2(n_526), .B(n_532), .Y(n_525) );
OR2x2_ASAP7_75t_L g263 ( .A(n_253), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g277 ( .A(n_253), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_253), .B(n_266), .Y(n_310) );
AND2x2_ASAP7_75t_L g359 ( .A(n_253), .B(n_303), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_253), .B(n_286), .Y(n_397) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_254), .B(n_286), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_268), .C(n_272), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_263), .A2(n_265), .B1(n_390), .B2(n_392), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_265), .A2(n_288), .B1(n_343), .B2(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_SL g417 ( .A(n_266), .Y(n_417) );
INVx1_ASAP7_75t_SL g317 ( .A(n_267), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_269), .B(n_289), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g330 ( .A1(n_269), .A2(n_310), .B1(n_317), .B2(n_331), .C1(n_335), .C2(n_341), .Y(n_330) );
AND2x2_ASAP7_75t_L g420 ( .A(n_269), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_270), .B(n_290), .Y(n_365) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_270), .Y(n_402) );
AND2x2_ASAP7_75t_L g405 ( .A(n_270), .B(n_314), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_270), .B(n_421), .Y(n_431) );
INVx1_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_273), .A2(n_414), .B(n_415), .C(n_418), .Y(n_413) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_275), .B(n_337), .C(n_340), .Y(n_336) );
OR2x2_ASAP7_75t_L g364 ( .A(n_275), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_275), .B(n_291), .Y(n_392) );
OR2x2_ASAP7_75t_L g297 ( .A(n_277), .B(n_298), .Y(n_297) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .B(n_287), .C(n_299), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_280), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g386 ( .A(n_281), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_282), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g300 ( .A(n_285), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_286), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g354 ( .A(n_286), .B(n_304), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_286), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_286), .B(n_303), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B1(n_293), .B2(n_297), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_289), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_291), .B(n_333), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_292), .A2(n_356), .B1(n_358), .B2(n_360), .C(n_362), .Y(n_355) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g410 ( .A(n_295), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g423 ( .A(n_295), .B(n_412), .Y(n_423) );
INVx1_ASAP7_75t_L g343 ( .A(n_296), .Y(n_343) );
INVx1_ASAP7_75t_L g414 ( .A(n_297), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_298), .A2(n_381), .B(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_302), .B(n_305), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_310), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g347 ( .A(n_308), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_309), .A2(n_395), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_394) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_317), .A2(n_407), .B1(n_408), .B2(n_410), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp67_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g387 ( .A(n_323), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_333), .B(n_357), .Y(n_409) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_339), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g425 ( .A(n_340), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_340), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI211xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_347), .B(n_348), .C(n_382), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_355), .C(n_374), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g435 ( .A(n_359), .Y(n_435) );
AND2x2_ASAP7_75t_L g372 ( .A(n_361), .B(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_370), .B2(n_372), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g380 ( .A(n_368), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI31xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .A3(n_377), .B(n_380), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .C(n_389), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g390 ( .A(n_391), .Y(n_390) );
NAND5xp2_ASAP7_75t_L g393 ( .A(n_394), .B(n_406), .C(n_413), .D(n_427), .E(n_430), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_405), .A2(n_431), .B1(n_432), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_SL g429 ( .A(n_407), .Y(n_429) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_424), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_437), .B(n_441), .C(n_723), .Y(n_440) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_710), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g716 ( .A(n_445), .Y(n_716) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR3x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_621), .C(n_668), .Y(n_448) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_567), .C(n_592), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_505), .B1(n_533), .B2(n_536), .C(n_544), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_473), .B(n_498), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_453), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_453), .B(n_549), .Y(n_665) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_464), .Y(n_453) );
AND2x2_ASAP7_75t_L g535 ( .A(n_454), .B(n_504), .Y(n_535) );
AND2x2_ASAP7_75t_L g585 ( .A(n_454), .B(n_503), .Y(n_585) );
AND2x2_ASAP7_75t_L g606 ( .A(n_454), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_454), .B(n_578), .Y(n_611) );
OR2x2_ASAP7_75t_L g619 ( .A(n_454), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g691 ( .A(n_454), .B(n_487), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_454), .B(n_640), .Y(n_705) );
INVx3_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g550 ( .A(n_455), .B(n_464), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_455), .B(n_487), .Y(n_551) );
AND2x4_ASAP7_75t_L g573 ( .A(n_455), .B(n_504), .Y(n_573) );
AND2x2_ASAP7_75t_L g603 ( .A(n_455), .B(n_475), .Y(n_603) );
AND2x2_ASAP7_75t_L g612 ( .A(n_455), .B(n_602), .Y(n_612) );
AND2x2_ASAP7_75t_L g628 ( .A(n_455), .B(n_488), .Y(n_628) );
OR2x2_ASAP7_75t_L g637 ( .A(n_455), .B(n_620), .Y(n_637) );
AND2x2_ASAP7_75t_L g643 ( .A(n_455), .B(n_578), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_455), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g657 ( .A(n_455), .B(n_500), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_455), .B(n_546), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_455), .B(n_607), .Y(n_696) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_462), .Y(n_455) );
INVx2_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
AND2x2_ASAP7_75t_L g602 ( .A(n_464), .B(n_487), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_464), .B(n_488), .Y(n_607) );
INVx1_ASAP7_75t_L g663 ( .A(n_464), .Y(n_663) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g572 ( .A(n_474), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_487), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_475), .B(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
OR2x2_ASAP7_75t_L g620 ( .A(n_475), .B(n_487), .Y(n_620) );
OR2x2_ASAP7_75t_L g681 ( .A(n_475), .B(n_588), .Y(n_681) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_486), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_477), .A2(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g501 ( .A(n_479), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_486), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_487), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g640 ( .A(n_487), .B(n_500), .Y(n_640) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g579 ( .A(n_488), .Y(n_579) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_499), .A2(n_685), .B1(n_689), .B2(n_692), .C(n_693), .Y(n_684) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_SL g547 ( .A(n_500), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_500), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g679 ( .A(n_500), .B(n_535), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_503), .B(n_549), .Y(n_671) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g582 ( .A(n_505), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_505), .B(n_588), .Y(n_618) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
AND2x2_ASAP7_75t_L g543 ( .A(n_506), .B(n_516), .Y(n_543) );
INVx4_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
BUFx3_ASAP7_75t_L g598 ( .A(n_506), .Y(n_598) );
AND3x2_ASAP7_75t_L g613 ( .A(n_506), .B(n_614), .C(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g695 ( .A(n_515), .B(n_609), .Y(n_695) );
AND2x2_ASAP7_75t_L g703 ( .A(n_515), .B(n_588), .Y(n_703) );
INVx1_ASAP7_75t_SL g708 ( .A(n_515), .Y(n_708) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
INVx1_ASAP7_75t_SL g566 ( .A(n_516), .Y(n_566) );
AND2x2_ASAP7_75t_L g589 ( .A(n_516), .B(n_555), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_516), .B(n_539), .Y(n_591) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_516), .Y(n_631) );
OR2x2_ASAP7_75t_L g636 ( .A(n_516), .B(n_555), .Y(n_636) );
INVx2_ASAP7_75t_L g541 ( .A(n_525), .Y(n_541) );
AND2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_556), .Y(n_576) );
OR2x2_ASAP7_75t_L g596 ( .A(n_525), .B(n_556), .Y(n_596) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_525), .Y(n_616) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_534), .A2(n_575), .B(n_667), .Y(n_666) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_536), .A2(n_546), .A3(n_573), .B1(n_703), .B2(n_704), .C1(n_706), .C2(n_709), .Y(n_702) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_538), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_539), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g565 ( .A(n_540), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g633 ( .A(n_541), .B(n_555), .Y(n_633) );
AND2x2_ASAP7_75t_L g700 ( .A(n_541), .B(n_556), .Y(n_700) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g641 ( .A(n_543), .B(n_595), .Y(n_641) );
AOI31xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .A3(n_551), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g600 ( .A(n_546), .B(n_578), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_546), .B(n_570), .Y(n_682) );
AND2x2_ASAP7_75t_L g701 ( .A(n_546), .B(n_606), .Y(n_701) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_549), .B(n_578), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_549), .B(n_607), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_549), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_549), .B(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_550), .B(n_607), .Y(n_639) );
INVx1_ASAP7_75t_L g683 ( .A(n_550), .Y(n_683) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_565), .Y(n_553) );
INVxp67_ASAP7_75t_L g635 ( .A(n_554), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_555), .B(n_566), .Y(n_571) );
INVx1_ASAP7_75t_L g677 ( .A(n_555), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_555), .B(n_654), .Y(n_688) );
BUFx3_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_556), .B(n_566), .Y(n_614) );
INVx2_ASAP7_75t_L g654 ( .A(n_556), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_565), .B(n_687), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .B(n_574), .C(n_583), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_569), .A2(n_618), .B(n_619), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_570), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_570), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g650 ( .A(n_571), .B(n_596), .Y(n_650) );
INVx3_ASAP7_75t_L g581 ( .A(n_573), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_577), .B1(n_580), .B2(n_582), .Y(n_574) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_576), .A2(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g625 ( .A(n_576), .B(n_589), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_576), .B(n_677), .Y(n_676) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g580 ( .A(n_579), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g649 ( .A(n_579), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_580), .A2(n_594), .B(n_599), .Y(n_593) );
OAI22xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_586), .B1(n_590), .B2(n_591), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_585), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_588), .B(n_631), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_604), .C(n_617), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_594), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g664 ( .A(n_596), .B(n_597), .Y(n_664) );
AND2x2_ASAP7_75t_L g672 ( .A(n_597), .B(n_653), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_598), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_SL g680 ( .A1(n_598), .A2(n_681), .B(n_682), .C(n_683), .Y(n_680) );
OR2x2_ASAP7_75t_L g707 ( .A(n_598), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B(n_610), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_606), .A2(n_643), .B(n_644), .C(n_647), .Y(n_642) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B(n_613), .Y(n_610) );
AND2x2_ASAP7_75t_L g675 ( .A(n_614), .B(n_633), .Y(n_675) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g653 ( .A(n_616), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_618), .Y(n_658) );
NAND3xp33_ASAP7_75t_SL g621 ( .A(n_622), .B(n_642), .C(n_655), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B(n_626), .C(n_634), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g692 ( .A(n_629), .Y(n_692) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g652 ( .A(n_631), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_631), .B(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_637), .C(n_638), .Y(n_634) );
INVx2_ASAP7_75t_SL g646 ( .A(n_636), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_637), .A2(n_648), .B1(n_650), .B2(n_651), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_640), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B(n_659), .C(n_666), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVxp33_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g709 ( .A(n_663), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_669), .B(n_684), .C(n_697), .D(n_702), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_673), .C(n_680), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_678), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_674), .A2(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_681), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g718 ( .A(n_710), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_712), .Y(n_719) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx3_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
endmodule