module fake_ibex_1941_n_3658 (n_151, n_85, n_599, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3658);

input n_151;
input n_85;
input n_599;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3658;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_2230;
wire n_1782;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2333;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3023;
wire n_784;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2451;
wire n_2166;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_3241;
wire n_1121;
wire n_2746;
wire n_2397;
wire n_2256;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2697;
wire n_2224;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_3416;
wire n_1031;
wire n_2962;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2971;
wire n_3578;
wire n_954;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2612;
wire n_2193;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_2263;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2923;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_3284;
wire n_2524;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_3314;
wire n_2997;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_3556;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2698;
wire n_2274;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_3162;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_2154;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1542;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2494;
wire n_2156;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3163;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2652;
wire n_2227;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_3015;
wire n_2588;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2303;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g778 ( 
.A(n_370),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_552),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_775),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_576),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_51),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_287),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_735),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_331),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_238),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_708),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_58),
.Y(n_789)
);

BUFx2_ASAP7_75t_SL g790 ( 
.A(n_604),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_444),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_206),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_668),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_670),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_668),
.Y(n_795)
);

BUFx10_ASAP7_75t_L g796 ( 
.A(n_559),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_257),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_571),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_572),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_695),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_428),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_411),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_77),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_129),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_301),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_757),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_452),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_691),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_677),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_154),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_198),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_429),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_720),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_472),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_167),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_667),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_453),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_584),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_553),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_506),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_299),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_638),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_350),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_463),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_698),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_524),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_625),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_688),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_418),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_769),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_542),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_582),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_686),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_103),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_509),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_375),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_269),
.B(n_436),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_769),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_89),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_37),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_433),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_605),
.Y(n_843)
);

INVxp33_ASAP7_75t_R g844 ( 
.A(n_131),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_181),
.B(n_26),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_9),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_647),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_134),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_341),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_295),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_154),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_65),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_170),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_594),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_1),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_383),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_521),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_168),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_321),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_748),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_592),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_31),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_726),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_463),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_564),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_605),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_680),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_152),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_109),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_404),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_599),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_701),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_29),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_610),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_699),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_473),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_276),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_3),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_651),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_202),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_481),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_709),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_632),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_223),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_598),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_393),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_247),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_301),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_214),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_502),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_704),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_69),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_645),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_590),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_190),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_380),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_4),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_761),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_700),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_80),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_216),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_717),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_426),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_7),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_103),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_127),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_643),
.B(n_727),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_537),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_454),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_109),
.Y(n_910)
);

CKINVDCx14_ASAP7_75t_R g911 ( 
.A(n_369),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_512),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_201),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_373),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_496),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_455),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_760),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_229),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_584),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_306),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_701),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_604),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_749),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_521),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_163),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_386),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_78),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_445),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_452),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_207),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_277),
.Y(n_931)
);

BUFx8_ASAP7_75t_SL g932 ( 
.A(n_149),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_618),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_397),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_69),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_160),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_299),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_143),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_149),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_203),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_210),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_316),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_139),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_65),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_308),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_586),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_229),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_18),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_615),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_66),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_483),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_763),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_618),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_120),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_436),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_183),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_88),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_324),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_440),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_242),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_690),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_26),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_30),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_706),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_703),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_581),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_36),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_35),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_569),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_734),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_340),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_466),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_695),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_471),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_96),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_338),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_585),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_544),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_126),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_251),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_507),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_758),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_415),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_368),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_615),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_430),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_776),
.Y(n_987)
);

BUFx10_ASAP7_75t_L g988 ( 
.A(n_80),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_220),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_68),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_433),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_302),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_582),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_602),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_217),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_472),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_603),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_157),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_663),
.Y(n_999)
);

CKINVDCx16_ASAP7_75t_R g1000 ( 
.A(n_542),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_438),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_644),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_451),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_319),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_683),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_706),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_626),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_408),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_234),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_365),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_563),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_166),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_354),
.Y(n_1013)
);

CKINVDCx11_ASAP7_75t_R g1014 ( 
.A(n_176),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_455),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_458),
.Y(n_1016)
);

XOR2xp5_ASAP7_75t_R g1017 ( 
.A(n_273),
.B(n_379),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_570),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_63),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_768),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_523),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_638),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_266),
.Y(n_1023)
);

BUFx5_ASAP7_75t_L g1024 ( 
.A(n_435),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_628),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_457),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_226),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_760),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_546),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_418),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_745),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_313),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_540),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_38),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_748),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_624),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_612),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_555),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_134),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_353),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_485),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_653),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_33),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_113),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_344),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_774),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_205),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_525),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_81),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_5),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_198),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_L g1052 ( 
.A(n_175),
.B(n_342),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_40),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_520),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_608),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_106),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_547),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_565),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_303),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_332),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_520),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_419),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_243),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_580),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_665),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_150),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_224),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_313),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_431),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_6),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_577),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_718),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_442),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_564),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_173),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_387),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_735),
.Y(n_1077)
);

BUFx10_ASAP7_75t_L g1078 ( 
.A(n_110),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_556),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_607),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_153),
.B(n_740),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_215),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_191),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_672),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_252),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_688),
.Y(n_1086)
);

CKINVDCx16_ASAP7_75t_R g1087 ( 
.A(n_71),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_226),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_286),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_571),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_750),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_448),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_685),
.Y(n_1093)
);

CKINVDCx14_ASAP7_75t_R g1094 ( 
.A(n_334),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_559),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_174),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_625),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_339),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_287),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_4),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_498),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_170),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_527),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_381),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_541),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_4),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_78),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_630),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_648),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_326),
.B(n_371),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_141),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_345),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_302),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_290),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_660),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_682),
.B(n_515),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_99),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_532),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_330),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_351),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_727),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_707),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_712),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_446),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_361),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_307),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_751),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_43),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_731),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_740),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_390),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_757),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_517),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_758),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_492),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_75),
.Y(n_1136)
);

BUFx2_ASAP7_75t_SL g1137 ( 
.A(n_50),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_828),
.B(n_0),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_849),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_796),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_839),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_911),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1106),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_849),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_911),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_849),
.Y(n_1146)
);

BUFx8_ASAP7_75t_L g1147 ( 
.A(n_827),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_828),
.Y(n_1148)
);

AND2x6_ASAP7_75t_L g1149 ( 
.A(n_835),
.B(n_0),
.Y(n_1149)
);

OAI22x1_ASAP7_75t_SL g1150 ( 
.A1(n_813),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_835),
.Y(n_1151)
);

BUFx8_ASAP7_75t_L g1152 ( 
.A(n_875),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_879),
.B(n_1),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_849),
.Y(n_1154)
);

INVxp33_ASAP7_75t_SL g1155 ( 
.A(n_975),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_879),
.B(n_2),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_796),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_843),
.B(n_2),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_892),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_796),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_849),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_809),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_846),
.B(n_3),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_918),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_809),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1094),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_918),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_922),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_809),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_786),
.A2(n_3),
.B(n_5),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_982),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_894),
.B(n_6),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1024),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_920),
.B(n_6),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1024),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_816),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_968),
.B(n_7),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_922),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_839),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1094),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1026),
.B(n_8),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1026),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_839),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_839),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1029),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_855),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1024),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_956),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_786),
.A2(n_9),
.B(n_10),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1029),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1024),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_909),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1044),
.B(n_10),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_909),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_878),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1044),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1024),
.Y(n_1197)
);

AOI22x1_ASAP7_75t_SL g1198 ( 
.A1(n_813),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_1198)
);

BUFx8_ASAP7_75t_SL g1199 ( 
.A(n_932),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_816),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_909),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1054),
.B(n_11),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_1055),
.B(n_14),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_897),
.B(n_14),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_909),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1055),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1004),
.B(n_15),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1058),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_904),
.B(n_15),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1058),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_936),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1089),
.B(n_16),
.Y(n_1212)
);

BUFx8_ASAP7_75t_SL g1213 ( 
.A(n_932),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1089),
.B(n_793),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_936),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_793),
.A2(n_16),
.B(n_17),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1050),
.B(n_17),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_936),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_959),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_802),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_819),
.Y(n_1221)
);

OAI22x1_ASAP7_75t_SL g1222 ( 
.A1(n_822),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_959),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_959),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1070),
.B(n_19),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_824),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1226)
);

AOI22x1_ASAP7_75t_SL g1227 ( 
.A1(n_822),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1227)
);

AOI22x1_ASAP7_75t_SL g1228 ( 
.A1(n_842),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_802),
.B(n_810),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_810),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1100),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1149),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1157),
.B(n_1046),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1166),
.B(n_1180),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1166),
.Y(n_1236)
);

OA22x2_ASAP7_75t_L g1237 ( 
.A1(n_1186),
.A2(n_826),
.B1(n_1098),
.B2(n_825),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1168),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1141),
.Y(n_1239)
);

CKINVDCx6p67_ASAP7_75t_R g1240 ( 
.A(n_1140),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1143),
.B(n_971),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1212),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1159),
.B(n_823),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_L g1244 ( 
.A(n_1149),
.B(n_971),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1212),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1206),
.B(n_1151),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1138),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1208),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1153),
.B(n_971),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1153),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1210),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1214),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1157),
.B(n_789),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1156),
.B(n_997),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1170),
.A2(n_781),
.B(n_778),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1186),
.A2(n_1000),
.B1(n_1009),
.B2(n_930),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1180),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1214),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1188),
.B(n_1027),
.Y(n_1259)
);

CKINVDCx16_ASAP7_75t_R g1260 ( 
.A(n_1160),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1156),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1181),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1181),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1145),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1231),
.Y(n_1265)
);

INVxp67_ASAP7_75t_SL g1266 ( 
.A(n_1163),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1215),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1193),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1162),
.B(n_1087),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1193),
.B(n_997),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1172),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1229),
.Y(n_1272)
);

NAND2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1207),
.B(n_907),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1139),
.B(n_997),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1229),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1162),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1164),
.B(n_831),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1172),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1144),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1146),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1154),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1174),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1165),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1174),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1161),
.Y(n_1285)
);

INVx8_ASAP7_75t_L g1286 ( 
.A(n_1176),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1141),
.Y(n_1287)
);

AND3x2_ASAP7_75t_L g1288 ( 
.A(n_1199),
.B(n_1017),
.C(n_844),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1163),
.B(n_997),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1173),
.B(n_1025),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1175),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1169),
.B(n_1123),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1177),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1191),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1197),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1158),
.Y(n_1297)
);

AOI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1187),
.A2(n_877),
.B(n_848),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1204),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1187),
.B(n_1025),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1184),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1167),
.B(n_779),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1184),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1178),
.B(n_1025),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1141),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1184),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1202),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1199),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1182),
.B(n_848),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1184),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1185),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1202),
.Y(n_1312)
);

NAND2xp33_ASAP7_75t_L g1313 ( 
.A(n_1149),
.B(n_1038),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1200),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1205),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1205),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1221),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1190),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1196),
.B(n_877),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1211),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1204),
.B(n_825),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1220),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1230),
.B(n_1038),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1179),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1203),
.Y(n_1325)
);

AO22x2_ASAP7_75t_L g1326 ( 
.A1(n_1198),
.A2(n_1137),
.B1(n_790),
.B2(n_901),
.Y(n_1326)
);

INVxp33_ASAP7_75t_SL g1327 ( 
.A(n_1209),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1217),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1155),
.B(n_882),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1179),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1217),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1189),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1225),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1225),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1155),
.B(n_887),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1149),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1183),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1213),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1149),
.B(n_888),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_L g1340 ( 
.A(n_1192),
.B(n_1038),
.Y(n_1340)
);

INVx8_ASAP7_75t_L g1341 ( 
.A(n_1213),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1147),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1171),
.B(n_780),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1195),
.B(n_888),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1216),
.Y(n_1345)
);

NOR2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1147),
.B(n_826),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1171),
.B(n_782),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1192),
.B(n_1051),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1152),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1194),
.B(n_917),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1201),
.B(n_791),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1218),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1152),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1219),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1219),
.B(n_1051),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1226),
.A2(n_929),
.B(n_921),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1223),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1223),
.B(n_792),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1224),
.B(n_954),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1224),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1224),
.Y(n_1362)
);

NOR2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1150),
.B(n_1098),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1195),
.B(n_954),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1227),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1228),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1222),
.B(n_1051),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1187),
.A2(n_966),
.B(n_962),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1212),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1187),
.A2(n_966),
.B(n_962),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1148),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1166),
.B(n_850),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1212),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1166),
.B(n_850),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1266),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1271),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1278),
.B(n_1282),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1255),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1284),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1265),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1293),
.B(n_979),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1294),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_L g1383 ( 
.A(n_1336),
.B(n_1091),
.Y(n_1383)
);

INVx8_ASAP7_75t_L g1384 ( 
.A(n_1286),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1307),
.B(n_799),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1314),
.B(n_25),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_1317),
.B(n_27),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1312),
.B(n_1328),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1331),
.B(n_800),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1333),
.B(n_801),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1334),
.B(n_803),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1259),
.B(n_1260),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_1336),
.B(n_1091),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1299),
.B(n_806),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1299),
.B(n_807),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1257),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_L g1397 ( 
.A(n_1353),
.B(n_1349),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1327),
.B(n_808),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1321),
.B(n_811),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1276),
.B(n_1283),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1265),
.B(n_988),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1311),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1311),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1247),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1232),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1250),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1342),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1261),
.B(n_829),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1353),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1262),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1286),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1235),
.B(n_988),
.Y(n_1412)
);

OR2x6_ASAP7_75t_L g1413 ( 
.A(n_1286),
.B(n_838),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1371),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1263),
.B(n_834),
.Y(n_1415)
);

INVx8_ASAP7_75t_L g1416 ( 
.A(n_1341),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1240),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1283),
.B(n_837),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1298),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1339),
.B(n_1095),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1268),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1343),
.B(n_991),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1236),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1368),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1264),
.B(n_1234),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1370),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1253),
.B(n_847),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1248),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1251),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1292),
.B(n_851),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1297),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1242),
.B(n_1095),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1292),
.B(n_852),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1246),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1245),
.B(n_1369),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1246),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1234),
.B(n_853),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1372),
.B(n_854),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1374),
.B(n_1373),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1269),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1344),
.A2(n_784),
.B1(n_787),
.B2(n_783),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1343),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1344),
.A2(n_788),
.B1(n_795),
.B2(n_794),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1322),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1318),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1252),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_L g1447 ( 
.A(n_1345),
.B(n_860),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_SL g1448 ( 
.A(n_1346),
.B(n_842),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1329),
.B(n_861),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1347),
.B(n_991),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1258),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1329),
.B(n_979),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1243),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1335),
.B(n_863),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1249),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1347),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1249),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1238),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_L g1459 ( 
.A(n_1332),
.B(n_1313),
.C(n_1244),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1302),
.B(n_865),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1254),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1254),
.B(n_996),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1270),
.B(n_996),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1270),
.B(n_999),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1300),
.A2(n_1290),
.B(n_1274),
.Y(n_1465)
);

AND2x2_ASAP7_75t_SL g1466 ( 
.A(n_1338),
.B(n_1014),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1244),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1289),
.B(n_999),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1277),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1325),
.B(n_870),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1309),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1272),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1275),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1237),
.A2(n_868),
.B1(n_872),
.B2(n_859),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1313),
.B(n_1110),
.C(n_798),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1364),
.B(n_805),
.C(n_797),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1364),
.B(n_859),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1273),
.B(n_871),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1289),
.B(n_1005),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1365),
.B(n_872),
.C(n_868),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1319),
.B(n_1267),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1351),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1279),
.B(n_814),
.C(n_812),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1280),
.B(n_1285),
.C(n_1281),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1351),
.B(n_1359),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1237),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1291),
.B(n_876),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1350),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1350),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1256),
.Y(n_1490)
);

AO221x1_ASAP7_75t_L g1491 ( 
.A1(n_1326),
.A2(n_893),
.B1(n_899),
.B2(n_891),
.C(n_889),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1326),
.A2(n_1130),
.B1(n_1133),
.B2(n_1125),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_1366),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1360),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1295),
.B(n_880),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_L g1496 ( 
.A(n_1296),
.B(n_881),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1241),
.B(n_883),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1360),
.B(n_817),
.C(n_815),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1356),
.B(n_884),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1326),
.B(n_991),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1363),
.B(n_889),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1301),
.B(n_1016),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1303),
.Y(n_1503)
);

NOR2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1341),
.B(n_1041),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1306),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1304),
.B(n_885),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1310),
.B(n_1016),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1315),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1367),
.B(n_804),
.C(n_785),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1316),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1323),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1304),
.B(n_886),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1367),
.B(n_890),
.Y(n_1513)
);

NAND2xp33_ASAP7_75t_SL g1514 ( 
.A(n_1308),
.B(n_891),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1300),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1274),
.B(n_895),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1320),
.B(n_1085),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1290),
.B(n_1085),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1288),
.B(n_1034),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1288),
.B(n_1034),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1341),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1239),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1348),
.B(n_1129),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1348),
.B(n_27),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1355),
.B(n_900),
.Y(n_1525)
);

NOR3xp33_ASAP7_75t_L g1526 ( 
.A(n_1355),
.B(n_858),
.C(n_820),
.Y(n_1526)
);

AND3x1_ASAP7_75t_L g1527 ( 
.A(n_1308),
.B(n_821),
.C(n_818),
.Y(n_1527)
);

OAI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1340),
.A2(n_950),
.B1(n_1082),
.B2(n_948),
.C(n_947),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1340),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1324),
.B(n_830),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1330),
.B(n_902),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_SL g1532 ( 
.A(n_1239),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1352),
.A2(n_833),
.B(n_836),
.C(n_832),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1354),
.B(n_1034),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1357),
.B(n_912),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1358),
.B(n_915),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1361),
.B(n_1099),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1362),
.A2(n_899),
.B1(n_905),
.B2(n_893),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_L g1539 ( 
.A(n_1239),
.B(n_840),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1239),
.B(n_1061),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1287),
.B(n_841),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1305),
.Y(n_1542)
);

BUFx10_ASAP7_75t_L g1543 ( 
.A(n_1305),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1337),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1337),
.B(n_926),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1233),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1266),
.B(n_927),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1271),
.B(n_928),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1266),
.B(n_931),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1266),
.B(n_934),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1266),
.B(n_1061),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1266),
.B(n_935),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1266),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1233),
.B(n_856),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1266),
.B(n_857),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1257),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1266),
.Y(n_1557)
);

INVx6_ASAP7_75t_L g1558 ( 
.A(n_1407),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1378),
.A2(n_864),
.B(n_862),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1380),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1384),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1377),
.B(n_938),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1546),
.B(n_939),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1442),
.B(n_1456),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1388),
.A2(n_867),
.B(n_866),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1546),
.B(n_941),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1557),
.B(n_942),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1538),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1376),
.A2(n_869),
.B(n_874),
.C(n_873),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1379),
.B(n_943),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1375),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1411),
.B(n_28),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1380),
.B(n_944),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1407),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1553),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1382),
.B(n_946),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1419),
.A2(n_898),
.B(n_896),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1405),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1384),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1490),
.A2(n_1440),
.B(n_1474),
.C(n_1486),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1425),
.A2(n_952),
.B1(n_953),
.B2(n_951),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1424),
.A2(n_908),
.B(n_903),
.Y(n_1582)
);

OR2x6_ASAP7_75t_L g1583 ( 
.A(n_1384),
.B(n_845),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1543),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1426),
.A2(n_913),
.B(n_910),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1411),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1439),
.A2(n_919),
.B(n_923),
.C(n_916),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1409),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1431),
.B(n_905),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1396),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1554),
.A2(n_925),
.B(n_924),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1389),
.A2(n_940),
.B(n_933),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1521),
.B(n_29),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1390),
.A2(n_949),
.B(n_945),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1453),
.A2(n_960),
.B(n_955),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1469),
.A2(n_1081),
.B(n_1052),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1423),
.B(n_906),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1391),
.A2(n_963),
.B(n_961),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1551),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1416),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1385),
.A2(n_970),
.B(n_967),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1417),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1416),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1392),
.B(n_906),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1471),
.Y(n_1605)
);

AO21x1_ASAP7_75t_L g1606 ( 
.A1(n_1499),
.A2(n_977),
.B(n_976),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1435),
.A2(n_980),
.B(n_978),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1434),
.B(n_958),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1481),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1447),
.A2(n_984),
.B(n_983),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1436),
.B(n_964),
.Y(n_1611)
);

OAI321xp33_ASAP7_75t_L g1612 ( 
.A1(n_1476),
.A2(n_1003),
.A3(n_989),
.B1(n_1006),
.B2(n_992),
.C(n_987),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1445),
.Y(n_1613)
);

AOI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1459),
.A2(n_1011),
.B(n_1007),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1444),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1484),
.A2(n_1023),
.B(n_1020),
.Y(n_1616)
);

AO21x1_ASAP7_75t_L g1617 ( 
.A1(n_1485),
.A2(n_1032),
.B(n_1028),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1547),
.A2(n_1036),
.B(n_1035),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1556),
.B(n_965),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1549),
.A2(n_1552),
.B(n_1550),
.Y(n_1620)
);

AND2x6_ASAP7_75t_L g1621 ( 
.A(n_1455),
.B(n_1039),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1504),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1398),
.B(n_914),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1543),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1555),
.B(n_969),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1402),
.A2(n_1043),
.B(n_1042),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1452),
.A2(n_1449),
.B(n_1454),
.C(n_1478),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1403),
.A2(n_1048),
.B(n_1047),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1395),
.A2(n_981),
.B(n_973),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1548),
.B(n_985),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1404),
.A2(n_937),
.B1(n_957),
.B2(n_914),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1381),
.A2(n_1057),
.B(n_1049),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1406),
.Y(n_1633)
);

AND2x2_ASAP7_75t_SL g1634 ( 
.A(n_1466),
.B(n_937),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1488),
.A2(n_1060),
.B(n_1059),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1510),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1489),
.A2(n_1065),
.B(n_1064),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1477),
.A2(n_990),
.B1(n_994),
.B2(n_986),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1410),
.B(n_998),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1401),
.B(n_1001),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1476),
.A2(n_972),
.B1(n_974),
.B2(n_957),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1494),
.A2(n_1069),
.B(n_1067),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1412),
.B(n_972),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1422),
.B(n_974),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1408),
.A2(n_1415),
.B(n_1457),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1461),
.A2(n_1076),
.B(n_1075),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1458),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1421),
.B(n_1002),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1450),
.B(n_993),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1475),
.A2(n_1088),
.B(n_1086),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1482),
.B(n_1008),
.Y(n_1651)
);

INVx8_ASAP7_75t_L g1652 ( 
.A(n_1416),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1394),
.B(n_993),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1510),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1538),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1475),
.A2(n_1093),
.B(n_1090),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1467),
.A2(n_1105),
.B(n_1096),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1500),
.A2(n_1012),
.B1(n_1030),
.B2(n_995),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1514),
.Y(n_1659)
);

AO21x1_ASAP7_75t_L g1660 ( 
.A1(n_1468),
.A2(n_1479),
.B(n_1400),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1542),
.Y(n_1661)
);

OR2x6_ASAP7_75t_SL g1662 ( 
.A(n_1448),
.B(n_1010),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1441),
.A2(n_1012),
.B1(n_1030),
.B2(n_995),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1428),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1397),
.B(n_1116),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1438),
.B(n_1031),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1399),
.B(n_1013),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1443),
.B(n_1031),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1501),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1498),
.A2(n_1115),
.B(n_1113),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1542),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1446),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1429),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1427),
.A2(n_1117),
.B(n_1120),
.Y(n_1674)
);

BUFx4f_ASAP7_75t_L g1675 ( 
.A(n_1413),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1430),
.A2(n_1124),
.B(n_1121),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1437),
.B(n_1037),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1433),
.A2(n_1127),
.B(n_1126),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1472),
.A2(n_1040),
.B1(n_1062),
.B2(n_1037),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_L g1680 ( 
.A(n_1515),
.B(n_1015),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1509),
.B(n_1496),
.C(n_1492),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1527),
.Y(n_1682)
);

NOR2xp67_ASAP7_75t_L g1683 ( 
.A(n_1480),
.B(n_30),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1460),
.B(n_1040),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1462),
.A2(n_1132),
.B(n_1131),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1463),
.A2(n_1136),
.B(n_1135),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1473),
.B(n_1018),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1493),
.B(n_1062),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1542),
.Y(n_1689)
);

INVx11_ASAP7_75t_L g1690 ( 
.A(n_1386),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1473),
.B(n_1019),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1464),
.A2(n_1022),
.B(n_1021),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1491),
.B(n_1072),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1451),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1534),
.B(n_1072),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1470),
.B(n_1102),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1413),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_L g1698 ( 
.A(n_1513),
.B(n_1112),
.C(n_1033),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1418),
.B(n_1045),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1413),
.B(n_1495),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_SL g1701 ( 
.A(n_1526),
.B(n_1114),
.C(n_1109),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1527),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1487),
.A2(n_1056),
.B(n_1053),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1519),
.B(n_1080),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1520),
.B(n_1080),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1387),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1483),
.B(n_1063),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1498),
.A2(n_1068),
.B(n_1071),
.C(n_1066),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1511),
.A2(n_1074),
.B(n_1073),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1483),
.B(n_1077),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1537),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1518),
.A2(n_1083),
.B(n_1079),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1540),
.B(n_1084),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1516),
.A2(n_1092),
.B1(n_1101),
.B2(n_1097),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1530),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1530),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1497),
.B(n_1084),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1506),
.B(n_1512),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1528),
.Y(n_1719)
);

NOR2xp67_ASAP7_75t_L g1720 ( 
.A(n_1518),
.B(n_31),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1414),
.A2(n_1107),
.B1(n_1109),
.B2(n_1103),
.Y(n_1721)
);

NAND2x1_ASAP7_75t_L g1722 ( 
.A(n_1539),
.B(n_1128),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1525),
.A2(n_1104),
.B1(n_1111),
.B2(n_1108),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1503),
.A2(n_1107),
.B1(n_1114),
.B2(n_1103),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1383),
.A2(n_1134),
.B(n_1118),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1505),
.B(n_1119),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1393),
.A2(n_1122),
.B(n_1119),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_R g1728 ( 
.A(n_1532),
.B(n_1078),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1508),
.B(n_1128),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1545),
.A2(n_32),
.B(n_34),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1533),
.B(n_34),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1502),
.B(n_35),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1523),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1507),
.B(n_39),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1517),
.B(n_776),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1535),
.B(n_41),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1536),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1432),
.A2(n_42),
.B(n_44),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1531),
.B(n_45),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1523),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1529),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1541),
.A2(n_49),
.B(n_52),
.Y(n_1742)
);

CKINVDCx6p67_ASAP7_75t_R g1743 ( 
.A(n_1532),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1544),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1465),
.A2(n_53),
.B(n_54),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1465),
.A2(n_54),
.B(n_55),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1524),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1522),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1378),
.A2(n_762),
.B(n_759),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1388),
.A2(n_61),
.B(n_62),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1411),
.B(n_61),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1411),
.B(n_63),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1377),
.B(n_64),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1546),
.B(n_64),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1388),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1388),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1377),
.B(n_67),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1384),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1377),
.B(n_70),
.Y(n_1759)
);

INVx11_ASAP7_75t_L g1760 ( 
.A(n_1407),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1388),
.A2(n_70),
.B(n_71),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1388),
.A2(n_72),
.B(n_73),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1377),
.B(n_72),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1546),
.B(n_73),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1380),
.B(n_773),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1377),
.B(n_74),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1388),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1384),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1380),
.B(n_773),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1388),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1377),
.B(n_75),
.Y(n_1771)
);

BUFx12f_ASAP7_75t_L g1772 ( 
.A(n_1407),
.Y(n_1772)
);

AOI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1420),
.A2(n_76),
.B(n_77),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1377),
.B(n_79),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1377),
.B(n_82),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1546),
.Y(n_1776)
);

A2O1A1Ixp33_ASAP7_75t_L g1777 ( 
.A1(n_1377),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1378),
.A2(n_83),
.B(n_85),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1377),
.B(n_85),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1388),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_SL g1781 ( 
.A1(n_1559),
.A2(n_86),
.B(n_87),
.Y(n_1781)
);

AO31x2_ASAP7_75t_L g1782 ( 
.A1(n_1606),
.A2(n_90),
.A3(n_87),
.B(n_88),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1574),
.Y(n_1783)
);

OAI22x1_ASAP7_75t_L g1784 ( 
.A1(n_1655),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1767),
.A2(n_91),
.B(n_92),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1645),
.A2(n_93),
.B(n_94),
.Y(n_1786)
);

AOI21x1_ASAP7_75t_L g1787 ( 
.A1(n_1660),
.A2(n_93),
.B(n_94),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1770),
.A2(n_95),
.B(n_96),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1760),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1780),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1661),
.Y(n_1791)
);

AND2x6_ASAP7_75t_L g1792 ( 
.A(n_1609),
.B(n_1768),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1713),
.B(n_95),
.Y(n_1793)
);

AOI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1596),
.A2(n_97),
.B(n_98),
.Y(n_1794)
);

CKINVDCx16_ASAP7_75t_R g1795 ( 
.A(n_1772),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1564),
.B(n_99),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1560),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1652),
.B(n_100),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1605),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1613),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1575),
.B(n_101),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1615),
.B(n_102),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1633),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1599),
.B(n_104),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1568),
.B(n_105),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1749),
.A2(n_105),
.B(n_106),
.Y(n_1806)
);

CKINVDCx8_ASAP7_75t_R g1807 ( 
.A(n_1652),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1558),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1595),
.B(n_107),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1577),
.A2(n_107),
.B(n_108),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1558),
.Y(n_1811)
);

A2O1A1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1627),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1625),
.B(n_111),
.Y(n_1813)
);

AO21x2_ASAP7_75t_L g1814 ( 
.A1(n_1745),
.A2(n_112),
.B(n_114),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1582),
.A2(n_115),
.B(n_116),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1585),
.A2(n_116),
.B(n_117),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1600),
.B(n_1758),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1578),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1746),
.B(n_1778),
.C(n_1681),
.Y(n_1819)
);

AOI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1773),
.A2(n_118),
.B(n_119),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1588),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1571),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1715),
.A2(n_1716),
.B1(n_1757),
.B2(n_1753),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1632),
.B(n_121),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1618),
.B(n_122),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1664),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1579),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1635),
.B(n_123),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1637),
.B(n_124),
.Y(n_1829)
);

OAI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1677),
.A2(n_124),
.B(n_125),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1642),
.B(n_128),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_SL g1832 ( 
.A1(n_1617),
.A2(n_128),
.B(n_129),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1565),
.B(n_130),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1672),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1561),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1592),
.A2(n_135),
.B(n_132),
.C(n_133),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1718),
.A2(n_1611),
.B(n_1608),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1661),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1652),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1694),
.B(n_1594),
.Y(n_1840)
);

AO21x1_ASAP7_75t_L g1841 ( 
.A1(n_1730),
.A2(n_136),
.B(n_137),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1598),
.B(n_137),
.Y(n_1842)
);

AND2x6_ASAP7_75t_SL g1843 ( 
.A(n_1604),
.B(n_138),
.Y(n_1843)
);

BUFx12f_ASAP7_75t_L g1844 ( 
.A(n_1602),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1622),
.Y(n_1845)
);

BUFx12f_ASAP7_75t_L g1846 ( 
.A(n_1600),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1584),
.B(n_140),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1601),
.B(n_142),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1711),
.B(n_142),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1759),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1603),
.B(n_143),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1661),
.A2(n_144),
.B(n_145),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1724),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_SL g1854 ( 
.A(n_1584),
.B(n_146),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1743),
.Y(n_1855)
);

OAI21x1_ASAP7_75t_SL g1856 ( 
.A1(n_1763),
.A2(n_147),
.B(n_148),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1671),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1580),
.B(n_147),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1624),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1616),
.A2(n_150),
.B(n_151),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1671),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1668),
.B(n_1726),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1650),
.A2(n_1656),
.B(n_1674),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1676),
.A2(n_155),
.B(n_156),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1717),
.B(n_157),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1766),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1717),
.B(n_158),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1771),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1624),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1671),
.Y(n_1870)
);

OR2x6_ASAP7_75t_L g1871 ( 
.A(n_1586),
.B(n_1659),
.Y(n_1871)
);

OA21x2_ASAP7_75t_L g1872 ( 
.A1(n_1739),
.A2(n_161),
.B(n_162),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1624),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1673),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1684),
.B(n_1678),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1670),
.A2(n_164),
.B(n_165),
.Y(n_1876)
);

AOI211x1_ASAP7_75t_L g1877 ( 
.A1(n_1750),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1587),
.A2(n_172),
.B(n_169),
.C(n_171),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1774),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1776),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1728),
.B(n_178),
.Y(n_1881)
);

BUFx8_ASAP7_75t_L g1882 ( 
.A(n_1682),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1657),
.A2(n_179),
.B(n_180),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1653),
.B(n_181),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1775),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_1885)
);

AND3x4_ASAP7_75t_L g1886 ( 
.A(n_1683),
.B(n_185),
.C(n_186),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1752),
.B(n_1590),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1720),
.A2(n_187),
.B(n_188),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1779),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1688),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1776),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1646),
.A2(n_189),
.B(n_190),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1736),
.A2(n_1610),
.B(n_1762),
.C(n_1761),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1662),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1765),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1626),
.A2(n_191),
.B(n_192),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1628),
.B(n_192),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1623),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1675),
.Y(n_1899)
);

AOI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1720),
.A2(n_195),
.B(n_196),
.Y(n_1900)
);

AND2x2_ASAP7_75t_SL g1901 ( 
.A(n_1634),
.B(n_196),
.Y(n_1901)
);

OR2x6_ASAP7_75t_L g1902 ( 
.A(n_1663),
.B(n_197),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1569),
.B(n_197),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1621),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1732),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1647),
.Y(n_1906)
);

OAI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1708),
.A2(n_199),
.B(n_200),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1732),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1666),
.B(n_200),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1777),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1612),
.A2(n_204),
.B(n_207),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1689),
.A2(n_208),
.B(n_209),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1734),
.Y(n_1913)
);

AO31x2_ASAP7_75t_L g1914 ( 
.A1(n_1741),
.A2(n_213),
.A3(n_211),
.B(n_212),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1621),
.B(n_212),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1689),
.A2(n_213),
.B(n_215),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1631),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1607),
.A2(n_216),
.B(n_217),
.Y(n_1918)
);

OAI21xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1572),
.A2(n_220),
.B(n_219),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1731),
.A2(n_222),
.B1(n_218),
.B2(n_221),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1702),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1570),
.A2(n_223),
.B(n_224),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1636),
.A2(n_225),
.B(n_227),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1695),
.B(n_228),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1744),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1679),
.B(n_228),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1695),
.B(n_230),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1722),
.A2(n_1764),
.B(n_1754),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1562),
.B(n_231),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1576),
.A2(n_232),
.B(n_233),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1621),
.Y(n_1931)
);

BUFx10_ASAP7_75t_L g1932 ( 
.A(n_1589),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1729),
.B(n_235),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1698),
.B(n_236),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1748),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1712),
.A2(n_239),
.B(n_240),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1563),
.B(n_240),
.Y(n_1937)
);

OR2x6_ASAP7_75t_L g1938 ( 
.A(n_1751),
.B(n_241),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1621),
.B(n_1639),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1734),
.Y(n_1940)
);

OAI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1591),
.A2(n_241),
.B(n_242),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1597),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_SL g1943 ( 
.A1(n_1747),
.A2(n_243),
.B(n_244),
.Y(n_1943)
);

BUFx5_ASAP7_75t_L g1944 ( 
.A(n_1735),
.Y(n_1944)
);

OAI21x1_ASAP7_75t_SL g1945 ( 
.A1(n_1756),
.A2(n_245),
.B(n_246),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1733),
.A2(n_247),
.B(n_248),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1572),
.Y(n_1947)
);

OR2x6_ASAP7_75t_L g1948 ( 
.A(n_1583),
.B(n_249),
.Y(n_1948)
);

AO21x1_ASAP7_75t_L g1949 ( 
.A1(n_1740),
.A2(n_249),
.B(n_250),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1648),
.B(n_250),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1636),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1769),
.B(n_252),
.Y(n_1952)
);

AO31x2_ASAP7_75t_L g1953 ( 
.A1(n_1737),
.A2(n_1742),
.A3(n_1686),
.B(n_1685),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1675),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1643),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1690),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1687),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1707),
.B(n_256),
.Y(n_1958)
);

AO31x2_ASAP7_75t_L g1959 ( 
.A1(n_1738),
.A2(n_260),
.A3(n_258),
.B(n_259),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1703),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1691),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1644),
.B(n_262),
.Y(n_1962)
);

OA22x2_ASAP7_75t_L g1963 ( 
.A1(n_1693),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1669),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1649),
.B(n_265),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1710),
.B(n_267),
.Y(n_1966)
);

AND3x4_ASAP7_75t_L g1967 ( 
.A(n_1593),
.B(n_267),
.C(n_268),
.Y(n_1967)
);

OAI22x1_ASAP7_75t_L g1968 ( 
.A1(n_1638),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1705),
.B(n_271),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1641),
.B(n_1658),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1709),
.A2(n_272),
.B(n_273),
.Y(n_1971)
);

INVx4_ASAP7_75t_L g1972 ( 
.A(n_1654),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1667),
.B(n_274),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1727),
.B(n_274),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1567),
.A2(n_275),
.B(n_276),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1700),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1654),
.Y(n_1977)
);

AOI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1699),
.A2(n_281),
.B(n_282),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1583),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1630),
.B(n_283),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1629),
.B(n_284),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1696),
.B(n_285),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1583),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1581),
.B(n_288),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1721),
.B(n_289),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1566),
.Y(n_1986)
);

AOI221xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1680),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.C(n_294),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1651),
.A2(n_292),
.B(n_293),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1640),
.A2(n_296),
.B(n_297),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1701),
.B(n_296),
.Y(n_1990)
);

AO31x2_ASAP7_75t_L g1991 ( 
.A1(n_1692),
.A2(n_300),
.A3(n_297),
.B(n_298),
.Y(n_1991)
);

AOI21xp33_ASAP7_75t_L g1992 ( 
.A1(n_1665),
.A2(n_298),
.B(n_303),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1706),
.A2(n_307),
.B1(n_304),
.B2(n_305),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1714),
.B(n_304),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_R g1995 ( 
.A(n_1697),
.B(n_305),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1619),
.A2(n_309),
.B(n_310),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1573),
.Y(n_1997)
);

INVx5_ASAP7_75t_L g1998 ( 
.A(n_1725),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1723),
.A2(n_309),
.B(n_310),
.Y(n_1999)
);

AOI21xp33_ASAP7_75t_L g2000 ( 
.A1(n_1704),
.A2(n_311),
.B(n_312),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1755),
.B(n_314),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1755),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1755),
.B(n_314),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1755),
.B(n_315),
.Y(n_2004)
);

O2A1O1Ixp5_ASAP7_75t_L g2005 ( 
.A1(n_1606),
.A2(n_319),
.B(n_317),
.C(n_318),
.Y(n_2005)
);

INVxp67_ASAP7_75t_SL g2006 ( 
.A(n_1755),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1755),
.B(n_320),
.Y(n_2007)
);

AO31x2_ASAP7_75t_L g2008 ( 
.A1(n_1606),
.A2(n_324),
.A3(n_322),
.B(n_323),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1755),
.B(n_322),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1755),
.Y(n_2010)
);

OAI22x1_ASAP7_75t_L g2011 ( 
.A1(n_1655),
.A2(n_326),
.B1(n_323),
.B2(n_325),
.Y(n_2011)
);

A2O1A1Ixp33_ASAP7_75t_L g2012 ( 
.A1(n_1620),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_2012)
);

AO31x2_ASAP7_75t_L g2013 ( 
.A1(n_1606),
.A2(n_331),
.A3(n_329),
.B(n_330),
.Y(n_2013)
);

O2A1O1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1719),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2014)
);

NOR2x1_ASAP7_75t_SL g2015 ( 
.A(n_1600),
.B(n_336),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1560),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1755),
.B(n_337),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1755),
.B(n_339),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1620),
.A2(n_340),
.B(n_341),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1760),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1713),
.B(n_343),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1760),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1755),
.Y(n_2023)
);

OAI21x1_ASAP7_75t_L g2024 ( 
.A1(n_1614),
.A2(n_345),
.B(n_346),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1620),
.A2(n_346),
.B(n_347),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_L g2026 ( 
.A(n_1574),
.B(n_347),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1620),
.A2(n_348),
.B(n_349),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1755),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1713),
.B(n_352),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1780),
.B(n_352),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1755),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1713),
.B(n_354),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1620),
.A2(n_355),
.B(n_356),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1755),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1755),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1755),
.Y(n_2036)
);

BUFx2_ASAP7_75t_L g2037 ( 
.A(n_1560),
.Y(n_2037)
);

INVx5_ASAP7_75t_L g2038 ( 
.A(n_1584),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_L g2039 ( 
.A(n_1596),
.B(n_357),
.C(n_358),
.Y(n_2039)
);

BUFx8_ASAP7_75t_L g2040 ( 
.A(n_1574),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1755),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1780),
.B(n_359),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1780),
.B(n_360),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1780),
.B(n_360),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1755),
.B(n_361),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1620),
.A2(n_362),
.B(n_363),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1755),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1755),
.B(n_364),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1755),
.B(n_366),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1564),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1755),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1780),
.B(n_372),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_SL g2053 ( 
.A(n_1634),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_SL g2054 ( 
.A1(n_1559),
.A2(n_373),
.B(n_374),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1755),
.Y(n_2055)
);

NOR2x1_ASAP7_75t_SL g2056 ( 
.A(n_1600),
.B(n_376),
.Y(n_2056)
);

AOI211x1_ASAP7_75t_L g2057 ( 
.A1(n_1617),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1620),
.A2(n_377),
.B(n_379),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1780),
.B(n_380),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1780),
.B(n_382),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1620),
.A2(n_383),
.B(n_384),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1780),
.B(n_384),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1755),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1620),
.A2(n_385),
.B(n_386),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1780),
.B(n_388),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1614),
.A2(n_389),
.B(n_391),
.Y(n_2066)
);

AOI221xp5_ASAP7_75t_L g2067 ( 
.A1(n_1564),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.C(n_395),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_1755),
.B(n_395),
.Y(n_2068)
);

NAND2x1p5_ASAP7_75t_L g2069 ( 
.A(n_1600),
.B(n_396),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_1574),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1620),
.A2(n_397),
.B(n_398),
.Y(n_2071)
);

NAND2x1p5_ASAP7_75t_L g2072 ( 
.A(n_1600),
.B(n_398),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1620),
.A2(n_399),
.B(n_400),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1620),
.A2(n_399),
.B(n_400),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1620),
.A2(n_401),
.B(n_402),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1760),
.Y(n_2076)
);

NAND2x1p5_ASAP7_75t_L g2077 ( 
.A(n_1600),
.B(n_401),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1755),
.B(n_402),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1620),
.A2(n_403),
.B(n_404),
.Y(n_2079)
);

INVx3_ASAP7_75t_SL g2080 ( 
.A(n_1558),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1755),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1620),
.A2(n_405),
.B(n_406),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1755),
.B(n_407),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1755),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1631),
.B(n_409),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_1652),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1755),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1578),
.Y(n_2088)
);

NOR2xp67_ASAP7_75t_L g2089 ( 
.A(n_1574),
.B(n_410),
.Y(n_2089)
);

AO21x1_ASAP7_75t_L g2090 ( 
.A1(n_1745),
.A2(n_412),
.B(n_413),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1755),
.B(n_413),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1755),
.B(n_414),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1755),
.B(n_416),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1564),
.A2(n_420),
.B1(n_417),
.B2(n_419),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1755),
.B(n_420),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_1620),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1620),
.A2(n_424),
.B(n_425),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_SL g2098 ( 
.A1(n_1559),
.A2(n_424),
.B(n_425),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1661),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_1620),
.A2(n_430),
.B(n_426),
.C(n_427),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1652),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1780),
.B(n_432),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1755),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1755),
.B(n_434),
.Y(n_2104)
);

BUFx6f_ASAP7_75t_L g2105 ( 
.A(n_1661),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1780),
.B(n_437),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1780),
.B(n_437),
.Y(n_2107)
);

OAI22x1_ASAP7_75t_L g2108 ( 
.A1(n_1655),
.A2(n_441),
.B1(n_438),
.B2(n_439),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1780),
.B(n_443),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1584),
.Y(n_2110)
);

OAI21x1_ASAP7_75t_SL g2111 ( 
.A1(n_1559),
.A2(n_443),
.B(n_444),
.Y(n_2111)
);

AO21x2_ASAP7_75t_L g2112 ( 
.A1(n_1745),
.A2(n_445),
.B(n_446),
.Y(n_2112)
);

AO31x2_ASAP7_75t_L g2113 ( 
.A1(n_1606),
.A2(n_450),
.A3(n_447),
.B(n_449),
.Y(n_2113)
);

NOR2xp67_ASAP7_75t_L g2114 ( 
.A(n_1574),
.B(n_449),
.Y(n_2114)
);

NAND2x1p5_ASAP7_75t_L g2115 ( 
.A(n_1600),
.B(n_454),
.Y(n_2115)
);

OAI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_1620),
.A2(n_456),
.B(n_457),
.Y(n_2116)
);

OR2x6_ASAP7_75t_L g2117 ( 
.A(n_1652),
.B(n_459),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1620),
.A2(n_459),
.B(n_460),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1755),
.B(n_460),
.Y(n_2119)
);

INVx5_ASAP7_75t_L g2120 ( 
.A(n_1584),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1755),
.B(n_461),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1713),
.B(n_462),
.Y(n_2122)
);

BUFx3_ASAP7_75t_L g2123 ( 
.A(n_1574),
.Y(n_2123)
);

AND3x4_ASAP7_75t_L g2124 ( 
.A(n_1683),
.B(n_464),
.C(n_465),
.Y(n_2124)
);

AOI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_1564),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_1560),
.Y(n_2126)
);

OA22x2_ASAP7_75t_L g2127 ( 
.A1(n_1655),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_2127)
);

AND3x4_ASAP7_75t_L g2128 ( 
.A(n_1683),
.B(n_469),
.C(n_470),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_SL g2129 ( 
.A1(n_1559),
.A2(n_470),
.B(n_471),
.Y(n_2129)
);

AO31x2_ASAP7_75t_L g2130 ( 
.A1(n_1606),
.A2(n_475),
.A3(n_473),
.B(n_474),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1755),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_1652),
.Y(n_2132)
);

OAI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1620),
.A2(n_476),
.B(n_477),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1755),
.B(n_476),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_1564),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_2135)
);

OAI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1620),
.A2(n_478),
.B(n_479),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1755),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_SL g2138 ( 
.A(n_1755),
.B(n_484),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_1846),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1859),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1790),
.Y(n_2141)
);

BUFx2_ASAP7_75t_R g2142 ( 
.A(n_1807),
.Y(n_2142)
);

INVx3_ASAP7_75t_L g2143 ( 
.A(n_2132),
.Y(n_2143)
);

NAND3xp33_ASAP7_75t_L g2144 ( 
.A(n_1877),
.B(n_485),
.C(n_486),
.Y(n_2144)
);

BUFx4f_ASAP7_75t_SL g2145 ( 
.A(n_2040),
.Y(n_2145)
);

AOI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_1917),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.C(n_490),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1859),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_2002),
.B(n_488),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2034),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1859),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_1798),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2047),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_2040),
.Y(n_2153)
);

AO21x2_ASAP7_75t_L g2154 ( 
.A1(n_1819),
.A2(n_491),
.B(n_493),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2010),
.B(n_494),
.Y(n_2155)
);

OA21x2_ASAP7_75t_L g2156 ( 
.A1(n_1819),
.A2(n_495),
.B(n_496),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_SL g2157 ( 
.A1(n_2025),
.A2(n_497),
.B(n_498),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2010),
.B(n_497),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_1783),
.Y(n_2159)
);

OA21x2_ASAP7_75t_L g2160 ( 
.A1(n_1806),
.A2(n_499),
.B(n_500),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1837),
.A2(n_499),
.B(n_500),
.Y(n_2161)
);

AOI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1787),
.A2(n_1823),
.B(n_1947),
.Y(n_2162)
);

OR2x6_ASAP7_75t_L g2163 ( 
.A(n_1798),
.B(n_501),
.Y(n_2163)
);

OR2x6_ASAP7_75t_L g2164 ( 
.A(n_1798),
.B(n_501),
.Y(n_2164)
);

AO21x2_ASAP7_75t_L g2165 ( 
.A1(n_2025),
.A2(n_502),
.B(n_503),
.Y(n_2165)
);

NAND3xp33_ASAP7_75t_L g2166 ( 
.A(n_1987),
.B(n_503),
.C(n_504),
.Y(n_2166)
);

BUFx12f_ASAP7_75t_L g2167 ( 
.A(n_1789),
.Y(n_2167)
);

AO21x2_ASAP7_75t_L g2168 ( 
.A1(n_2046),
.A2(n_504),
.B(n_505),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2006),
.B(n_508),
.Y(n_2169)
);

INVx1_ASAP7_75t_SL g2170 ( 
.A(n_1797),
.Y(n_2170)
);

INVx4_ASAP7_75t_L g2171 ( 
.A(n_1859),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_L g2172 ( 
.A(n_1987),
.B(n_1893),
.C(n_2057),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2051),
.Y(n_2173)
);

NAND2x1p5_ASAP7_75t_L g2174 ( 
.A(n_2038),
.B(n_510),
.Y(n_2174)
);

OR2x6_ASAP7_75t_L g2175 ( 
.A(n_2117),
.B(n_510),
.Y(n_2175)
);

AO21x2_ASAP7_75t_L g2176 ( 
.A1(n_2046),
.A2(n_511),
.B(n_512),
.Y(n_2176)
);

OA21x2_ASAP7_75t_L g2177 ( 
.A1(n_2116),
.A2(n_511),
.B(n_513),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_1797),
.B(n_513),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2038),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_2117),
.B(n_1839),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_1862),
.B(n_514),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_2038),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2055),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1863),
.A2(n_1840),
.B(n_2136),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_2123),
.Y(n_2185)
);

INVx1_ASAP7_75t_SL g2186 ( 
.A(n_2016),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_1977),
.A2(n_514),
.B(n_515),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_SL g2188 ( 
.A1(n_2116),
.A2(n_516),
.B(n_517),
.Y(n_2188)
);

INVx4_ASAP7_75t_L g2189 ( 
.A(n_2038),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_1821),
.B(n_516),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_1977),
.A2(n_518),
.B(n_519),
.Y(n_2191)
);

OA21x2_ASAP7_75t_L g2192 ( 
.A1(n_2118),
.A2(n_518),
.B(n_522),
.Y(n_2192)
);

AOI21xp33_ASAP7_75t_L g2193 ( 
.A1(n_1858),
.A2(n_522),
.B(n_523),
.Y(n_2193)
);

BUFx2_ASAP7_75t_R g2194 ( 
.A(n_2020),
.Y(n_2194)
);

NOR2x1_ASAP7_75t_R g2195 ( 
.A(n_2022),
.B(n_526),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2081),
.B(n_527),
.Y(n_2196)
);

INVx3_ASAP7_75t_L g2197 ( 
.A(n_2120),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_2120),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2084),
.B(n_528),
.Y(n_2199)
);

CKINVDCx11_ASAP7_75t_R g2200 ( 
.A(n_2070),
.Y(n_2200)
);

NAND2x1_ASAP7_75t_L g2201 ( 
.A(n_1792),
.B(n_528),
.Y(n_2201)
);

OA21x2_ASAP7_75t_L g2202 ( 
.A1(n_2118),
.A2(n_529),
.B(n_530),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_2023),
.B(n_531),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_2028),
.B(n_531),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1970),
.B(n_533),
.Y(n_2205)
);

BUFx3_ASAP7_75t_L g2206 ( 
.A(n_2120),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_2031),
.B(n_534),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2087),
.B(n_534),
.Y(n_2208)
);

OA21x2_ASAP7_75t_L g2209 ( 
.A1(n_2133),
.A2(n_535),
.B(n_536),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2035),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_1820),
.A2(n_537),
.B(n_538),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2036),
.B(n_538),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_2120),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2041),
.B(n_539),
.Y(n_2214)
);

AO21x2_ASAP7_75t_L g2215 ( 
.A1(n_2133),
.A2(n_541),
.B(n_543),
.Y(n_2215)
);

OA21x2_ASAP7_75t_L g2216 ( 
.A1(n_2136),
.A2(n_545),
.B(n_546),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_SL g2217 ( 
.A1(n_1785),
.A2(n_545),
.B(n_548),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2063),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_1795),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1875),
.A2(n_549),
.B(n_550),
.Y(n_2220)
);

NAND3xp33_ASAP7_75t_L g2221 ( 
.A(n_1812),
.B(n_551),
.C(n_552),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_2117),
.Y(n_2222)
);

INVx4_ASAP7_75t_SL g2223 ( 
.A(n_1792),
.Y(n_2223)
);

OA21x2_ASAP7_75t_L g2224 ( 
.A1(n_2090),
.A2(n_551),
.B(n_553),
.Y(n_2224)
);

INVx3_ASAP7_75t_SL g2225 ( 
.A(n_2076),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1791),
.Y(n_2226)
);

BUFx8_ASAP7_75t_L g2227 ( 
.A(n_2053),
.Y(n_2227)
);

BUFx12f_ASAP7_75t_L g2228 ( 
.A(n_1808),
.Y(n_2228)
);

OR2x6_ASAP7_75t_L g2229 ( 
.A(n_1902),
.B(n_554),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2103),
.Y(n_2230)
);

AO21x2_ASAP7_75t_L g2231 ( 
.A1(n_1814),
.A2(n_555),
.B(n_556),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2131),
.B(n_557),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1818),
.B(n_558),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1799),
.B(n_1800),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1803),
.B(n_560),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2001),
.Y(n_2236)
);

AOI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_1850),
.A2(n_561),
.B(n_562),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_2037),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_1869),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2001),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1942),
.B(n_561),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1838),
.Y(n_2242)
);

OA21x2_ASAP7_75t_L g2243 ( 
.A1(n_2024),
.A2(n_565),
.B(n_566),
.Y(n_2243)
);

AO21x2_ASAP7_75t_L g2244 ( 
.A1(n_1814),
.A2(n_566),
.B(n_567),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_2126),
.Y(n_2245)
);

BUFx3_ASAP7_75t_L g2246 ( 
.A(n_1873),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_1901),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1869),
.Y(n_2248)
);

OR2x6_ASAP7_75t_L g2249 ( 
.A(n_1902),
.B(n_573),
.Y(n_2249)
);

OR2x6_ASAP7_75t_L g2250 ( 
.A(n_1902),
.B(n_574),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2053),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_2251)
);

AOI22x1_ASAP7_75t_L g2252 ( 
.A1(n_2019),
.A2(n_575),
.B1(n_577),
.B2(n_578),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_2066),
.A2(n_578),
.B(n_579),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2003),
.Y(n_2254)
);

CKINVDCx6p67_ASAP7_75t_R g2255 ( 
.A(n_2080),
.Y(n_2255)
);

NOR2x1_ASAP7_75t_L g2256 ( 
.A(n_1967),
.B(n_583),
.Y(n_2256)
);

INVx5_ASAP7_75t_SL g2257 ( 
.A(n_1948),
.Y(n_2257)
);

NAND2x1p5_ASAP7_75t_L g2258 ( 
.A(n_2086),
.B(n_583),
.Y(n_2258)
);

OAI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_1863),
.A2(n_585),
.B(n_586),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_1868),
.A2(n_587),
.B(n_588),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_1853),
.B(n_588),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_1792),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_1855),
.Y(n_2263)
);

NAND2x1p5_ASAP7_75t_L g2264 ( 
.A(n_2101),
.B(n_589),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_1817),
.B(n_589),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_SL g2266 ( 
.A1(n_1785),
.A2(n_590),
.B(n_591),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_1817),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2004),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1845),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_SL g2270 ( 
.A1(n_1788),
.A2(n_593),
.B(n_594),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2110),
.Y(n_2271)
);

CKINVDCx11_ASAP7_75t_R g2272 ( 
.A(n_1844),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1857),
.Y(n_2273)
);

AO21x2_ASAP7_75t_L g2274 ( 
.A1(n_2112),
.A2(n_595),
.B(n_596),
.Y(n_2274)
);

NAND3x1_ASAP7_75t_L g2275 ( 
.A(n_1990),
.B(n_596),
.C(n_597),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2004),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1889),
.B(n_600),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2009),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2009),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2017),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_1811),
.Y(n_2281)
);

INVx2_ASAP7_75t_SL g2282 ( 
.A(n_1827),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_2110),
.Y(n_2283)
);

INVx6_ASAP7_75t_L g2284 ( 
.A(n_1882),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2017),
.Y(n_2285)
);

A2O1A1Ixp33_ASAP7_75t_L g2286 ( 
.A1(n_1936),
.A2(n_1816),
.B(n_1788),
.C(n_1876),
.Y(n_2286)
);

CKINVDCx11_ASAP7_75t_R g2287 ( 
.A(n_1948),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1834),
.B(n_606),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1905),
.B(n_609),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2027),
.A2(n_610),
.B(n_611),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2091),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1861),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2091),
.Y(n_2293)
);

INVx5_ASAP7_75t_L g2294 ( 
.A(n_1861),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2007),
.A2(n_613),
.B1(n_614),
.B2(n_616),
.Y(n_2295)
);

BUFx3_ASAP7_75t_L g2296 ( 
.A(n_1880),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2033),
.A2(n_617),
.B(n_619),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_1908),
.B(n_620),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_2088),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2092),
.Y(n_2300)
);

CKINVDCx11_ASAP7_75t_R g2301 ( 
.A(n_1948),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2092),
.Y(n_2302)
);

AO21x2_ASAP7_75t_L g2303 ( 
.A1(n_2112),
.A2(n_621),
.B(n_622),
.Y(n_2303)
);

BUFx2_ASAP7_75t_L g2304 ( 
.A(n_1835),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_1904),
.B(n_623),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_1851),
.Y(n_2306)
);

OAI21x1_ASAP7_75t_SL g2307 ( 
.A1(n_1816),
.A2(n_2056),
.B(n_2015),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_1851),
.Y(n_2308)
);

OAI22x1_ASAP7_75t_L g2309 ( 
.A1(n_1894),
.A2(n_627),
.B1(n_628),
.B2(n_629),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2093),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2093),
.Y(n_2311)
);

CKINVDCx20_ASAP7_75t_R g2312 ( 
.A(n_1882),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_1880),
.Y(n_2313)
);

OAI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2058),
.A2(n_631),
.B(n_632),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2007),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2121),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_1891),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_1924),
.B(n_633),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2018),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2121),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2018),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.Y(n_2321)
);

BUFx3_ASAP7_75t_L g2322 ( 
.A(n_1891),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_R g2323 ( 
.A(n_1954),
.B(n_637),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2061),
.A2(n_639),
.B(n_640),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_1927),
.B(n_639),
.Y(n_2325)
);

CKINVDCx20_ASAP7_75t_R g2326 ( 
.A(n_1995),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_1964),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_1913),
.B(n_640),
.Y(n_2328)
);

AO21x2_ASAP7_75t_L g2329 ( 
.A1(n_1781),
.A2(n_641),
.B(n_642),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1972),
.Y(n_2330)
);

INVx2_ASAP7_75t_SL g2331 ( 
.A(n_2068),
.Y(n_2331)
);

OAI21x1_ASAP7_75t_L g2332 ( 
.A1(n_1888),
.A2(n_642),
.B(n_643),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_1900),
.A2(n_644),
.B(n_645),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_1870),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1957),
.B(n_646),
.Y(n_2335)
);

OA21x2_ASAP7_75t_L g2336 ( 
.A1(n_1907),
.A2(n_646),
.B(n_647),
.Y(n_2336)
);

OR2x6_ASAP7_75t_L g2337 ( 
.A(n_2068),
.B(n_648),
.Y(n_2337)
);

AOI22x1_ASAP7_75t_L g2338 ( 
.A1(n_2064),
.A2(n_649),
.B1(n_650),
.B2(n_651),
.Y(n_2338)
);

AO21x2_ASAP7_75t_L g2339 ( 
.A1(n_2054),
.A2(n_652),
.B(n_653),
.Y(n_2339)
);

INVx6_ASAP7_75t_L g2340 ( 
.A(n_1972),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1870),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_2095),
.B(n_654),
.Y(n_2342)
);

AO21x2_ASAP7_75t_L g2343 ( 
.A1(n_2098),
.A2(n_655),
.B(n_656),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_1931),
.B(n_657),
.Y(n_2344)
);

NOR2x1_ASAP7_75t_SL g2345 ( 
.A(n_1938),
.B(n_657),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1961),
.B(n_658),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2134),
.Y(n_2347)
);

NOR2xp67_ASAP7_75t_L g2348 ( 
.A(n_1899),
.B(n_658),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_1982),
.B(n_659),
.Y(n_2349)
);

AO21x2_ASAP7_75t_L g2350 ( 
.A1(n_2111),
.A2(n_661),
.B(n_662),
.Y(n_2350)
);

NAND2x1p5_ASAP7_75t_L g2351 ( 
.A(n_2095),
.B(n_663),
.Y(n_2351)
);

NOR2xp67_ASAP7_75t_SL g2352 ( 
.A(n_1890),
.B(n_664),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_1985),
.B(n_666),
.Y(n_2353)
);

AO21x2_ASAP7_75t_L g2354 ( 
.A1(n_2129),
.A2(n_669),
.B(n_670),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_1940),
.B(n_669),
.Y(n_2355)
);

INVx5_ASAP7_75t_L g2356 ( 
.A(n_2099),
.Y(n_2356)
);

INVx4_ASAP7_75t_L g2357 ( 
.A(n_2069),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2119),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1822),
.B(n_671),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1944),
.B(n_671),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2071),
.A2(n_672),
.B(n_673),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_1895),
.B(n_673),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1944),
.B(n_674),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2045),
.B(n_675),
.Y(n_2364)
);

HB1xp67_ASAP7_75t_L g2365 ( 
.A(n_2119),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2073),
.A2(n_676),
.B(n_677),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_1895),
.B(n_678),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1944),
.B(n_679),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2134),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1802),
.Y(n_2370)
);

OAI21x1_ASAP7_75t_L g2371 ( 
.A1(n_1928),
.A2(n_681),
.B(n_682),
.Y(n_2371)
);

AO21x2_ASAP7_75t_L g2372 ( 
.A1(n_1856),
.A2(n_684),
.B(n_686),
.Y(n_2372)
);

AO21x2_ASAP7_75t_L g2373 ( 
.A1(n_1832),
.A2(n_684),
.B(n_687),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_1944),
.B(n_689),
.Y(n_2374)
);

OA21x2_ASAP7_75t_L g2375 ( 
.A1(n_2074),
.A2(n_689),
.B(n_690),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2138),
.B(n_691),
.Y(n_2376)
);

INVx4_ASAP7_75t_L g2377 ( 
.A(n_2069),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_1969),
.A2(n_692),
.B1(n_693),
.B2(n_694),
.Y(n_2378)
);

OR2x6_ASAP7_75t_L g2379 ( 
.A(n_2072),
.B(n_696),
.Y(n_2379)
);

OAI21x1_ASAP7_75t_L g2380 ( 
.A1(n_2075),
.A2(n_697),
.B(n_698),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_1982),
.B(n_697),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_2099),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_1871),
.Y(n_2383)
);

AOI22x1_ASAP7_75t_L g2384 ( 
.A1(n_2079),
.A2(n_702),
.B1(n_703),
.B2(n_704),
.Y(n_2384)
);

INVx2_ASAP7_75t_SL g2385 ( 
.A(n_2072),
.Y(n_2385)
);

OAI21x1_ASAP7_75t_L g2386 ( 
.A1(n_2082),
.A2(n_702),
.B(n_705),
.Y(n_2386)
);

INVx6_ASAP7_75t_L g2387 ( 
.A(n_1932),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1802),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_1865),
.B(n_705),
.Y(n_2389)
);

CKINVDCx14_ASAP7_75t_R g2390 ( 
.A(n_1938),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2048),
.Y(n_2391)
);

OAI21x1_ASAP7_75t_L g2392 ( 
.A1(n_2097),
.A2(n_710),
.B(n_711),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2049),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2078),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_2083),
.Y(n_2395)
);

BUFx5_ASAP7_75t_L g2396 ( 
.A(n_2104),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_SL g2397 ( 
.A(n_1956),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1801),
.Y(n_2398)
);

INVx6_ASAP7_75t_L g2399 ( 
.A(n_1932),
.Y(n_2399)
);

NAND2x1p5_ASAP7_75t_L g2400 ( 
.A(n_2105),
.B(n_713),
.Y(n_2400)
);

INVx3_ASAP7_75t_SL g2401 ( 
.A(n_1938),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1801),
.Y(n_2402)
);

NOR2x1_ASAP7_75t_R g2403 ( 
.A(n_1933),
.B(n_714),
.Y(n_2403)
);

AND2x6_ASAP7_75t_L g2404 ( 
.A(n_2105),
.B(n_1951),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_1965),
.A2(n_715),
.B1(n_716),
.B2(n_717),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_1843),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1944),
.B(n_719),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_1921),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_1826),
.Y(n_2409)
);

AO21x1_ASAP7_75t_L g2410 ( 
.A1(n_2138),
.A2(n_720),
.B(n_721),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2077),
.Y(n_2411)
);

OAI21x1_ASAP7_75t_SL g2412 ( 
.A1(n_1860),
.A2(n_722),
.B(n_723),
.Y(n_2412)
);

AOI21xp33_ASAP7_75t_L g2413 ( 
.A1(n_1805),
.A2(n_724),
.B(n_725),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_1973),
.B(n_725),
.Y(n_2414)
);

CKINVDCx20_ASAP7_75t_R g2415 ( 
.A(n_1983),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2115),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2115),
.Y(n_2417)
);

INVx5_ASAP7_75t_SL g2418 ( 
.A(n_1871),
.Y(n_2418)
);

OA21x2_ASAP7_75t_L g2419 ( 
.A1(n_2012),
.A2(n_728),
.B(n_729),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_1871),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1973),
.B(n_729),
.Y(n_2421)
);

AO21x2_ASAP7_75t_L g2422 ( 
.A1(n_1975),
.A2(n_730),
.B(n_731),
.Y(n_2422)
);

AO31x2_ASAP7_75t_L g2423 ( 
.A1(n_1841),
.A2(n_730),
.A3(n_732),
.B(n_733),
.Y(n_2423)
);

AO21x2_ASAP7_75t_L g2424 ( 
.A1(n_1975),
.A2(n_732),
.B(n_733),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_1933),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2030),
.Y(n_2426)
);

OAI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_1958),
.A2(n_736),
.B(n_737),
.Y(n_2427)
);

OAI21x1_ASAP7_75t_L g2428 ( 
.A1(n_1978),
.A2(n_738),
.B(n_739),
.Y(n_2428)
);

AOI22x1_ASAP7_75t_L g2429 ( 
.A1(n_1786),
.A2(n_741),
.B1(n_742),
.B2(n_743),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2042),
.B(n_741),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2043),
.Y(n_2431)
);

AOI22xp33_ASAP7_75t_L g2432 ( 
.A1(n_2000),
.A2(n_742),
.B1(n_743),
.B2(n_744),
.Y(n_2432)
);

AO21x1_ASAP7_75t_L g2433 ( 
.A1(n_1910),
.A2(n_746),
.B(n_747),
.Y(n_2433)
);

BUFx12f_ASAP7_75t_L g2434 ( 
.A(n_1979),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_1939),
.A2(n_747),
.B(n_750),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_1958),
.A2(n_751),
.B(n_752),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_1912),
.A2(n_753),
.B(n_754),
.Y(n_2437)
);

OAI21x1_ASAP7_75t_L g2438 ( 
.A1(n_1916),
.A2(n_754),
.B(n_755),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_1966),
.A2(n_755),
.B(n_756),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_1925),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_1937),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1874),
.Y(n_2442)
);

AO21x2_ASAP7_75t_L g2443 ( 
.A1(n_2096),
.A2(n_762),
.B(n_763),
.Y(n_2443)
);

AOI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2000),
.A2(n_764),
.B1(n_765),
.B2(n_766),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2044),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2052),
.Y(n_2446)
);

NOR2x1_ASAP7_75t_R g2447 ( 
.A(n_1937),
.B(n_765),
.Y(n_2447)
);

NAND2x1p5_ASAP7_75t_L g2448 ( 
.A(n_1887),
.B(n_766),
.Y(n_2448)
);

AO21x2_ASAP7_75t_L g2449 ( 
.A1(n_2100),
.A2(n_767),
.B(n_768),
.Y(n_2449)
);

OAI21x1_ASAP7_75t_SL g2450 ( 
.A1(n_1876),
.A2(n_767),
.B(n_770),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_1925),
.B(n_770),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_1867),
.B(n_771),
.Y(n_2452)
);

O2A1O1Ixp33_ASAP7_75t_L g2453 ( 
.A1(n_1878),
.A2(n_777),
.B(n_772),
.C(n_775),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_1997),
.B(n_771),
.Y(n_2454)
);

BUFx2_ASAP7_75t_R g2455 ( 
.A(n_1881),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2059),
.Y(n_2456)
);

INVx8_ASAP7_75t_L g2457 ( 
.A(n_1986),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2060),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_1986),
.B(n_772),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2062),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_1966),
.A2(n_1824),
.B(n_2005),
.Y(n_2461)
);

OAI21x1_ASAP7_75t_SL g2462 ( 
.A1(n_1999),
.A2(n_1911),
.B(n_1915),
.Y(n_2462)
);

OAI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_1915),
.A2(n_1809),
.B1(n_1999),
.B2(n_2137),
.Y(n_2463)
);

OA21x2_ASAP7_75t_L g2464 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1971),
.Y(n_2464)
);

AO21x2_ASAP7_75t_L g2465 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1971),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2085),
.B(n_1926),
.Y(n_2466)
);

CKINVDCx14_ASAP7_75t_R g2467 ( 
.A(n_2137),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_1986),
.B(n_2065),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_1911),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2102),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2467),
.A2(n_2127),
.B1(n_1963),
.B2(n_2039),
.Y(n_2471)
);

AOI21x1_ASAP7_75t_L g2472 ( 
.A1(n_2162),
.A2(n_1854),
.B(n_1872),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2171),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2181),
.B(n_1796),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_2145),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2141),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2467),
.A2(n_2127),
.B1(n_1963),
.B2(n_2039),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2140),
.Y(n_2478)
);

BUFx4f_ASAP7_75t_SL g2479 ( 
.A(n_2255),
.Y(n_2479)
);

BUFx8_ASAP7_75t_SL g2480 ( 
.A(n_2153),
.Y(n_2480)
);

INVx3_ASAP7_75t_L g2481 ( 
.A(n_2171),
.Y(n_2481)
);

INVx2_ASAP7_75t_SL g2482 ( 
.A(n_2145),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2149),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2152),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2139),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2173),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2409),
.Y(n_2487)
);

AO21x2_ASAP7_75t_L g2488 ( 
.A1(n_2184),
.A2(n_1943),
.B(n_1945),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2183),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2409),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2234),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2189),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2170),
.B(n_1962),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2234),
.Y(n_2494)
);

HB1xp67_ASAP7_75t_L g2495 ( 
.A(n_2170),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2163),
.B(n_1990),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2442),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2210),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2218),
.Y(n_2499)
);

AOI22xp33_ASAP7_75t_L g2500 ( 
.A1(n_2229),
.A2(n_2250),
.B1(n_2249),
.B2(n_2287),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2230),
.Y(n_2501)
);

BUFx3_ASAP7_75t_L g2502 ( 
.A(n_2140),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2196),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2196),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2199),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2199),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2163),
.B(n_1784),
.Y(n_2507)
);

AO21x2_ASAP7_75t_L g2508 ( 
.A1(n_2462),
.A2(n_1883),
.B(n_1864),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_L g2509 ( 
.A1(n_2229),
.A2(n_2128),
.B1(n_1886),
.B2(n_2124),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2208),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2208),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2163),
.B(n_2011),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2235),
.Y(n_2513)
);

HB1xp67_ASAP7_75t_L g2514 ( 
.A(n_2315),
.Y(n_2514)
);

AO21x1_ASAP7_75t_SL g2515 ( 
.A1(n_2411),
.A2(n_1896),
.B(n_1918),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2189),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2235),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2229),
.A2(n_1794),
.B1(n_1949),
.B2(n_1830),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2288),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2180),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2249),
.A2(n_1794),
.B1(n_1993),
.B2(n_1935),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2164),
.B(n_2108),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2288),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2160),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2164),
.B(n_1849),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2236),
.B(n_2106),
.Y(n_2526)
);

OA21x2_ASAP7_75t_L g2527 ( 
.A1(n_2172),
.A2(n_1892),
.B(n_1941),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2299),
.B(n_1804),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2179),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2232),
.Y(n_2530)
);

OA21x2_ASAP7_75t_L g2531 ( 
.A1(n_2172),
.A2(n_1892),
.B(n_1941),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2160),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2249),
.A2(n_1920),
.B1(n_1898),
.B2(n_1955),
.Y(n_2533)
);

BUFx2_ASAP7_75t_L g2534 ( 
.A(n_2180),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2232),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2158),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2315),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2179),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2358),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2158),
.Y(n_2540)
);

BUFx2_ASAP7_75t_R g2541 ( 
.A(n_2153),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2250),
.A2(n_1993),
.B1(n_1935),
.B2(n_1910),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2359),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2359),
.Y(n_2544)
);

INVx2_ASAP7_75t_SL g2545 ( 
.A(n_2284),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2335),
.Y(n_2546)
);

NAND2x1_ASAP7_75t_L g2547 ( 
.A(n_2404),
.B(n_1852),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2335),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2358),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2346),
.Y(n_2550)
);

INVx1_ASAP7_75t_SL g2551 ( 
.A(n_2186),
.Y(n_2551)
);

AOI221xp5_ASAP7_75t_L g2552 ( 
.A1(n_2247),
.A2(n_1885),
.B1(n_1866),
.B2(n_1920),
.C(n_2067),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2164),
.B(n_1934),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2346),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_2180),
.Y(n_2555)
);

HB1xp67_ASAP7_75t_L g2556 ( 
.A(n_2365),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2198),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2365),
.Y(n_2558)
);

INVx3_ASAP7_75t_L g2559 ( 
.A(n_2198),
.Y(n_2559)
);

AOI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2390),
.A2(n_1981),
.B1(n_1909),
.B2(n_1994),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2147),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2203),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2203),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2147),
.Y(n_2564)
);

OAI21xp5_ASAP7_75t_L g2565 ( 
.A1(n_2286),
.A2(n_1825),
.B(n_1842),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2206),
.Y(n_2566)
);

CKINVDCx11_ASAP7_75t_R g2567 ( 
.A(n_2200),
.Y(n_2567)
);

BUFx12f_ASAP7_75t_L g2568 ( 
.A(n_2200),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2204),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2204),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2207),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2207),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_SL g2573 ( 
.A1(n_2390),
.A2(n_1866),
.B1(n_1885),
.B2(n_1988),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2212),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2175),
.B(n_1994),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2206),
.Y(n_2576)
);

INVx6_ASAP7_75t_L g2577 ( 
.A(n_2294),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2250),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2212),
.Y(n_2579)
);

INVx3_ASAP7_75t_L g2580 ( 
.A(n_2357),
.Y(n_2580)
);

AO21x2_ASAP7_75t_L g2581 ( 
.A1(n_2286),
.A2(n_1896),
.B(n_1988),
.Y(n_2581)
);

NAND2x1p5_ASAP7_75t_L g2582 ( 
.A(n_2357),
.B(n_1793),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2214),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2337),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2214),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2287),
.A2(n_1968),
.B1(n_1909),
.B2(n_1903),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2301),
.A2(n_1903),
.B1(n_1992),
.B2(n_1980),
.Y(n_2587)
);

BUFx5_ASAP7_75t_L g2588 ( 
.A(n_2404),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2301),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2277),
.Y(n_2590)
);

BUFx2_ASAP7_75t_L g2591 ( 
.A(n_2143),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2277),
.Y(n_2592)
);

BUFx2_ASAP7_75t_L g2593 ( 
.A(n_2143),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2178),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2289),
.Y(n_2595)
);

BUFx10_ASAP7_75t_L g2596 ( 
.A(n_2284),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_2186),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2466),
.B(n_1884),
.Y(n_2598)
);

OR2x6_ASAP7_75t_L g2599 ( 
.A(n_2175),
.B(n_2337),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2150),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2175),
.A2(n_1992),
.B1(n_1974),
.B2(n_1946),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2289),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2451),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2451),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2463),
.A2(n_1825),
.B(n_1842),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2463),
.A2(n_2166),
.B(n_2461),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2258),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2377),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2258),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2205),
.A2(n_2050),
.B1(n_2125),
.B2(n_1952),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2264),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2264),
.Y(n_2612)
);

INVx3_ASAP7_75t_SL g2613 ( 
.A(n_2225),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2169),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2169),
.Y(n_2615)
);

BUFx4f_ASAP7_75t_SL g2616 ( 
.A(n_2167),
.Y(n_2616)
);

HB1xp67_ASAP7_75t_L g2617 ( 
.A(n_2337),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2223),
.B(n_1998),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2226),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2379),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2379),
.Y(n_2621)
);

NOR2x1_ASAP7_75t_L g2622 ( 
.A(n_2379),
.B(n_2026),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2155),
.Y(n_2623)
);

AO21x1_ASAP7_75t_SL g2624 ( 
.A1(n_2411),
.A2(n_1833),
.B(n_1831),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2273),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2265),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2265),
.Y(n_2627)
);

BUFx12f_ASAP7_75t_L g2628 ( 
.A(n_2272),
.Y(n_2628)
);

INVx1_ASAP7_75t_SL g2629 ( 
.A(n_2245),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2273),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2351),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2351),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2148),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2273),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2243),
.Y(n_2635)
);

BUFx2_ASAP7_75t_L g2636 ( 
.A(n_2150),
.Y(n_2636)
);

INVx4_ASAP7_75t_SL g2637 ( 
.A(n_2401),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2148),
.Y(n_2638)
);

AOI21x1_ASAP7_75t_L g2639 ( 
.A1(n_2469),
.A2(n_1847),
.B(n_1929),
.Y(n_2639)
);

OR2x6_ASAP7_75t_L g2640 ( 
.A(n_2342),
.B(n_1923),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2240),
.B(n_2109),
.Y(n_2641)
);

INVx2_ASAP7_75t_SL g2642 ( 
.A(n_2284),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2233),
.Y(n_2643)
);

OR2x6_ASAP7_75t_L g2644 ( 
.A(n_2342),
.B(n_2014),
.Y(n_2644)
);

BUFx3_ASAP7_75t_L g2645 ( 
.A(n_2182),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2355),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2355),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2253),
.Y(n_2648)
);

AOI21x1_ASAP7_75t_L g2649 ( 
.A1(n_2469),
.A2(n_1813),
.B(n_1950),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2253),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2142),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2190),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_2342),
.B(n_1906),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2254),
.B(n_2107),
.Y(n_2654)
);

INVx2_ASAP7_75t_SL g2655 ( 
.A(n_2387),
.Y(n_2655)
);

BUFx2_ASAP7_75t_L g2656 ( 
.A(n_2182),
.Y(n_2656)
);

OAI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2144),
.A2(n_1848),
.B(n_1828),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2362),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2205),
.A2(n_2135),
.B1(n_2094),
.B2(n_1848),
.Y(n_2659)
);

OR2x2_ASAP7_75t_L g2660 ( 
.A(n_2299),
.B(n_2245),
.Y(n_2660)
);

CKINVDCx20_ASAP7_75t_R g2661 ( 
.A(n_2312),
.Y(n_2661)
);

AO21x2_ASAP7_75t_L g2662 ( 
.A1(n_2157),
.A2(n_1879),
.B(n_1960),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_L g2663 ( 
.A1(n_2433),
.A2(n_1828),
.B1(n_1829),
.B2(n_1831),
.Y(n_2663)
);

OAI21x1_ASAP7_75t_SL g2664 ( 
.A1(n_2345),
.A2(n_1922),
.B(n_1930),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2362),
.Y(n_2665)
);

BUFx3_ASAP7_75t_L g2666 ( 
.A(n_2197),
.Y(n_2666)
);

OR2x6_ASAP7_75t_L g2667 ( 
.A(n_2262),
.B(n_2021),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2367),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2367),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2321),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2321),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2294),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2197),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2459),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2223),
.B(n_1998),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2459),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2174),
.Y(n_2677)
);

HB1xp67_ASAP7_75t_L g2678 ( 
.A(n_2294),
.Y(n_2678)
);

OR2x6_ASAP7_75t_L g2679 ( 
.A(n_2377),
.B(n_2122),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2174),
.Y(n_2680)
);

OAI21xp5_ASAP7_75t_L g2681 ( 
.A1(n_2144),
.A2(n_1829),
.B(n_1897),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2305),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2305),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2425),
.B(n_2306),
.Y(n_2684)
);

INVx1_ASAP7_75t_SL g2685 ( 
.A(n_2267),
.Y(n_2685)
);

BUFx2_ASAP7_75t_L g2686 ( 
.A(n_2420),
.Y(n_2686)
);

INVx1_ASAP7_75t_SL g2687 ( 
.A(n_2267),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2344),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2239),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2364),
.Y(n_2690)
);

OR2x6_ASAP7_75t_L g2691 ( 
.A(n_2201),
.B(n_2029),
.Y(n_2691)
);

INVxp33_ASAP7_75t_L g2692 ( 
.A(n_2403),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2238),
.B(n_1984),
.Y(n_2693)
);

BUFx2_ASAP7_75t_L g2694 ( 
.A(n_2420),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2308),
.B(n_2114),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2364),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2448),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2294),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2448),
.Y(n_2699)
);

OAI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2401),
.A2(n_1976),
.B1(n_1897),
.B2(n_1836),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2241),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2356),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2241),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2423),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2423),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_2408),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2387),
.Y(n_2707)
);

INVx2_ASAP7_75t_SL g2708 ( 
.A(n_2387),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2408),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2348),
.Y(n_2710)
);

INVxp67_ASAP7_75t_L g2711 ( 
.A(n_2376),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2391),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2393),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2142),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2223),
.B(n_1998),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2242),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2399),
.Y(n_2717)
);

OR2x2_ASAP7_75t_SL g2718 ( 
.A(n_2399),
.B(n_2089),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2394),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2414),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2268),
.B(n_1914),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2247),
.A2(n_2032),
.B1(n_1919),
.B2(n_1989),
.Y(n_2722)
);

OAI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2221),
.A2(n_1996),
.B(n_1998),
.Y(n_2723)
);

BUFx12f_ASAP7_75t_L g2724 ( 
.A(n_2272),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2414),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2421),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2389),
.B(n_2130),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2421),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2239),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2261),
.Y(n_2730)
);

CKINVDCx14_ASAP7_75t_R g2731 ( 
.A(n_2312),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2261),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2356),
.Y(n_2733)
);

NAND2x1p5_ASAP7_75t_L g2734 ( 
.A(n_2356),
.B(n_1914),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2298),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2282),
.B(n_2113),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2257),
.A2(n_1782),
.B1(n_2008),
.B2(n_2013),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2239),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2298),
.Y(n_2739)
);

BUFx2_ASAP7_75t_L g2740 ( 
.A(n_2213),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2328),
.Y(n_2741)
);

BUFx4f_ASAP7_75t_SL g2742 ( 
.A(n_2228),
.Y(n_2742)
);

OAI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2221),
.A2(n_1953),
.B(n_1782),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2328),
.Y(n_2744)
);

OAI22x1_ASAP7_75t_L g2745 ( 
.A1(n_2151),
.A2(n_2222),
.B1(n_2256),
.B2(n_2406),
.Y(n_2745)
);

OR2x6_ASAP7_75t_L g2746 ( 
.A(n_2331),
.B(n_1782),
.Y(n_2746)
);

OAI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2295),
.A2(n_2008),
.B1(n_2013),
.B2(n_2113),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2349),
.Y(n_2748)
);

INVx2_ASAP7_75t_SL g2749 ( 
.A(n_2399),
.Y(n_2749)
);

OAI21x1_ASAP7_75t_L g2750 ( 
.A1(n_2292),
.A2(n_1959),
.B(n_1953),
.Y(n_2750)
);

OAI21x1_ASAP7_75t_L g2751 ( 
.A1(n_2341),
.A2(n_1959),
.B(n_1953),
.Y(n_2751)
);

AO21x2_ASAP7_75t_L g2752 ( 
.A1(n_2188),
.A2(n_2008),
.B(n_2013),
.Y(n_2752)
);

AOI22xp33_ASAP7_75t_L g2753 ( 
.A1(n_2257),
.A2(n_2113),
.B1(n_1991),
.B2(n_1959),
.Y(n_2753)
);

AOI22xp33_ASAP7_75t_SL g2754 ( 
.A1(n_2257),
.A2(n_2441),
.B1(n_2418),
.B2(n_2307),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2356),
.Y(n_2755)
);

OAI222xp33_ASAP7_75t_L g2756 ( 
.A1(n_2319),
.A2(n_1991),
.B1(n_2352),
.B2(n_2260),
.C1(n_2237),
.C2(n_2378),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2340),
.Y(n_2757)
);

AOI22xp33_ASAP7_75t_SL g2758 ( 
.A1(n_2418),
.A2(n_2326),
.B1(n_2217),
.B2(n_2270),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2381),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2416),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2476),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2479),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2483),
.Y(n_2763)
);

INVxp67_ASAP7_75t_SL g2764 ( 
.A(n_2524),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2660),
.B(n_2551),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2551),
.B(n_2395),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2474),
.B(n_2318),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2484),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2495),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_SL g2770 ( 
.A1(n_2584),
.A2(n_2418),
.B1(n_2326),
.B2(n_2383),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2493),
.B(n_2325),
.Y(n_2771)
);

OAI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2500),
.A2(n_2395),
.B1(n_2464),
.B2(n_2444),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2643),
.B(n_2452),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_L g2774 ( 
.A1(n_2542),
.A2(n_2146),
.B1(n_2454),
.B2(n_2396),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2692),
.B(n_2406),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2652),
.B(n_2353),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2597),
.B(n_2246),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_SL g2778 ( 
.A1(n_2584),
.A2(n_2266),
.B1(n_2464),
.B2(n_2336),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2597),
.B(n_2440),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2629),
.B(n_2500),
.Y(n_2780)
);

INVxp67_ASAP7_75t_SL g2781 ( 
.A(n_2524),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2577),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2670),
.B(n_2370),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2629),
.B(n_2246),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2637),
.B(n_2248),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2671),
.B(n_2388),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2486),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2594),
.B(n_2309),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2495),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2514),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2740),
.B(n_2440),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2489),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2514),
.Y(n_2793)
);

HB1xp67_ASAP7_75t_L g2794 ( 
.A(n_2537),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2498),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2507),
.B(n_2454),
.Y(n_2796)
);

HB1xp67_ASAP7_75t_L g2797 ( 
.A(n_2537),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2499),
.Y(n_2798)
);

INVxp67_ASAP7_75t_SL g2799 ( 
.A(n_2532),
.Y(n_2799)
);

BUFx2_ASAP7_75t_L g2800 ( 
.A(n_2599),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2637),
.B(n_2599),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2512),
.B(n_2248),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2539),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2491),
.B(n_2398),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2501),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2522),
.B(n_2417),
.Y(n_2806)
);

INVxp67_ASAP7_75t_L g2807 ( 
.A(n_2624),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2712),
.B(n_2146),
.Y(n_2808)
);

NOR2x1_ASAP7_75t_SL g2809 ( 
.A(n_2599),
.B(n_2385),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2494),
.B(n_2402),
.Y(n_2810)
);

INVx4_ASAP7_75t_R g2811 ( 
.A(n_2475),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2487),
.Y(n_2812)
);

BUFx2_ASAP7_75t_L g2813 ( 
.A(n_2561),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2487),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2542),
.A2(n_2396),
.B1(n_2276),
.B2(n_2279),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2713),
.B(n_2427),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2692),
.B(n_2219),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2719),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2760),
.Y(n_2819)
);

HB1xp67_ASAP7_75t_L g2820 ( 
.A(n_2539),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2479),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2706),
.B(n_2427),
.Y(n_2822)
);

AOI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2533),
.A2(n_2396),
.B1(n_2347),
.B2(n_2280),
.Y(n_2823)
);

INVx2_ASAP7_75t_SL g2824 ( 
.A(n_2596),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2709),
.B(n_2360),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2637),
.B(n_2330),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2620),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2490),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2549),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2621),
.Y(n_2830)
);

AOI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2509),
.A2(n_2251),
.B1(n_2369),
.B2(n_2320),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2521),
.A2(n_2432),
.B1(n_2444),
.B2(n_2259),
.Y(n_2832)
);

BUFx2_ASAP7_75t_L g2833 ( 
.A(n_2566),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2684),
.B(n_2436),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2623),
.B(n_2436),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2533),
.A2(n_2396),
.B1(n_2278),
.B2(n_2302),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2748),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2759),
.Y(n_2838)
);

AOI22xp33_ASAP7_75t_L g2839 ( 
.A1(n_2573),
.A2(n_2396),
.B1(n_2285),
.B2(n_2291),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2509),
.A2(n_2521),
.B1(n_2573),
.B2(n_2552),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2736),
.Y(n_2841)
);

INVxp67_ASAP7_75t_SL g2842 ( 
.A(n_2532),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2553),
.B(n_2439),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2577),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2653),
.B(n_2439),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2727),
.B(n_2293),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2720),
.B(n_2300),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2575),
.B(n_2432),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2577),
.Y(n_2849)
);

OR2x6_ASAP7_75t_L g2850 ( 
.A(n_2640),
.B(n_2400),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2496),
.B(n_2405),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2690),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2696),
.Y(n_2853)
);

BUFx3_ASAP7_75t_L g2854 ( 
.A(n_2661),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2655),
.B(n_2373),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2707),
.B(n_2373),
.Y(n_2856)
);

INVx2_ASAP7_75t_SL g2857 ( 
.A(n_2596),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2549),
.Y(n_2858)
);

BUFx3_ASAP7_75t_L g2859 ( 
.A(n_2661),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2725),
.B(n_2310),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2471),
.A2(n_2161),
.B1(n_2275),
.B2(n_2216),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2480),
.Y(n_2862)
);

OAI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2471),
.A2(n_2202),
.B1(n_2209),
.B2(n_2192),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2708),
.B(n_2426),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2617),
.B(n_2363),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2717),
.B(n_2431),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2556),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2617),
.B(n_2368),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2580),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2749),
.B(n_2445),
.Y(n_2870)
);

AOI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2552),
.A2(n_2396),
.B1(n_2316),
.B2(n_2311),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2497),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2614),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2686),
.B(n_2446),
.Y(n_2874)
);

AOI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2644),
.A2(n_2410),
.B1(n_2458),
.B2(n_2456),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2694),
.B(n_2578),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2615),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2480),
.Y(n_2878)
);

AND2x4_ASAP7_75t_L g2879 ( 
.A(n_2473),
.B(n_2330),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2726),
.B(n_2465),
.Y(n_2880)
);

OAI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2477),
.A2(n_2177),
.B1(n_2202),
.B2(n_2216),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2728),
.B(n_2465),
.Y(n_2882)
);

OR2x2_ASAP7_75t_L g2883 ( 
.A(n_2578),
.B(n_2368),
.Y(n_2883)
);

AOI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2644),
.A2(n_2470),
.B1(n_2460),
.B2(n_2215),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2591),
.B(n_2372),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2485),
.B(n_2323),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2593),
.B(n_2372),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2600),
.B(n_2468),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2644),
.A2(n_2468),
.B1(n_2429),
.B2(n_2413),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2503),
.B(n_2374),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2556),
.Y(n_2891)
);

AOI22xp33_ASAP7_75t_L g2892 ( 
.A1(n_2477),
.A2(n_2215),
.B1(n_2165),
.B2(n_2168),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2558),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2504),
.B(n_2374),
.Y(n_2894)
);

INVxp67_ASAP7_75t_L g2895 ( 
.A(n_2515),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2558),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2505),
.B(n_2407),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2626),
.Y(n_2898)
);

OAI21xp33_ASAP7_75t_SL g2899 ( 
.A1(n_2640),
.A2(n_2407),
.B(n_2191),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2627),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2750),
.Y(n_2901)
);

CKINVDCx14_ASAP7_75t_R g2902 ( 
.A(n_2731),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2631),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_2473),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2632),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2506),
.B(n_2165),
.Y(n_2906)
);

OAI21xp33_ASAP7_75t_L g2907 ( 
.A1(n_2737),
.A2(n_2297),
.B(n_2290),
.Y(n_2907)
);

BUFx4f_ASAP7_75t_SL g2908 ( 
.A(n_2568),
.Y(n_2908)
);

NAND2x1_ASAP7_75t_L g2909 ( 
.A(n_2580),
.B(n_2404),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2633),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2638),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2510),
.B(n_2511),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2562),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2636),
.B(n_2296),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2563),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2656),
.B(n_2296),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2569),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2567),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2672),
.Y(n_2919)
);

INVx3_ASAP7_75t_L g2920 ( 
.A(n_2481),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2613),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2481),
.Y(n_2922)
);

INVx3_ASAP7_75t_L g2923 ( 
.A(n_2492),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2730),
.B(n_2322),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2598),
.A2(n_2415),
.B1(n_2430),
.B2(n_2227),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2570),
.Y(n_2926)
);

BUFx2_ASAP7_75t_L g2927 ( 
.A(n_2672),
.Y(n_2927)
);

AND2x4_ASAP7_75t_SL g2928 ( 
.A(n_2482),
.B(n_2608),
.Y(n_2928)
);

HB1xp67_ASAP7_75t_L g2929 ( 
.A(n_2751),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2732),
.B(n_2322),
.Y(n_2930)
);

AND2x4_ASAP7_75t_L g2931 ( 
.A(n_2492),
.B(n_2334),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2571),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2613),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2572),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2513),
.B(n_2168),
.Y(n_2935)
);

INVxp67_ASAP7_75t_SL g2936 ( 
.A(n_2635),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2598),
.A2(n_2176),
.B1(n_2422),
.B2(n_2424),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2574),
.Y(n_2938)
);

AOI222xp33_ASAP7_75t_L g2939 ( 
.A1(n_2701),
.A2(n_2447),
.B1(n_2195),
.B2(n_2227),
.C1(n_2361),
.C2(n_2366),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2579),
.Y(n_2940)
);

BUFx2_ASAP7_75t_L g2941 ( 
.A(n_2678),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2703),
.B(n_2693),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2583),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2528),
.B(n_2413),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2585),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2607),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2609),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2586),
.A2(n_2587),
.B1(n_2518),
.B2(n_2640),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2611),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2612),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2678),
.Y(n_2951)
);

NAND2x1p5_ASAP7_75t_L g2952 ( 
.A(n_2608),
.B(n_2334),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2698),
.Y(n_2953)
);

HB1xp67_ASAP7_75t_L g2954 ( 
.A(n_2734),
.Y(n_2954)
);

BUFx4f_ASAP7_75t_L g2955 ( 
.A(n_2628),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2698),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2517),
.B(n_2176),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2702),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2519),
.B(n_2220),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2516),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2689),
.B(n_2327),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2586),
.A2(n_2252),
.B1(n_2384),
.B2(n_2338),
.Y(n_2962)
);

AOI22xp33_ASAP7_75t_L g2963 ( 
.A1(n_2587),
.A2(n_2193),
.B1(n_2412),
.B2(n_2450),
.Y(n_2963)
);

INVx1_ASAP7_75t_SL g2964 ( 
.A(n_2702),
.Y(n_2964)
);

AND2x4_ASAP7_75t_L g2965 ( 
.A(n_2516),
.B(n_2382),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2733),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2645),
.B(n_2666),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2689),
.B(n_2327),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2478),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2757),
.B(n_2658),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2755),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2478),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2757),
.B(n_2271),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2595),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2502),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2665),
.B(n_2271),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2602),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2536),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2668),
.B(n_2283),
.Y(n_2979)
);

INVx4_ASAP7_75t_R g2980 ( 
.A(n_2731),
.Y(n_2980)
);

HB1xp67_ASAP7_75t_L g2981 ( 
.A(n_2734),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2540),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2523),
.B(n_2422),
.Y(n_2983)
);

BUFx3_ASAP7_75t_L g2984 ( 
.A(n_2742),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2710),
.Y(n_2985)
);

OAI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2560),
.A2(n_2177),
.B1(n_2209),
.B2(n_2192),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2546),
.B(n_2424),
.Y(n_2987)
);

BUFx2_ASAP7_75t_L g2988 ( 
.A(n_2502),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2669),
.B(n_2564),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2567),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2603),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2564),
.B(n_2283),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2604),
.Y(n_2993)
);

INVx5_ASAP7_75t_L g2994 ( 
.A(n_2716),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2646),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2635),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2647),
.Y(n_2997)
);

INVx4_ASAP7_75t_L g2998 ( 
.A(n_2576),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2576),
.B(n_2313),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2525),
.B(n_2695),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2548),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2550),
.Y(n_3002)
);

INVx4_ASAP7_75t_L g3003 ( 
.A(n_2666),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2554),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2685),
.B(n_2304),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2673),
.B(n_2313),
.Y(n_3006)
);

INVx3_ASAP7_75t_L g3007 ( 
.A(n_2673),
.Y(n_3007)
);

BUFx3_ASAP7_75t_L g3008 ( 
.A(n_2742),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2685),
.B(n_2317),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2687),
.B(n_2317),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2687),
.B(n_2329),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2729),
.B(n_2329),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2590),
.B(n_2592),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_2616),
.Y(n_3014)
);

OAI222xp33_ASAP7_75t_L g3015 ( 
.A1(n_2758),
.A2(n_2260),
.B1(n_2237),
.B2(n_2435),
.C1(n_2400),
.C2(n_2453),
.Y(n_3015)
);

INVx1_ASAP7_75t_SL g3016 ( 
.A(n_2557),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2729),
.B(n_2339),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2738),
.B(n_2339),
.Y(n_3018)
);

INVx3_ASAP7_75t_L g3019 ( 
.A(n_2618),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2648),
.Y(n_3020)
);

OR2x2_ASAP7_75t_L g3021 ( 
.A(n_2520),
.B(n_2534),
.Y(n_3021)
);

INVx3_ASAP7_75t_L g3022 ( 
.A(n_2618),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_2650),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2682),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2518),
.A2(n_2663),
.B1(n_2601),
.B2(n_2610),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2529),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2683),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2738),
.B(n_2343),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2735),
.B(n_2343),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_2555),
.B(n_2457),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2688),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2610),
.A2(n_2193),
.B1(n_2361),
.B2(n_2297),
.Y(n_3032)
);

OR2x2_ASAP7_75t_L g3033 ( 
.A(n_2543),
.B(n_2457),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2761),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_3000),
.B(n_2746),
.Y(n_3035)
);

NAND3xp33_ASAP7_75t_L g3036 ( 
.A(n_2840),
.B(n_2737),
.C(n_2753),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2763),
.Y(n_3037)
);

HB1xp67_ASAP7_75t_L g3038 ( 
.A(n_2790),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2771),
.B(n_2806),
.Y(n_3039)
);

BUFx2_ASAP7_75t_SL g3040 ( 
.A(n_2984),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2768),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2787),
.Y(n_3042)
);

HB1xp67_ASAP7_75t_L g3043 ( 
.A(n_2790),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2792),
.Y(n_3044)
);

OAI222xp33_ASAP7_75t_L g3045 ( 
.A1(n_2948),
.A2(n_2754),
.B1(n_2758),
.B2(n_2746),
.C1(n_2711),
.C2(n_2622),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2840),
.A2(n_2739),
.B1(n_2744),
.B2(n_2741),
.Y(n_3046)
);

HB1xp67_ASAP7_75t_L g3047 ( 
.A(n_2793),
.Y(n_3047)
);

BUFx2_ASAP7_75t_L g3048 ( 
.A(n_2869),
.Y(n_3048)
);

NOR2xp67_ASAP7_75t_SL g3049 ( 
.A(n_2762),
.B(n_2589),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2942),
.B(n_2746),
.Y(n_3050)
);

OR2x2_ASAP7_75t_L g3051 ( 
.A(n_2765),
.B(n_2721),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2795),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2798),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2805),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2818),
.Y(n_3055)
);

BUFx3_ASAP7_75t_L g3056 ( 
.A(n_3008),
.Y(n_3056)
);

INVxp67_ASAP7_75t_L g3057 ( 
.A(n_2919),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_SL g3058 ( 
.A(n_2807),
.B(n_2541),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2807),
.B(n_2675),
.Y(n_3059)
);

OR2x2_ASAP7_75t_L g3060 ( 
.A(n_2766),
.B(n_2721),
.Y(n_3060)
);

OAI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_2832),
.A2(n_2700),
.B1(n_2679),
.B2(n_2680),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_SL g3062 ( 
.A1(n_2948),
.A2(n_2677),
.B1(n_2606),
.B2(n_2508),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_2767),
.B(n_2674),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2819),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2837),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2838),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_3001),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_3029),
.B(n_2704),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_3014),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3002),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2796),
.B(n_2676),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3004),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2978),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_2869),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2802),
.B(n_2488),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2939),
.A2(n_2700),
.B1(n_2659),
.B2(n_2544),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2783),
.B(n_2786),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2982),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2812),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2854),
.B(n_2859),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2841),
.B(n_2705),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2880),
.B(n_2605),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2846),
.B(n_2530),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2895),
.B(n_2754),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2876),
.B(n_2488),
.Y(n_3085)
);

INVxp67_ASAP7_75t_L g3086 ( 
.A(n_2927),
.Y(n_3086)
);

BUFx2_ASAP7_75t_L g3087 ( 
.A(n_3003),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2912),
.Y(n_3088)
);

AOI22xp33_ASAP7_75t_L g3089 ( 
.A1(n_2939),
.A2(n_2659),
.B1(n_2745),
.B2(n_2535),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2912),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3013),
.Y(n_3091)
);

OR2x2_ASAP7_75t_L g3092 ( 
.A(n_2846),
.B(n_2545),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_2777),
.B(n_2711),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2784),
.B(n_2538),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2822),
.B(n_2538),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2814),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_3013),
.Y(n_3097)
);

OR2x2_ASAP7_75t_L g3098 ( 
.A(n_2813),
.B(n_2642),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2828),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2827),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_3025),
.A2(n_2699),
.B1(n_2697),
.B2(n_2722),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2830),
.Y(n_3102)
);

OR2x2_ASAP7_75t_L g3103 ( 
.A(n_2833),
.B(n_2589),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2873),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2877),
.Y(n_3105)
);

INVxp67_ASAP7_75t_SL g3106 ( 
.A(n_2996),
.Y(n_3106)
);

BUFx2_ASAP7_75t_L g3107 ( 
.A(n_3003),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2985),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2891),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2893),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2780),
.B(n_2559),
.Y(n_3111)
);

INVx2_ASAP7_75t_SL g3112 ( 
.A(n_2811),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2970),
.B(n_2559),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2880),
.B(n_2605),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2874),
.B(n_2753),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2896),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2793),
.Y(n_3117)
);

OAI221xp5_ASAP7_75t_L g3118 ( 
.A1(n_3025),
.A2(n_2601),
.B1(n_2663),
.B2(n_2606),
.C(n_2722),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_2773),
.B(n_2752),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_2776),
.B(n_2752),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2974),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2977),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2989),
.B(n_2941),
.Y(n_3123)
);

INVxp67_ASAP7_75t_SL g3124 ( 
.A(n_2996),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2964),
.B(n_2350),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2964),
.B(n_2350),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2898),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2900),
.Y(n_3128)
);

INVxp67_ASAP7_75t_SL g3129 ( 
.A(n_3020),
.Y(n_3129)
);

INVxp67_ASAP7_75t_SL g3130 ( 
.A(n_3020),
.Y(n_3130)
);

HB1xp67_ASAP7_75t_L g3131 ( 
.A(n_2794),
.Y(n_3131)
);

AND2x4_ASAP7_75t_SL g3132 ( 
.A(n_2801),
.B(n_2415),
.Y(n_3132)
);

BUFx2_ASAP7_75t_L g3133 ( 
.A(n_2998),
.Y(n_3133)
);

AND2x4_ASAP7_75t_L g3134 ( 
.A(n_2895),
.B(n_2675),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2924),
.B(n_2354),
.Y(n_3135)
);

AND2x4_ASAP7_75t_L g3136 ( 
.A(n_2801),
.B(n_2715),
.Y(n_3136)
);

NAND2x1p5_ASAP7_75t_L g3137 ( 
.A(n_2909),
.B(n_2715),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2872),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2930),
.B(n_2354),
.Y(n_3139)
);

INVx3_ASAP7_75t_L g3140 ( 
.A(n_2998),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2788),
.B(n_2565),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2832),
.A2(n_2581),
.B1(n_2508),
.B2(n_2662),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2791),
.B(n_2864),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2852),
.Y(n_3144)
);

AOI22xp33_ASAP7_75t_L g3145 ( 
.A1(n_2851),
.A2(n_2581),
.B1(n_2662),
.B2(n_2443),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2866),
.B(n_2565),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2870),
.B(n_2619),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_2772),
.A2(n_2443),
.B1(n_2449),
.B2(n_2681),
.Y(n_3148)
);

INVxp67_ASAP7_75t_SL g3149 ( 
.A(n_3023),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2772),
.A2(n_2449),
.B1(n_2681),
.B2(n_2657),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2825),
.B(n_2619),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_2794),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2976),
.B(n_2625),
.Y(n_3153)
);

BUFx3_ASAP7_75t_L g3154 ( 
.A(n_2821),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_2797),
.B(n_2526),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2979),
.B(n_2625),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2888),
.B(n_2630),
.Y(n_3157)
);

AND2x4_ASAP7_75t_SL g3158 ( 
.A(n_2785),
.B(n_2159),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2882),
.B(n_2747),
.Y(n_3159)
);

OR2x2_ASAP7_75t_L g3160 ( 
.A(n_2797),
.B(n_2803),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2853),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2991),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2882),
.B(n_2747),
.Y(n_3163)
);

INVxp67_ASAP7_75t_SL g3164 ( 
.A(n_3023),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2993),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2951),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2843),
.B(n_2630),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2953),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2816),
.B(n_2743),
.Y(n_3169)
);

NOR2x1_ASAP7_75t_R g3170 ( 
.A(n_2862),
.B(n_2724),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2921),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2956),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2958),
.Y(n_3173)
);

NOR2x1_ASAP7_75t_L g3174 ( 
.A(n_2933),
.B(n_2679),
.Y(n_3174)
);

NOR2x1_ASAP7_75t_L g3175 ( 
.A(n_2878),
.B(n_2679),
.Y(n_3175)
);

BUFx3_ASAP7_75t_L g3176 ( 
.A(n_2928),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_2848),
.A2(n_2657),
.B1(n_2527),
.B2(n_2531),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2966),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2944),
.B(n_2743),
.Y(n_3179)
);

OAI222xp33_ASAP7_75t_L g3180 ( 
.A1(n_2861),
.A2(n_2667),
.B1(n_2691),
.B2(n_2714),
.C1(n_2651),
.C2(n_2582),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2971),
.Y(n_3181)
);

INVxp33_ASAP7_75t_L g3182 ( 
.A(n_2886),
.Y(n_3182)
);

OAI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_3032),
.A2(n_2453),
.B(n_2756),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2803),
.B(n_2820),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_2834),
.B(n_2634),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_3024),
.B(n_3027),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2820),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2829),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_3031),
.B(n_2231),
.Y(n_3189)
);

INVx2_ASAP7_75t_SL g3190 ( 
.A(n_2980),
.Y(n_3190)
);

INVxp67_ASAP7_75t_SL g3191 ( 
.A(n_2764),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2914),
.B(n_2231),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2829),
.B(n_2527),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2858),
.B(n_2867),
.Y(n_3194)
);

INVxp67_ASAP7_75t_SL g3195 ( 
.A(n_2764),
.Y(n_3195)
);

AND2x4_ASAP7_75t_SL g3196 ( 
.A(n_2785),
.B(n_2185),
.Y(n_3196)
);

OR2x2_ASAP7_75t_SL g3197 ( 
.A(n_3005),
.B(n_2541),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_2858),
.B(n_2526),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2916),
.B(n_2244),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_2946),
.B(n_2244),
.Y(n_3200)
);

AND2x2_ASAP7_75t_L g3201 ( 
.A(n_2947),
.B(n_2274),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2949),
.B(n_2274),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2817),
.B(n_2281),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2867),
.B(n_2531),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2910),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2779),
.B(n_2641),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2911),
.Y(n_3207)
);

OR2x2_ASAP7_75t_L g3208 ( 
.A(n_2865),
.B(n_2641),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2950),
.B(n_2903),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2913),
.Y(n_3210)
);

INVx3_ASAP7_75t_L g3211 ( 
.A(n_2904),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2905),
.B(n_2303),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_2845),
.B(n_2988),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_3079),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3108),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3034),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_3096),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3160),
.B(n_2769),
.Y(n_3218)
);

OR2x2_ASAP7_75t_L g3219 ( 
.A(n_3184),
.B(n_2769),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3119),
.B(n_3011),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3037),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3120),
.B(n_2789),
.Y(n_3222)
);

OR2x2_ASAP7_75t_L g3223 ( 
.A(n_3184),
.B(n_2789),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3041),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3042),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3213),
.B(n_2800),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3099),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3141),
.B(n_2835),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_3048),
.B(n_2899),
.Y(n_3229)
);

OR2x2_ASAP7_75t_L g3230 ( 
.A(n_3194),
.B(n_2868),
.Y(n_3230)
);

BUFx2_ASAP7_75t_L g3231 ( 
.A(n_3087),
.Y(n_3231)
);

NAND2x1p5_ASAP7_75t_L g3232 ( 
.A(n_3074),
.B(n_2826),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3044),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3085),
.B(n_3012),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3052),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3053),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3075),
.B(n_3017),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_3107),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_3111),
.B(n_2954),
.Y(n_3239)
);

HB1xp67_ASAP7_75t_L g3240 ( 
.A(n_3106),
.Y(n_3240)
);

OR2x2_ASAP7_75t_L g3241 ( 
.A(n_3194),
.B(n_3051),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3185),
.B(n_3018),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3167),
.B(n_3028),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3054),
.Y(n_3244)
);

OR2x2_ASAP7_75t_L g3245 ( 
.A(n_3060),
.B(n_2883),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3192),
.B(n_2901),
.Y(n_3246)
);

HB1xp67_ASAP7_75t_L g3247 ( 
.A(n_3106),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3199),
.B(n_2901),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3143),
.B(n_2885),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3055),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_3123),
.B(n_2887),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3039),
.B(n_3093),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3088),
.B(n_3090),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3050),
.B(n_3009),
.Y(n_3254)
);

OR2x2_ASAP7_75t_L g3255 ( 
.A(n_3155),
.B(n_2906),
.Y(n_3255)
);

HB1xp67_ASAP7_75t_L g3256 ( 
.A(n_3124),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3035),
.B(n_3010),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3091),
.B(n_3097),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_3133),
.B(n_2967),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_3124),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3095),
.B(n_2855),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3064),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_3134),
.B(n_2954),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3146),
.B(n_2856),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3094),
.B(n_3021),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3065),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3179),
.B(n_2929),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3179),
.B(n_2929),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3083),
.B(n_2915),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3135),
.B(n_2781),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3206),
.B(n_2917),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_3198),
.B(n_2906),
.Y(n_3272)
);

INVx2_ASAP7_75t_SL g3273 ( 
.A(n_3074),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_3129),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3066),
.Y(n_3275)
);

OR2x2_ASAP7_75t_L g3276 ( 
.A(n_3057),
.B(n_2935),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3139),
.B(n_2781),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3067),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_3115),
.B(n_2799),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3208),
.B(n_2926),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3070),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3166),
.B(n_2932),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3072),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3071),
.B(n_3157),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3073),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3168),
.B(n_2934),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3078),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3153),
.B(n_3016),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_3156),
.B(n_3016),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3100),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3102),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3151),
.B(n_3019),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3063),
.B(n_3019),
.Y(n_3293)
);

OR2x2_ASAP7_75t_L g3294 ( 
.A(n_3057),
.B(n_2935),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3172),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_3089),
.B(n_2925),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3173),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3169),
.B(n_2799),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3169),
.B(n_2842),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3125),
.B(n_2842),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3178),
.B(n_2938),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_3126),
.B(n_2936),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3181),
.Y(n_3303)
);

OR2x2_ASAP7_75t_L g3304 ( 
.A(n_3086),
.B(n_2957),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3109),
.B(n_2940),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3215),
.Y(n_3306)
);

OAI22xp33_ASAP7_75t_SL g3307 ( 
.A1(n_3229),
.A2(n_3058),
.B1(n_3084),
.B2(n_3140),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3249),
.B(n_3086),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3216),
.Y(n_3309)
);

INVx1_ASAP7_75t_SL g3310 ( 
.A(n_3238),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3238),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3267),
.B(n_3110),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3221),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3224),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3225),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3267),
.B(n_3268),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_3251),
.B(n_3038),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3268),
.B(n_3116),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3233),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3235),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3265),
.B(n_3038),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3236),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3244),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3250),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3262),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3266),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3229),
.A2(n_3045),
.B(n_3061),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3228),
.B(n_3187),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3275),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3296),
.A2(n_3089),
.B1(n_3061),
.B2(n_3036),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3278),
.Y(n_3331)
);

INVxp67_ASAP7_75t_L g3332 ( 
.A(n_3231),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3257),
.B(n_3254),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3281),
.Y(n_3334)
);

AND2x4_ASAP7_75t_L g3335 ( 
.A(n_3263),
.B(n_3188),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3259),
.A2(n_3045),
.B(n_3180),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3283),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3285),
.Y(n_3338)
);

OAI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3296),
.A2(n_3076),
.B(n_2861),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3252),
.B(n_3043),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_SL g3341 ( 
.A(n_3232),
.B(n_3058),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3240),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3298),
.B(n_3142),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3287),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3284),
.B(n_3043),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3290),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3298),
.B(n_3142),
.Y(n_3347)
);

CKINVDCx16_ASAP7_75t_R g3348 ( 
.A(n_3263),
.Y(n_3348)
);

OR2x2_ASAP7_75t_L g3349 ( 
.A(n_3241),
.B(n_3047),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3269),
.B(n_2902),
.Y(n_3350)
);

HB1xp67_ASAP7_75t_L g3351 ( 
.A(n_3240),
.Y(n_3351)
);

NOR3xp33_ASAP7_75t_L g3352 ( 
.A(n_3259),
.B(n_3180),
.C(n_3118),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3291),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3237),
.B(n_3242),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3222),
.B(n_3186),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3295),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3237),
.B(n_3047),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3299),
.B(n_3117),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3299),
.B(n_3117),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3247),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3222),
.B(n_3131),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3297),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_3245),
.B(n_3131),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3247),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3256),
.Y(n_3365)
);

INVxp67_ASAP7_75t_SL g3366 ( 
.A(n_3256),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3242),
.B(n_3243),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_3260),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3303),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3219),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3255),
.B(n_3152),
.Y(n_3371)
);

OAI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3232),
.A2(n_3076),
.B(n_3183),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3260),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3264),
.B(n_3209),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_3263),
.B(n_3140),
.Y(n_3375)
);

BUFx3_ASAP7_75t_L g3376 ( 
.A(n_3273),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3223),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3274),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3274),
.Y(n_3379)
);

NOR3xp33_ASAP7_75t_L g3380 ( 
.A(n_3273),
.B(n_3118),
.C(n_3015),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3220),
.B(n_3152),
.Y(n_3381)
);

INVx1_ASAP7_75t_SL g3382 ( 
.A(n_3310),
.Y(n_3382)
);

OR2x2_ASAP7_75t_L g3383 ( 
.A(n_3358),
.B(n_3230),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3358),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3359),
.Y(n_3385)
);

AOI32xp33_ASAP7_75t_L g3386 ( 
.A1(n_3352),
.A2(n_3132),
.A3(n_3175),
.B1(n_3174),
.B2(n_3112),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3359),
.Y(n_3387)
);

AOI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3330),
.A2(n_3046),
.B1(n_3036),
.B2(n_3062),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3336),
.A2(n_3197),
.B1(n_3062),
.B2(n_3190),
.Y(n_3389)
);

OAI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3341),
.A2(n_2850),
.B1(n_3171),
.B2(n_3176),
.Y(n_3390)
);

NAND4xp25_ASAP7_75t_L g3391 ( 
.A(n_3327),
.B(n_3046),
.C(n_2770),
.D(n_2839),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3371),
.Y(n_3392)
);

OAI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3341),
.A2(n_2850),
.B1(n_3211),
.B2(n_3103),
.Y(n_3393)
);

HB1xp67_ASAP7_75t_L g3394 ( 
.A(n_3351),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3343),
.B(n_3220),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3348),
.B(n_3288),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_SL g3397 ( 
.A(n_3307),
.B(n_3170),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3354),
.B(n_3289),
.Y(n_3398)
);

OR2x2_ASAP7_75t_L g3399 ( 
.A(n_3316),
.B(n_3276),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3371),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3357),
.B(n_3234),
.Y(n_3401)
);

O2A1O1Ixp33_ASAP7_75t_SL g3402 ( 
.A1(n_3310),
.A2(n_3098),
.B(n_3080),
.C(n_2824),
.Y(n_3402)
);

AOI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_3339),
.A2(n_2823),
.B1(n_2836),
.B2(n_3101),
.Y(n_3403)
);

INVxp67_ASAP7_75t_L g3404 ( 
.A(n_3350),
.Y(n_3404)
);

OAI21xp33_ASAP7_75t_SL g3405 ( 
.A1(n_3366),
.A2(n_3195),
.B(n_3191),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3361),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3361),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3349),
.Y(n_3408)
);

OAI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3372),
.A2(n_3339),
.B(n_3332),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3375),
.B(n_3134),
.Y(n_3410)
);

OAI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3372),
.A2(n_2770),
.B1(n_3239),
.B2(n_3059),
.Y(n_3411)
);

OR2x2_ASAP7_75t_L g3412 ( 
.A(n_3316),
.B(n_3381),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3312),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3380),
.A2(n_3239),
.B1(n_3183),
.B2(n_3226),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3312),
.Y(n_3415)
);

INVx1_ASAP7_75t_SL g3416 ( 
.A(n_3376),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_3374),
.B(n_3182),
.Y(n_3417)
);

NAND3xp33_ASAP7_75t_L g3418 ( 
.A(n_3368),
.B(n_3177),
.C(n_3150),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3318),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3375),
.A2(n_2809),
.B(n_3059),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3343),
.B(n_3234),
.Y(n_3421)
);

NAND2x1p5_ASAP7_75t_L g3422 ( 
.A(n_3311),
.B(n_3049),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3318),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3363),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_3347),
.A2(n_3015),
.B(n_2775),
.C(n_3056),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3306),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3309),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3313),
.Y(n_3428)
);

NAND2x1_ASAP7_75t_L g3429 ( 
.A(n_3335),
.B(n_3239),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3347),
.B(n_3294),
.Y(n_3430)
);

AO22x1_ASAP7_75t_L g3431 ( 
.A1(n_3335),
.A2(n_3136),
.B1(n_2990),
.B2(n_2918),
.Y(n_3431)
);

BUFx2_ASAP7_75t_L g3432 ( 
.A(n_3345),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3342),
.A2(n_3130),
.B(n_3129),
.Y(n_3433)
);

HB1xp67_ASAP7_75t_L g3434 ( 
.A(n_3360),
.Y(n_3434)
);

INVxp67_ASAP7_75t_L g3435 ( 
.A(n_3314),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_SL g3436 ( 
.A1(n_3364),
.A2(n_3195),
.B(n_3191),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3315),
.Y(n_3437)
);

AOI211xp5_ASAP7_75t_L g3438 ( 
.A1(n_3370),
.A2(n_2714),
.B(n_2651),
.C(n_3069),
.Y(n_3438)
);

OR2x2_ASAP7_75t_L g3439 ( 
.A(n_3355),
.B(n_3304),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3365),
.Y(n_3440)
);

A2O1A1Ixp33_ASAP7_75t_SL g3441 ( 
.A1(n_3379),
.A2(n_3203),
.B(n_2844),
.C(n_2849),
.Y(n_3441)
);

OAI22xp33_ASAP7_75t_SL g3442 ( 
.A1(n_3319),
.A2(n_3154),
.B1(n_3137),
.B2(n_2850),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3320),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3322),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3323),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_3377),
.B(n_3272),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3373),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3324),
.Y(n_3448)
);

AOI211xp5_ASAP7_75t_L g3449 ( 
.A1(n_3389),
.A2(n_2907),
.B(n_2756),
.C(n_2881),
.Y(n_3449)
);

AOI31xp33_ASAP7_75t_L g3450 ( 
.A1(n_3402),
.A2(n_3137),
.A3(n_2857),
.B(n_3040),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_3405),
.B(n_3378),
.Y(n_3451)
);

AOI221xp5_ASAP7_75t_L g3452 ( 
.A1(n_3409),
.A2(n_3325),
.B1(n_3331),
.B2(n_3329),
.C(n_3326),
.Y(n_3452)
);

AOI322xp5_ASAP7_75t_L g3453 ( 
.A1(n_3414),
.A2(n_3340),
.A3(n_3308),
.B1(n_3367),
.B2(n_3321),
.C1(n_3317),
.C2(n_3333),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3429),
.B(n_3432),
.Y(n_3454)
);

INVxp67_ASAP7_75t_L g3455 ( 
.A(n_3397),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3392),
.Y(n_3456)
);

OAI221xp5_ASAP7_75t_L g3457 ( 
.A1(n_3411),
.A2(n_3328),
.B1(n_2875),
.B2(n_2889),
.C(n_2884),
.Y(n_3457)
);

OR2x2_ASAP7_75t_L g3458 ( 
.A(n_3430),
.B(n_3218),
.Y(n_3458)
);

AOI32xp33_ASAP7_75t_L g3459 ( 
.A1(n_3405),
.A2(n_3293),
.A3(n_3196),
.B1(n_3158),
.B2(n_3292),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3400),
.Y(n_3460)
);

OAI221xp5_ASAP7_75t_L g3461 ( 
.A1(n_3386),
.A2(n_2884),
.B1(n_2955),
.B2(n_3150),
.C(n_2963),
.Y(n_3461)
);

OAI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3425),
.A2(n_3436),
.B(n_3388),
.Y(n_3462)
);

OAI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_3388),
.A2(n_3211),
.B1(n_3130),
.B2(n_3164),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3391),
.A2(n_3418),
.B1(n_3424),
.B2(n_3408),
.Y(n_3464)
);

AOI21xp33_ASAP7_75t_L g3465 ( 
.A1(n_3441),
.A2(n_2955),
.B(n_2961),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3406),
.Y(n_3466)
);

O2A1O1Ixp33_ASAP7_75t_L g3467 ( 
.A1(n_3390),
.A2(n_3337),
.B(n_3338),
.C(n_3334),
.Y(n_3467)
);

AOI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3431),
.A2(n_3353),
.B1(n_3356),
.B2(n_3346),
.C(n_3344),
.Y(n_3468)
);

AOI211xp5_ASAP7_75t_L g3469 ( 
.A1(n_3442),
.A2(n_2881),
.B(n_2863),
.C(n_2986),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3407),
.Y(n_3470)
);

OAI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3382),
.A2(n_3148),
.B(n_3145),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_SL g3472 ( 
.A(n_3393),
.B(n_2908),
.Y(n_3472)
);

AOI221xp5_ASAP7_75t_L g3473 ( 
.A1(n_3435),
.A2(n_3369),
.B1(n_3362),
.B2(n_3271),
.C(n_3280),
.Y(n_3473)
);

XOR2x2_ASAP7_75t_SL g3474 ( 
.A(n_3422),
.B(n_3136),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3384),
.A2(n_3248),
.B1(n_3246),
.B2(n_3279),
.Y(n_3475)
);

OAI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3416),
.A2(n_3148),
.B(n_3145),
.Y(n_3476)
);

OAI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_3420),
.A2(n_3164),
.B1(n_3149),
.B2(n_2981),
.Y(n_3477)
);

AOI21xp33_ASAP7_75t_L g3478 ( 
.A1(n_3438),
.A2(n_3092),
.B(n_2968),
.Y(n_3478)
);

XOR2x2_ASAP7_75t_L g3479 ( 
.A(n_3417),
.B(n_2908),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3403),
.A2(n_3385),
.B1(n_3387),
.B2(n_3413),
.Y(n_3480)
);

AOI21xp33_ASAP7_75t_L g3481 ( 
.A1(n_3404),
.A2(n_2434),
.B(n_2831),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_SL g3482 ( 
.A1(n_3396),
.A2(n_3279),
.B1(n_3248),
.B2(n_3246),
.Y(n_3482)
);

NAND2xp33_ASAP7_75t_L g3483 ( 
.A(n_3410),
.B(n_2263),
.Y(n_3483)
);

AOI21xp33_ASAP7_75t_L g3484 ( 
.A1(n_3394),
.A2(n_2959),
.B(n_3253),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3415),
.B(n_2616),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3433),
.A2(n_2863),
.B(n_2962),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3426),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3421),
.B(n_3419),
.Y(n_3488)
);

OAI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_3403),
.A2(n_3177),
.B(n_2892),
.Y(n_3489)
);

NAND3xp33_ASAP7_75t_L g3490 ( 
.A(n_3427),
.B(n_2892),
.C(n_2778),
.Y(n_3490)
);

O2A1O1Ixp5_ASAP7_75t_L g3491 ( 
.A1(n_3428),
.A2(n_3258),
.B(n_3286),
.C(n_3282),
.Y(n_3491)
);

OAI311xp33_ASAP7_75t_L g3492 ( 
.A1(n_3462),
.A2(n_2774),
.A3(n_2815),
.B1(n_3395),
.C1(n_2871),
.Y(n_3492)
);

O2A1O1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3455),
.A2(n_3437),
.B(n_3444),
.C(n_3443),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3464),
.A2(n_3412),
.B1(n_3383),
.B2(n_3399),
.Y(n_3494)
);

O2A1O1Ixp33_ASAP7_75t_L g3495 ( 
.A1(n_3472),
.A2(n_3445),
.B(n_3448),
.C(n_3434),
.Y(n_3495)
);

OAI211xp5_ASAP7_75t_L g3496 ( 
.A1(n_3465),
.A2(n_3423),
.B(n_2778),
.C(n_2937),
.Y(n_3496)
);

AOI211xp5_ASAP7_75t_L g3497 ( 
.A1(n_3465),
.A2(n_3463),
.B(n_3461),
.C(n_3489),
.Y(n_3497)
);

OA22x2_ASAP7_75t_L g3498 ( 
.A1(n_3480),
.A2(n_3398),
.B1(n_3401),
.B2(n_3440),
.Y(n_3498)
);

AOI22x1_ASAP7_75t_L g3499 ( 
.A1(n_3474),
.A2(n_2263),
.B1(n_2826),
.B2(n_2225),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3479),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3487),
.Y(n_3501)
);

OAI221xp5_ASAP7_75t_L g3502 ( 
.A1(n_3459),
.A2(n_3468),
.B1(n_3467),
.B2(n_3453),
.C(n_3450),
.Y(n_3502)
);

AOI221xp5_ASAP7_75t_L g3503 ( 
.A1(n_3452),
.A2(n_3447),
.B1(n_3446),
.B2(n_3439),
.C(n_3305),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3483),
.A2(n_3301),
.B(n_3149),
.Y(n_3504)
);

OAI21xp5_ASAP7_75t_SL g3505 ( 
.A1(n_3477),
.A2(n_2808),
.B(n_2967),
.Y(n_3505)
);

AOI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3449),
.A2(n_3261),
.B1(n_3113),
.B2(n_3147),
.Y(n_3506)
);

OAI221xp5_ASAP7_75t_L g3507 ( 
.A1(n_3451),
.A2(n_3077),
.B1(n_2937),
.B2(n_3163),
.C(n_3159),
.Y(n_3507)
);

NAND3xp33_ASAP7_75t_L g3508 ( 
.A(n_3486),
.B(n_2314),
.C(n_2290),
.Y(n_3508)
);

AOI221xp5_ASAP7_75t_L g3509 ( 
.A1(n_3473),
.A2(n_3105),
.B1(n_3122),
.B2(n_3121),
.C(n_3104),
.Y(n_3509)
);

INVxp67_ASAP7_75t_L g3510 ( 
.A(n_3485),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3456),
.B(n_3243),
.Y(n_3511)
);

XOR2xp5_ASAP7_75t_L g3512 ( 
.A(n_3476),
.B(n_2194),
.Y(n_3512)
);

OAI221xp5_ASAP7_75t_L g3513 ( 
.A1(n_3457),
.A2(n_3077),
.B1(n_3163),
.B2(n_3159),
.C(n_2314),
.Y(n_3513)
);

OAI221xp5_ASAP7_75t_SL g3514 ( 
.A1(n_3469),
.A2(n_3302),
.B1(n_3300),
.B2(n_3277),
.C(n_3270),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3488),
.B(n_2718),
.Y(n_3515)
);

NAND3xp33_ASAP7_75t_SL g3516 ( 
.A(n_3454),
.B(n_2269),
.C(n_2952),
.Y(n_3516)
);

AOI211x1_ASAP7_75t_L g3517 ( 
.A1(n_3478),
.A2(n_3128),
.B(n_3144),
.C(n_3127),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3491),
.Y(n_3518)
);

NAND4xp75_ASAP7_75t_L g3519 ( 
.A(n_3471),
.B(n_2959),
.C(n_2366),
.D(n_2324),
.Y(n_3519)
);

NAND3xp33_ASAP7_75t_SL g3520 ( 
.A(n_3482),
.B(n_3490),
.C(n_3475),
.Y(n_3520)
);

OAI21xp33_ASAP7_75t_L g3521 ( 
.A1(n_3484),
.A2(n_3470),
.B(n_3466),
.Y(n_3521)
);

AO22x1_ASAP7_75t_L g3522 ( 
.A1(n_3460),
.A2(n_2920),
.B1(n_2922),
.B2(n_2904),
.Y(n_3522)
);

OAI221xp5_ASAP7_75t_L g3523 ( 
.A1(n_3481),
.A2(n_2324),
.B1(n_3204),
.B2(n_3193),
.C(n_3068),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3481),
.A2(n_3277),
.B1(n_3270),
.B2(n_3200),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3458),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3455),
.B(n_3161),
.Y(n_3526)
);

OAI21xp33_ASAP7_75t_L g3527 ( 
.A1(n_3462),
.A2(n_3068),
.B(n_3300),
.Y(n_3527)
);

OAI211xp5_ASAP7_75t_SL g3528 ( 
.A1(n_3462),
.A2(n_2860),
.B(n_2847),
.C(n_2890),
.Y(n_3528)
);

NAND3xp33_ASAP7_75t_L g3529 ( 
.A(n_3462),
.B(n_3201),
.C(n_3189),
.Y(n_3529)
);

OAI221xp5_ASAP7_75t_L g3530 ( 
.A1(n_3462),
.A2(n_3204),
.B1(n_3193),
.B2(n_3082),
.C(n_3114),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3487),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3464),
.B(n_3202),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3450),
.A2(n_2879),
.B(n_3081),
.Y(n_3533)
);

O2A1O1Ixp5_ASAP7_75t_L g3534 ( 
.A1(n_3462),
.A2(n_3138),
.B(n_3081),
.C(n_3162),
.Y(n_3534)
);

NAND3xp33_ASAP7_75t_L g3535 ( 
.A(n_3462),
.B(n_3212),
.C(n_2987),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_SL g3536 ( 
.A1(n_3450),
.A2(n_2397),
.B(n_2269),
.Y(n_3536)
);

NOR3xp33_ASAP7_75t_L g3537 ( 
.A(n_3462),
.B(n_2922),
.C(n_2920),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3474),
.B(n_3214),
.Y(n_3538)
);

O2A1O1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3492),
.A2(n_2664),
.B(n_2582),
.C(n_2654),
.Y(n_3539)
);

AOI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3520),
.A2(n_3302),
.B1(n_3165),
.B2(n_3207),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3518),
.B(n_3205),
.Y(n_3541)
);

NAND4xp25_ASAP7_75t_L g3542 ( 
.A(n_3497),
.B(n_2860),
.C(n_2847),
.D(n_2804),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3525),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3500),
.B(n_2194),
.Y(n_3544)
);

NAND4xp25_ASAP7_75t_L g3545 ( 
.A(n_3502),
.B(n_2810),
.C(n_2804),
.D(n_2890),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3503),
.B(n_3210),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3501),
.Y(n_3547)
);

NAND3xp33_ASAP7_75t_SL g3548 ( 
.A(n_3537),
.B(n_2952),
.C(n_2547),
.Y(n_3548)
);

NOR2x1_ASAP7_75t_L g3549 ( 
.A(n_3536),
.B(n_2923),
.Y(n_3549)
);

NOR3x1_ASAP7_75t_L g3550 ( 
.A(n_3516),
.B(n_3030),
.C(n_2810),
.Y(n_3550)
);

NOR3xp33_ASAP7_75t_L g3551 ( 
.A(n_3528),
.B(n_2649),
.C(n_2430),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3510),
.B(n_3214),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3531),
.Y(n_3553)
);

AOI221xp5_ASAP7_75t_L g3554 ( 
.A1(n_3530),
.A2(n_2986),
.B1(n_2945),
.B2(n_2995),
.C(n_2943),
.Y(n_3554)
);

NAND4xp25_ASAP7_75t_L g3555 ( 
.A(n_3527),
.B(n_2897),
.C(n_2894),
.D(n_3033),
.Y(n_3555)
);

OAI211xp5_ASAP7_75t_L g3556 ( 
.A1(n_3499),
.A2(n_2844),
.B(n_2849),
.C(n_2782),
.Y(n_3556)
);

NAND3xp33_ASAP7_75t_L g3557 ( 
.A(n_3535),
.B(n_2224),
.C(n_2419),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3517),
.B(n_3217),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_SL g3559 ( 
.A(n_3498),
.B(n_2994),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3512),
.B(n_2397),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3534),
.B(n_2994),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3495),
.A2(n_3538),
.B(n_3493),
.Y(n_3562)
);

NAND4xp25_ASAP7_75t_L g3563 ( 
.A(n_3529),
.B(n_2894),
.C(n_2897),
.D(n_2973),
.Y(n_3563)
);

NAND4xp25_ASAP7_75t_L g3564 ( 
.A(n_3508),
.B(n_2782),
.C(n_2997),
.D(n_2879),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3509),
.B(n_3494),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3511),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3515),
.B(n_2455),
.Y(n_3567)
);

NAND5xp2_ASAP7_75t_L g3568 ( 
.A(n_3505),
.B(n_2455),
.C(n_2723),
.D(n_2999),
.E(n_2992),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3526),
.Y(n_3569)
);

NOR3xp33_ASAP7_75t_L g3570 ( 
.A(n_3545),
.B(n_3565),
.C(n_3562),
.Y(n_3570)
);

NAND3xp33_ASAP7_75t_L g3571 ( 
.A(n_3540),
.B(n_3496),
.C(n_3514),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3552),
.Y(n_3572)
);

INVxp67_ASAP7_75t_SL g3573 ( 
.A(n_3544),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3541),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3543),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3547),
.Y(n_3576)
);

NOR3xp33_ASAP7_75t_L g3577 ( 
.A(n_3542),
.B(n_3523),
.C(n_3513),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3553),
.Y(n_3578)
);

OAI211xp5_ASAP7_75t_L g3579 ( 
.A1(n_3549),
.A2(n_3521),
.B(n_3533),
.C(n_3507),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3566),
.B(n_3569),
.Y(n_3580)
);

NOR2x1_ASAP7_75t_SL g3581 ( 
.A(n_3556),
.B(n_3519),
.Y(n_3581)
);

NOR3x1_ASAP7_75t_L g3582 ( 
.A(n_3559),
.B(n_3564),
.C(n_3548),
.Y(n_3582)
);

NOR3xp33_ASAP7_75t_L g3583 ( 
.A(n_3568),
.B(n_3522),
.C(n_3532),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3558),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3546),
.Y(n_3585)
);

NAND5xp2_ASAP7_75t_L g3586 ( 
.A(n_3560),
.B(n_3504),
.C(n_3492),
.D(n_3524),
.E(n_3506),
.Y(n_3586)
);

NOR3xp33_ASAP7_75t_L g3587 ( 
.A(n_3568),
.B(n_2187),
.C(n_2654),
.Y(n_3587)
);

NAND4xp25_ASAP7_75t_L g3588 ( 
.A(n_3550),
.B(n_2923),
.C(n_2960),
.D(n_3006),
.Y(n_3588)
);

INVxp67_ASAP7_75t_L g3589 ( 
.A(n_3567),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_L g3590 ( 
.A(n_3555),
.B(n_2960),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3561),
.B(n_3217),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_3563),
.B(n_3007),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3539),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3580),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3572),
.Y(n_3595)
);

NOR3x2_ASAP7_75t_L g3596 ( 
.A(n_3581),
.B(n_3582),
.C(n_3586),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3575),
.Y(n_3597)
);

NOR2x1_ASAP7_75t_L g3598 ( 
.A(n_3593),
.B(n_3557),
.Y(n_3598)
);

NOR2x1_ASAP7_75t_L g3599 ( 
.A(n_3586),
.B(n_2154),
.Y(n_3599)
);

NAND4xp75_ASAP7_75t_L g3600 ( 
.A(n_3584),
.B(n_3585),
.C(n_3578),
.D(n_3576),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3574),
.Y(n_3601)
);

NOR2x1_ASAP7_75t_L g3602 ( 
.A(n_3579),
.B(n_2154),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3570),
.B(n_3554),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3573),
.Y(n_3604)
);

NAND3xp33_ASAP7_75t_SL g3605 ( 
.A(n_3577),
.B(n_3551),
.C(n_2723),
.Y(n_3605)
);

NOR3x1_ASAP7_75t_L g3606 ( 
.A(n_3571),
.B(n_3026),
.C(n_2386),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3592),
.B(n_3590),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3589),
.B(n_3227),
.Y(n_3608)
);

NOR3xp33_ASAP7_75t_L g3609 ( 
.A(n_3588),
.B(n_2438),
.C(n_2437),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3591),
.Y(n_3610)
);

NOR2x1_ASAP7_75t_L g3611 ( 
.A(n_3583),
.B(n_2303),
.Y(n_3611)
);

OAI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_3587),
.A2(n_3022),
.B1(n_3114),
.B2(n_3082),
.Y(n_3612)
);

NAND3xp33_ASAP7_75t_L g3613 ( 
.A(n_3570),
.B(n_2224),
.C(n_2375),
.Y(n_3613)
);

INVxp67_ASAP7_75t_SL g3614 ( 
.A(n_3604),
.Y(n_3614)
);

XNOR2xp5_ASAP7_75t_L g3615 ( 
.A(n_3596),
.B(n_2931),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3594),
.B(n_3022),
.Y(n_3616)
);

NOR3xp33_ASAP7_75t_L g3617 ( 
.A(n_3605),
.B(n_2371),
.C(n_2333),
.Y(n_3617)
);

NAND2xp33_ASAP7_75t_L g3618 ( 
.A(n_3595),
.B(n_2588),
.Y(n_3618)
);

NOR2x1_ASAP7_75t_L g3619 ( 
.A(n_3600),
.B(n_3597),
.Y(n_3619)
);

XOR2x1_ASAP7_75t_L g3620 ( 
.A(n_3601),
.B(n_2156),
.Y(n_3620)
);

NAND4xp75_ASAP7_75t_L g3621 ( 
.A(n_3606),
.B(n_2156),
.C(n_2336),
.D(n_2375),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3608),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3610),
.B(n_2931),
.Y(n_3623)
);

NOR4xp75_ASAP7_75t_L g3624 ( 
.A(n_3603),
.B(n_2639),
.C(n_3007),
.D(n_2472),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3598),
.Y(n_3625)
);

AND2x4_ASAP7_75t_L g3626 ( 
.A(n_3607),
.B(n_2965),
.Y(n_3626)
);

NOR2x1_ASAP7_75t_L g3627 ( 
.A(n_3611),
.B(n_2691),
.Y(n_3627)
);

OR2x6_ASAP7_75t_L g3628 ( 
.A(n_3619),
.B(n_3625),
.Y(n_3628)
);

NOR2xp67_ASAP7_75t_L g3629 ( 
.A(n_3615),
.B(n_3612),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3614),
.B(n_3609),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3622),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3615),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3616),
.Y(n_3633)
);

AOI22xp5_ASAP7_75t_L g3634 ( 
.A1(n_3626),
.A2(n_3599),
.B1(n_3602),
.B2(n_3613),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3623),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_3627),
.B(n_2965),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3620),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3624),
.Y(n_3638)
);

XOR2x2_ASAP7_75t_L g3639 ( 
.A(n_3621),
.B(n_2419),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3628),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_3628),
.Y(n_3641)
);

AOI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3632),
.A2(n_3618),
.B1(n_3617),
.B2(n_2667),
.Y(n_3642)
);

INVx1_ASAP7_75t_SL g3643 ( 
.A(n_3631),
.Y(n_3643)
);

INVx2_ASAP7_75t_SL g3644 ( 
.A(n_3635),
.Y(n_3644)
);

OAI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3630),
.A2(n_2392),
.B(n_2380),
.Y(n_3645)
);

AO22x2_ASAP7_75t_L g3646 ( 
.A1(n_3633),
.A2(n_2972),
.B1(n_2975),
.B2(n_2969),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3638),
.B(n_3227),
.Y(n_3647)
);

XNOR2x1_ASAP7_75t_L g3648 ( 
.A(n_3640),
.B(n_3629),
.Y(n_3648)
);

OA22x2_ASAP7_75t_L g3649 ( 
.A1(n_3644),
.A2(n_3637),
.B1(n_3634),
.B2(n_3636),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3646),
.Y(n_3650)
);

XNOR2x1_ASAP7_75t_L g3651 ( 
.A(n_3649),
.B(n_3641),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3648),
.A2(n_3643),
.B1(n_3647),
.B2(n_3642),
.Y(n_3652)
);

AOI311xp33_ASAP7_75t_L g3653 ( 
.A1(n_3650),
.A2(n_3645),
.A3(n_3646),
.B(n_3639),
.C(n_2983),
.Y(n_3653)
);

INVxp67_ASAP7_75t_L g3654 ( 
.A(n_3651),
.Y(n_3654)
);

AO21x2_ASAP7_75t_L g3655 ( 
.A1(n_3654),
.A2(n_3652),
.B(n_3653),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3655),
.A2(n_2428),
.B(n_2211),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3656),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3657),
.A2(n_2457),
.B(n_2332),
.Y(n_3658)
);


endmodule