module real_aes_954_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g244 ( .A(n_0), .B(n_151), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_1), .B(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_2), .B(n_140), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_3), .B(n_149), .Y(n_475) );
INVx1_ASAP7_75t_L g139 ( .A(n_4), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_5), .B(n_140), .Y(n_197) );
NAND2xp33_ASAP7_75t_SL g190 ( .A(n_6), .B(n_146), .Y(n_190) );
INVx1_ASAP7_75t_L g170 ( .A(n_7), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_8), .Y(n_760) );
AND2x2_ASAP7_75t_L g195 ( .A(n_9), .B(n_130), .Y(n_195) );
AND2x2_ASAP7_75t_L g468 ( .A(n_10), .B(n_187), .Y(n_468) );
AND2x2_ASAP7_75t_L g477 ( .A(n_11), .B(n_162), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_12), .Y(n_763) );
INVx2_ASAP7_75t_L g131 ( .A(n_13), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_14), .B(n_149), .Y(n_530) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_15), .B(n_759), .C(n_761), .Y(n_758) );
AOI221x1_ASAP7_75t_L g184 ( .A1(n_16), .A2(n_134), .B1(n_185), .B2(n_187), .C(n_189), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_17), .B(n_140), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_18), .B(n_140), .Y(n_515) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_20), .A2(n_88), .B1(n_140), .B2(n_172), .Y(n_456) );
AOI221xp5_ASAP7_75t_SL g133 ( .A1(n_21), .A2(n_35), .B1(n_134), .B2(n_140), .C(n_147), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_22), .A2(n_134), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_23), .B(n_151), .Y(n_200) );
OR2x2_ASAP7_75t_L g132 ( .A(n_24), .B(n_87), .Y(n_132) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_24), .A2(n_87), .B(n_131), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_25), .B(n_149), .Y(n_161) );
INVxp67_ASAP7_75t_L g183 ( .A(n_26), .Y(n_183) );
AND2x2_ASAP7_75t_L g233 ( .A(n_27), .B(n_129), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_28), .A2(n_134), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_29), .A2(n_187), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_30), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_31), .A2(n_134), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_32), .B(n_149), .Y(n_510) );
AND2x2_ASAP7_75t_L g135 ( .A(n_33), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g146 ( .A(n_33), .B(n_139), .Y(n_146) );
INVx1_ASAP7_75t_L g179 ( .A(n_33), .Y(n_179) );
OR2x6_ASAP7_75t_L g115 ( .A(n_34), .B(n_116), .Y(n_115) );
INVxp67_ASAP7_75t_L g761 ( .A(n_34), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_36), .B(n_140), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_37), .A2(n_80), .B1(n_134), .B2(n_177), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_38), .B(n_149), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_39), .B(n_140), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_40), .B(n_151), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_41), .A2(n_134), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g247 ( .A(n_42), .B(n_129), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_43), .B(n_151), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_44), .B(n_129), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_45), .B(n_140), .Y(n_527) );
INVx1_ASAP7_75t_L g138 ( .A(n_46), .Y(n_138) );
INVx1_ASAP7_75t_L g143 ( .A(n_46), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_47), .B(n_149), .Y(n_466) );
AND2x2_ASAP7_75t_L g496 ( .A(n_48), .B(n_129), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_49), .B(n_140), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_50), .B(n_151), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_51), .B(n_151), .Y(n_509) );
AND2x2_ASAP7_75t_L g211 ( .A(n_52), .B(n_129), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_53), .B(n_140), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_54), .B(n_149), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_55), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_56), .B(n_140), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_57), .A2(n_134), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_58), .B(n_130), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_59), .B(n_151), .Y(n_208) );
AND2x2_ASAP7_75t_L g521 ( .A(n_60), .B(n_130), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_61), .A2(n_134), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_62), .B(n_149), .Y(n_201) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_63), .B(n_162), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_64), .B(n_151), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_65), .B(n_151), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_66), .A2(n_90), .B1(n_134), .B2(n_177), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_67), .A2(n_745), .B1(n_746), .B2(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_67), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_68), .B(n_149), .Y(n_518) );
OAI222xp33_ASAP7_75t_L g120 ( .A1(n_69), .A2(n_121), .B1(n_730), .B2(n_731), .C1(n_735), .C2(n_738), .Y(n_120) );
INVx1_ASAP7_75t_L g730 ( .A(n_69), .Y(n_730) );
INVx1_ASAP7_75t_L g136 ( .A(n_70), .Y(n_136) );
INVx1_ASAP7_75t_L g145 ( .A(n_70), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_71), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_72), .B(n_151), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_73), .A2(n_134), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_74), .A2(n_134), .B(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_75), .A2(n_134), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g512 ( .A(n_76), .B(n_130), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_77), .B(n_129), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_78), .B(n_140), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_79), .A2(n_82), .B1(n_140), .B2(n_172), .Y(n_216) );
INVx1_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_81), .B(n_117), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_83), .B(n_151), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_84), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g489 ( .A(n_85), .B(n_162), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_86), .A2(n_134), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_89), .B(n_149), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_91), .A2(n_134), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_92), .B(n_149), .Y(n_487) );
INVxp67_ASAP7_75t_L g186 ( .A(n_93), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_94), .B(n_140), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_95), .B(n_149), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_96), .A2(n_134), .B(n_159), .Y(n_158) );
BUFx2_ASAP7_75t_L g520 ( .A(n_97), .Y(n_520) );
BUFx2_ASAP7_75t_L g105 ( .A(n_98), .Y(n_105) );
BUFx2_ASAP7_75t_SL g742 ( .A(n_98), .Y(n_742) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_752), .B(n_762), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_120), .B(n_739), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_107), .A2(n_744), .B(n_749), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_119), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_R g751 ( .A(n_112), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_SL g443 ( .A(n_113), .B(n_115), .Y(n_443) );
OR2x6_ASAP7_75t_SL g729 ( .A(n_113), .B(n_114), .Y(n_729) );
OR2x2_ASAP7_75t_L g737 ( .A(n_113), .B(n_115), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_440), .B1(n_444), .B2(n_727), .Y(n_122) );
INVx2_ASAP7_75t_L g732 ( .A(n_123), .Y(n_732) );
INVx4_ASAP7_75t_L g747 ( .A(n_123), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_123), .Y(n_748) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_353), .Y(n_123) );
NAND3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_263), .C(n_303), .Y(n_124) );
O2A1O1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_165), .B(n_192), .C(n_219), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_126), .B(n_268), .Y(n_302) );
NOR2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_154), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g238 ( .A(n_128), .Y(n_238) );
INVx2_ASAP7_75t_L g254 ( .A(n_128), .Y(n_254) );
OR2x2_ASAP7_75t_L g266 ( .A(n_128), .B(n_155), .Y(n_266) );
AND2x2_ASAP7_75t_L g280 ( .A(n_128), .B(n_239), .Y(n_280) );
INVx1_ASAP7_75t_L g308 ( .A(n_128), .Y(n_308) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_128), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_128), .B(n_155), .Y(n_414) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_153), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_129), .Y(n_210) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_129), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_129), .A2(n_484), .B(n_485), .Y(n_483) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x4_ASAP7_75t_L g171 ( .A(n_131), .B(n_132), .Y(n_171) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
AND2x6_ASAP7_75t_L g151 ( .A(n_136), .B(n_142), .Y(n_151) );
INVx2_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
AND2x4_ASAP7_75t_L g177 ( .A(n_137), .B(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g149 ( .A(n_138), .B(n_144), .Y(n_149) );
INVx2_ASAP7_75t_L g174 ( .A(n_138), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_152), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_151), .B(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_152), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_152), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_152), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_152), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_152), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_152), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_152), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_152), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_152), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_152), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_152), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_152), .A2(n_530), .B(n_531), .Y(n_529) );
OR2x2_ASAP7_75t_L g235 ( .A(n_154), .B(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_154), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_154), .B(n_237), .Y(n_375) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g165 ( .A(n_155), .B(n_166), .Y(n_165) );
OR2x2_ASAP7_75t_L g234 ( .A(n_155), .B(n_167), .Y(n_234) );
OR2x2_ASAP7_75t_L g253 ( .A(n_155), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g282 ( .A(n_155), .Y(n_282) );
AND2x4_ASAP7_75t_SL g321 ( .A(n_155), .B(n_167), .Y(n_321) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_155), .Y(n_325) );
OR2x2_ASAP7_75t_L g342 ( .A(n_155), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g352 ( .A(n_155), .B(n_259), .Y(n_352) );
INVx1_ASAP7_75t_L g381 ( .A(n_155), .Y(n_381) );
OR2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_164), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_162), .Y(n_156) );
INVx2_ASAP7_75t_SL g214 ( .A(n_162), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_162), .A2(n_515), .B(n_516), .Y(n_514) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_165), .B(n_310), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_166), .B(n_239), .Y(n_256) );
AND2x2_ASAP7_75t_L g268 ( .A(n_166), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g286 ( .A(n_166), .B(n_253), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_166), .B(n_307), .Y(n_306) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g259 ( .A(n_167), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g281 ( .A(n_167), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g316 ( .A(n_167), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_167), .B(n_239), .Y(n_340) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B1(n_177), .B2(n_182), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_171), .B(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_171), .B(n_186), .Y(n_185) );
NOR3xp33_ASAP7_75t_L g189 ( .A(n_171), .B(n_190), .C(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_171), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_171), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_171), .A2(n_527), .B(n_528), .Y(n_526) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_176), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2x1p5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g505 ( .A(n_187), .Y(n_505) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_188), .A2(n_241), .B(n_247), .Y(n_240) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_188), .A2(n_462), .B(n_468), .Y(n_461) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_193), .B(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g289 ( .A(n_193), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_193), .B(n_203), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_193), .B(n_310), .C(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g357 ( .A(n_193), .B(n_262), .Y(n_357) );
INVx5_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g224 ( .A(n_194), .B(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_SL g261 ( .A(n_194), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
OR2x2_ASAP7_75t_L g300 ( .A(n_194), .B(n_290), .Y(n_300) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_194), .Y(n_317) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_194), .B(n_223), .Y(n_335) );
AND2x4_ASAP7_75t_L g350 ( .A(n_194), .B(n_226), .Y(n_350) );
AND2x2_ASAP7_75t_L g364 ( .A(n_194), .B(n_203), .Y(n_364) );
OR2x2_ASAP7_75t_L g385 ( .A(n_194), .B(n_212), .Y(n_385) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
AND2x2_ASAP7_75t_L g439 ( .A(n_202), .B(n_317), .Y(n_439) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_212), .Y(n_202) );
AND2x4_ASAP7_75t_L g262 ( .A(n_203), .B(n_225), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_203), .B(n_223), .Y(n_278) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_203), .Y(n_311) );
OR2x2_ASAP7_75t_L g334 ( .A(n_203), .B(n_226), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_203), .B(n_226), .Y(n_337) );
INVx1_ASAP7_75t_L g346 ( .A(n_203), .Y(n_346) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_210), .A2(n_227), .B(n_233), .Y(n_226) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_210), .A2(n_227), .B(n_233), .Y(n_290) );
AOI21x1_ASAP7_75t_L g470 ( .A1(n_210), .A2(n_471), .B(n_477), .Y(n_470) );
AND2x2_ASAP7_75t_L g249 ( .A(n_212), .B(n_226), .Y(n_249) );
BUFx2_ASAP7_75t_L g298 ( .A(n_212), .Y(n_298) );
AND2x2_ASAP7_75t_L g393 ( .A(n_212), .B(n_273), .Y(n_393) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
AOI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_218), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
OAI221xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_234), .B1(n_235), .B2(n_248), .C(n_250), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
NOR2x1_ASAP7_75t_L g295 ( .A(n_222), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_222), .B(n_289), .Y(n_329) );
OR2x2_ASAP7_75t_L g341 ( .A(n_222), .B(n_337), .Y(n_341) );
OR2x2_ASAP7_75t_L g344 ( .A(n_222), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g433 ( .A(n_222), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g272 ( .A(n_223), .B(n_273), .Y(n_272) );
OA33x2_ASAP7_75t_L g305 ( .A1(n_223), .A2(n_266), .A3(n_306), .B1(n_309), .B2(n_312), .B3(n_315), .Y(n_305) );
OR2x2_ASAP7_75t_L g336 ( .A(n_223), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g360 ( .A(n_223), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g368 ( .A(n_223), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g388 ( .A(n_223), .B(n_262), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_223), .B(n_277), .Y(n_426) );
INVx2_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
AOI322xp5_ASAP7_75t_L g366 ( .A1(n_224), .A2(n_279), .A3(n_367), .B1(n_370), .B2(n_371), .C1(n_373), .C2(n_375), .Y(n_366) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_226), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_232), .Y(n_227) );
OR2x2_ASAP7_75t_L g348 ( .A(n_234), .B(n_327), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_234), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g421 ( .A(n_234), .Y(n_421) );
INVx1_ASAP7_75t_SL g287 ( .A(n_235), .Y(n_287) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g320 ( .A(n_237), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
INVx1_ASAP7_75t_L g269 ( .A(n_239), .Y(n_269) );
INVx1_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
OR2x2_ASAP7_75t_L g327 ( .A(n_239), .B(n_254), .Y(n_327) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_239), .Y(n_402) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_246), .Y(n_241) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_249), .B(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_257), .B(n_261), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_251), .A2(n_325), .B(n_326), .C(n_328), .Y(n_324) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g389 ( .A(n_253), .B(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_254), .Y(n_258) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g413 ( .A(n_256), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_259), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g390 ( .A(n_259), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_259), .B(n_381), .Y(n_398) );
INVx3_ASAP7_75t_SL g323 ( .A(n_262), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_270), .B1(n_274), .B2(n_279), .C(n_283), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_269), .Y(n_314) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_272), .A2(n_299), .B(n_371), .Y(n_377) );
AND2x2_ASAP7_75t_L g403 ( .A(n_272), .B(n_350), .Y(n_403) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_277), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g412 ( .A(n_277), .B(n_334), .Y(n_412) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g361 ( .A(n_280), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B(n_292), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx2_ASAP7_75t_L g434 ( .A(n_289), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_290), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g363 ( .A(n_290), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_291), .B(n_313), .Y(n_312) );
OAI31xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .A3(n_297), .B(n_301), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_296), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g374 ( .A(n_298), .B(n_300), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_298), .B(n_350), .Y(n_429) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR5xp2_ASAP7_75t_L g303 ( .A(n_304), .B(n_318), .C(n_330), .D(n_339), .E(n_347), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_308), .B(n_310), .Y(n_343) );
INVx1_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_308), .Y(n_420) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVxp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI321xp33_ASAP7_75t_L g355 ( .A1(n_316), .A2(n_356), .A3(n_358), .B1(n_362), .B2(n_365), .C(n_366), .Y(n_355) );
INVx1_ASAP7_75t_L g409 ( .A(n_317), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_324), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_320), .A2(n_393), .B1(n_400), .B2(n_403), .Y(n_399) );
AND2x2_ASAP7_75t_L g428 ( .A(n_321), .B(n_402), .Y(n_428) );
INVx1_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_337), .A2(n_348), .B1(n_349), .B2(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_342), .B2(n_344), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_346), .B(n_350), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_348), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_430), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_348), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_349), .A2(n_406), .B1(n_413), .B2(n_415), .C(n_416), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_351), .A2(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_404), .Y(n_353) );
NOR3xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_376), .C(n_394), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_357), .Y(n_423) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g422 ( .A(n_365), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_367), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g415 ( .A(n_375), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_384), .B(n_386), .Y(n_378) );
INVxp67_ASAP7_75t_L g436 ( .A(n_379), .Y(n_436) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_SL g391 ( .A(n_382), .Y(n_391) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_391), .B2(n_392), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_399), .Y(n_394) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_424), .C(n_435), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_422), .B(n_423), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_428), .A2(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx4_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
CKINVDCx6p67_ASAP7_75t_R g733 ( .A(n_441), .Y(n_733) );
INVx3_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g734 ( .A(n_444), .Y(n_734) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_664), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_580), .C(n_617), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_548), .C(n_563), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_493), .B1(n_522), .B2(n_534), .C(n_535), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_450), .B(n_478), .Y(n_449) );
OAI22xp33_ASAP7_75t_SL g608 ( .A1(n_450), .A2(n_572), .B1(n_609), .B2(n_612), .Y(n_608) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .Y(n_450) );
OAI21xp33_ASAP7_75t_SL g618 ( .A1(n_451), .A2(n_619), .B(n_625), .Y(n_618) );
OR2x2_ASAP7_75t_L g647 ( .A(n_451), .B(n_480), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_451), .B(n_567), .Y(n_648) );
INVx2_ASAP7_75t_L g679 ( .A(n_451), .Y(n_679) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_452), .B(n_539), .Y(n_660) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_461), .Y(n_534) );
BUFx3_ASAP7_75t_L g560 ( .A(n_453), .Y(n_560) );
AND2x2_ASAP7_75t_L g696 ( .A(n_453), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g719 ( .A(n_453), .B(n_481), .Y(n_719) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x4_ASAP7_75t_L g492 ( .A(n_454), .B(n_455), .Y(n_492) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_459), .B(n_481), .Y(n_639) );
INVx1_ASAP7_75t_L g676 ( .A(n_459), .Y(n_676) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_469), .Y(n_459) );
AND2x2_ASAP7_75t_L g491 ( .A(n_460), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g697 ( .A(n_460), .Y(n_697) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g540 ( .A(n_461), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_461), .B(n_469), .Y(n_541) );
AND2x2_ASAP7_75t_L g562 ( .A(n_461), .B(n_482), .Y(n_562) );
AND2x2_ASAP7_75t_L g644 ( .A(n_461), .B(n_470), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
AND2x4_ASAP7_75t_SL g537 ( .A(n_469), .B(n_482), .Y(n_537) );
INVx1_ASAP7_75t_L g568 ( .A(n_469), .Y(n_568) );
INVx2_ASAP7_75t_L g576 ( .A(n_469), .Y(n_576) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_469), .Y(n_600) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_470), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
AND2x2_ASAP7_75t_L g715 ( .A(n_479), .B(n_578), .Y(n_715) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_481), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g626 ( .A(n_481), .B(n_541), .Y(n_626) );
AND2x2_ASAP7_75t_L g643 ( .A(n_481), .B(n_644), .Y(n_643) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g567 ( .A(n_482), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g583 ( .A(n_482), .Y(n_583) );
AND2x2_ASAP7_75t_L g627 ( .A(n_482), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g634 ( .A(n_482), .B(n_635), .Y(n_634) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_482), .B(n_540), .Y(n_649) );
BUFx2_ASAP7_75t_L g659 ( .A(n_482), .Y(n_659) );
AND2x2_ASAP7_75t_L g684 ( .A(n_482), .B(n_644), .Y(n_684) );
AND2x2_ASAP7_75t_L g705 ( .A(n_482), .B(n_706), .Y(n_705) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .Y(n_482) );
INVx1_ASAP7_75t_L g636 ( .A(n_490), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_491), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g666 ( .A(n_491), .B(n_537), .Y(n_666) );
INVx3_ASAP7_75t_L g573 ( .A(n_492), .Y(n_573) );
AND2x2_ASAP7_75t_L g706 ( .A(n_492), .B(n_628), .Y(n_706) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_494), .A2(n_536), .B1(n_541), .B2(n_542), .Y(n_535) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx4_ASAP7_75t_L g533 ( .A(n_495), .Y(n_533) );
INVx2_ASAP7_75t_L g570 ( .A(n_495), .Y(n_570) );
NAND2x1_ASAP7_75t_L g596 ( .A(n_495), .B(n_513), .Y(n_596) );
OR2x2_ASAP7_75t_L g611 ( .A(n_495), .B(n_546), .Y(n_611) );
OR2x2_ASAP7_75t_SL g638 ( .A(n_495), .B(n_610), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_495), .B(n_525), .Y(n_651) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_495), .Y(n_672) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g551 ( .A(n_503), .Y(n_551) );
AND2x2_ASAP7_75t_L g683 ( .A(n_503), .B(n_657), .Y(n_683) );
NOR2x1_ASAP7_75t_SL g503 ( .A(n_504), .B(n_513), .Y(n_503) );
AND2x2_ASAP7_75t_L g524 ( .A(n_504), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g700 ( .A(n_504), .B(n_623), .Y(n_700) );
AO21x1_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_504) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
OR2x2_ASAP7_75t_L g532 ( .A(n_513), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g543 ( .A(n_513), .B(n_533), .Y(n_543) );
AND2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_546), .Y(n_589) );
OR2x2_ASAP7_75t_L g610 ( .A(n_513), .B(n_525), .Y(n_610) );
INVx2_ASAP7_75t_SL g616 ( .A(n_513), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_513), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g632 ( .A(n_513), .B(n_615), .Y(n_632) );
BUFx2_ASAP7_75t_L g654 ( .A(n_513), .Y(n_654) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_521), .Y(n_513) );
INVx2_ASAP7_75t_L g701 ( .A(n_522), .Y(n_701) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
OR2x2_ASAP7_75t_L g726 ( .A(n_523), .B(n_570), .Y(n_726) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_524), .B(n_533), .Y(n_592) );
AND2x2_ASAP7_75t_L g663 ( .A(n_524), .B(n_543), .Y(n_663) );
INVx1_ASAP7_75t_L g545 ( .A(n_525), .Y(n_545) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_525), .Y(n_554) );
INVx1_ASAP7_75t_L g587 ( .A(n_525), .Y(n_587) );
INVx2_ASAP7_75t_L g623 ( .A(n_525), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g553 ( .A(n_533), .B(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g613 ( .A(n_533), .Y(n_613) );
INVx2_ASAP7_75t_SL g689 ( .A(n_534), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_536), .A2(n_591), .B1(n_593), .B2(n_597), .Y(n_590) );
AND2x2_ASAP7_75t_SL g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g717 ( .A(n_537), .B(n_573), .Y(n_717) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_539), .B(n_583), .Y(n_662) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g628 ( .A(n_540), .B(n_576), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_541), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g571 ( .A(n_542), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_542), .A2(n_686), .B1(n_690), .B2(n_692), .C(n_694), .Y(n_685) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g555 ( .A(n_543), .B(n_556), .Y(n_555) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_543), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_543), .B(n_586), .Y(n_641) );
INVx1_ASAP7_75t_SL g637 ( .A(n_544), .Y(n_637) );
AOI221xp5_ASAP7_75t_SL g665 ( .A1(n_544), .A2(n_555), .B1(n_666), .B2(n_667), .C(n_670), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_544), .A2(n_616), .A3(n_643), .B1(n_699), .B2(n_701), .C1(n_702), .C2(n_705), .Y(n_698) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
BUFx2_ASAP7_75t_L g565 ( .A(n_545), .Y(n_565) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_546), .Y(n_557) );
INVx2_ASAP7_75t_L g615 ( .A(n_546), .Y(n_615) );
AND2x2_ASAP7_75t_L g656 ( .A(n_546), .B(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OA21x2_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_555), .B(n_558), .Y(n_548) );
AOI211xp5_ASAP7_75t_L g718 ( .A1(n_549), .A2(n_719), .B(n_720), .C(n_724), .Y(n_718) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OR2x2_ASAP7_75t_L g607 ( .A(n_551), .B(n_569), .Y(n_607) );
OR2x2_ASAP7_75t_L g691 ( .A(n_551), .B(n_586), .Y(n_691) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g631 ( .A(n_553), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g709 ( .A(n_556), .Y(n_709) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g595 ( .A(n_557), .Y(n_595) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
OR2x2_ASAP7_75t_L g564 ( .A(n_560), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g599 ( .A(n_562), .B(n_600), .Y(n_599) );
OAI322xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .A3(n_569), .B1(n_571), .B2(n_572), .C1(n_577), .C2(n_579), .Y(n_563) );
INVx1_ASAP7_75t_L g605 ( .A(n_564), .Y(n_605) );
OR2x2_ASAP7_75t_L g577 ( .A(n_566), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_566), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g588 ( .A(n_570), .B(n_589), .Y(n_588) );
OAI32xp33_ASAP7_75t_L g633 ( .A1(n_570), .A2(n_634), .A3(n_637), .B1(n_638), .B2(n_639), .Y(n_633) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g578 ( .A(n_573), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_573), .B(n_636), .Y(n_635) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_573), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g699 ( .A(n_573), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g620 ( .A(n_574), .Y(n_620) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_578), .B(n_644), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_601), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_590), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_SL g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g650 ( .A(n_589), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_592), .A2(n_612), .B1(n_714), .B2(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_594), .A2(n_641), .B(n_642), .C(n_645), .Y(n_640) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx3_ASAP7_75t_L g722 ( .A(n_596), .Y(n_722) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g603 ( .A(n_600), .Y(n_603) );
AO21x1_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B(n_608), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g668 ( .A(n_603), .Y(n_668) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_609), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g624 ( .A(n_611), .Y(n_624) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g681 ( .A(n_614), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_640), .C(n_652), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_621), .A2(n_683), .B(n_684), .Y(n_682) );
AND2x4_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
O2A1O1Ixp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_627), .B(n_629), .C(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_635), .Y(n_725) );
INVx2_ASAP7_75t_L g710 ( .A(n_638), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g724 ( .A1(n_639), .A2(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g704 ( .A(n_644), .Y(n_704) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .A3(n_649), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g723 ( .A(n_651), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_658), .B(n_661), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
BUFx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g673 ( .A(n_656), .Y(n_673) );
AOI21xp33_ASAP7_75t_SL g720 ( .A1(n_658), .A2(n_721), .B(n_723), .Y(n_720) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g688 ( .A(n_659), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_659), .B(n_679), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_659), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g669 ( .A(n_660), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_665), .B(n_685), .C(n_698), .D(n_707), .E(n_718), .Y(n_664) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_677), .B2(n_680), .C(n_682), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_713), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OA22x2_ASAP7_75t_L g731 ( .A1(n_727), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
CKINVDCx11_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g764 ( .A(n_755), .Y(n_764) );
INVx3_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
endmodule