module real_aes_3392_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
HB1xp67_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
AND2x4_ASAP7_75t_L g29 ( .A(n_0), .B(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_1), .B(n_4), .Y(n_18) );
INVx1_ASAP7_75t_L g23 ( .A(n_2), .Y(n_23) );
INVx2_ASAP7_75t_SL g27 ( .A(n_3), .Y(n_27) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
BUFx3_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
O2A1O1Ixp33_ASAP7_75t_SL g6 ( .A1(n_7), .A2(n_19), .B(n_24), .C(n_28), .Y(n_6) );
AOI21xp33_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_11), .B(n_16), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
BUFx3_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVxp33_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_13), .B(n_14), .Y(n_12) );
INVxp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
NAND2xp33_ASAP7_75t_L g19 ( .A(n_20), .B(n_21), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
endmodule