module fake_jpeg_26851_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_5),
.B1(n_10),
.B2(n_7),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_13),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_1),
.C(n_2),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_25),
.B2(n_4),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_29),
.B(n_28),
.Y(n_32)
);

OAI221xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_3),
.B1(n_23),
.B2(n_12),
.C(n_6),
.Y(n_33)
);


endmodule