module fake_jpeg_16114_n_386 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_5),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_41),
.B(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_45),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_5),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_57),
.Y(n_81)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_21),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_13),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_66),
.B(n_67),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_31),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_35),
.B1(n_18),
.B2(n_15),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_84),
.B1(n_98),
.B2(n_100),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_2),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_35),
.B1(n_15),
.B2(n_18),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_82),
.A2(n_86),
.B1(n_102),
.B2(n_90),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_35),
.B1(n_18),
.B2(n_15),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_87),
.B(n_101),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_39),
.A2(n_31),
.B1(n_32),
.B2(n_16),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_96),
.B1(n_104),
.B2(n_112),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_115),
.B1(n_14),
.B2(n_6),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_94),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_37),
.B1(n_22),
.B2(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_103),
.B(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_42),
.A2(n_22),
.B1(n_17),
.B2(n_28),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_55),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_21),
.C(n_33),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_83),
.Y(n_135)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_50),
.A2(n_37),
.B1(n_28),
.B2(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_116),
.B1(n_81),
.B2(n_91),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_38),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_54),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_33),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_3),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_47),
.A2(n_24),
.B1(n_19),
.B2(n_23),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_19),
.B1(n_23),
.B2(n_33),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_19),
.B1(n_57),
.B2(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_121),
.A2(n_145),
.B1(n_146),
.B2(n_89),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_135),
.Y(n_191)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_127),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_14),
.B(n_5),
.C(n_8),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_94),
.B(n_152),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_4),
.B1(n_12),
.B2(n_11),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_129),
.A2(n_139),
.B1(n_148),
.B2(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_130),
.A2(n_74),
.B1(n_80),
.B2(n_94),
.Y(n_192)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_140),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_4),
.B1(n_11),
.B2(n_8),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_4),
.B1(n_11),
.B2(n_8),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_3),
.B1(n_13),
.B2(n_2),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_90),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_156),
.B1(n_142),
.B2(n_166),
.Y(n_200)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_71),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_1),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_67),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_162),
.Y(n_171)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_73),
.B(n_1),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_2),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_74),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_85),
.A2(n_75),
.B1(n_77),
.B2(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_106),
.B(n_79),
.C(n_89),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_85),
.A2(n_75),
.B1(n_77),
.B2(n_99),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_81),
.B1(n_99),
.B2(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_169),
.B(n_190),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_176),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_174),
.B1(n_213),
.B2(n_204),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_101),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_173),
.A2(n_126),
.B(n_138),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_113),
.C(n_80),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_187),
.C(n_169),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_181),
.B(n_202),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_124),
.A2(n_87),
.B1(n_79),
.B2(n_89),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_184),
.A2(n_192),
.B1(n_194),
.B2(n_196),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_117),
.C(n_162),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g194 ( 
.A1(n_120),
.A2(n_94),
.B1(n_132),
.B2(n_134),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_186),
.B(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_137),
.A2(n_122),
.B1(n_132),
.B2(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_202),
.B1(n_207),
.B2(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_150),
.B1(n_127),
.B2(n_159),
.Y(n_202)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_128),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_143),
.A2(n_154),
.B1(n_155),
.B2(n_131),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_145),
.B(n_158),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_156),
.A2(n_131),
.B1(n_123),
.B2(n_140),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_141),
.A2(n_160),
.B1(n_151),
.B2(n_144),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_149),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_SL g260 ( 
.A(n_216),
.B(n_225),
.C(n_227),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_220),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_118),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_222),
.B(n_224),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_223),
.A2(n_239),
.B(n_240),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_119),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_228),
.Y(n_288)
);

BUFx12f_ASAP7_75t_SL g227 ( 
.A(n_204),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_231),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_227),
.B1(n_249),
.B2(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_236),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_241),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_178),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_250),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_180),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_171),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_173),
.C(n_187),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_246),
.Y(n_275)
);

BUFx24_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_191),
.C(n_181),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_188),
.B(n_191),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_200),
.C(n_194),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_254),
.A2(n_256),
.B1(n_250),
.B2(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_194),
.A2(n_183),
.B1(n_172),
.B2(n_195),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_172),
.B1(n_190),
.B2(n_211),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_258),
.A2(n_261),
.B1(n_262),
.B2(n_278),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_172),
.B1(n_184),
.B2(n_215),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_201),
.B1(n_252),
.B2(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_285),
.B1(n_290),
.B2(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_235),
.B1(n_233),
.B2(n_237),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_216),
.B(n_236),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_225),
.A2(n_235),
.B(n_232),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_271),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_237),
.A2(n_234),
.B1(n_240),
.B2(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_218),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_220),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_225),
.B1(n_242),
.B2(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_294),
.B(n_310),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_298),
.B1(n_303),
.B2(n_305),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_223),
.B(n_225),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_301),
.B(n_317),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_241),
.B1(n_239),
.B2(n_222),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_272),
.A2(n_226),
.B(n_247),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_274),
.B1(n_286),
.B2(n_280),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_247),
.B(n_231),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_231),
.B1(n_247),
.B2(n_260),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_302),
.A2(n_311),
.B1(n_312),
.B2(n_268),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_258),
.B1(n_283),
.B2(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_275),
.C(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_277),
.C(n_267),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_285),
.B1(n_261),
.B2(n_260),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_284),
.B1(n_259),
.B2(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_308),
.B1(n_316),
.B2(n_317),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_264),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_277),
.A3(n_270),
.B1(n_288),
.B2(n_267),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_313),
.B(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_257),
.B(n_263),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_327),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_299),
.B(n_315),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_263),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_325),
.C(n_331),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_268),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_326),
.A2(n_330),
.B1(n_329),
.B2(n_331),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_303),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_334),
.Y(n_345)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_302),
.A2(n_301),
.B1(n_305),
.B2(n_300),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_318),
.C(n_314),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_307),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_318),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_339),
.Y(n_352)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_312),
.B(n_297),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g351 ( 
.A1(n_338),
.A2(n_326),
.B(n_330),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_291),
.C(n_299),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_333),
.B(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_356),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_297),
.B1(n_309),
.B2(n_292),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_354),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_320),
.B(n_324),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_348),
.B(n_355),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_353),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_356),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_R g357 ( 
.A1(n_351),
.A2(n_328),
.B1(n_322),
.B2(n_319),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_335),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_327),
.B1(n_336),
.B2(n_325),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_363),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_340),
.C(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_364),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_343),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_346),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_345),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_354),
.C(n_345),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_366),
.A2(n_348),
.B(n_347),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_372),
.B(n_362),
.Y(n_378)
);

OAI321xp33_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_342),
.A3(n_341),
.B1(n_344),
.B2(n_347),
.C(n_350),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_367),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_374),
.B(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_375),
.Y(n_379)
);

AOI31xp33_ASAP7_75t_SL g380 ( 
.A1(n_376),
.A2(n_377),
.A3(n_378),
.B(n_361),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_361),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_380),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_379),
.Y(n_382)
);

OAI311xp33_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_365),
.A3(n_373),
.B1(n_377),
.C1(n_360),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_366),
.B1(n_358),
.B2(n_371),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_363),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_364),
.Y(n_386)
);


endmodule