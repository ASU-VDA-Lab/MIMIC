module real_aes_18203_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g836 ( .A(n_0), .Y(n_836) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_2), .A2(n_161), .B1(n_386), .B2(n_395), .Y(n_573) );
OAI22xp33_ASAP7_75t_SL g589 ( .A1(n_2), .A2(n_161), .B1(n_405), .B2(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g690 ( .A(n_3), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_3), .A2(n_575), .B(n_695), .C(n_696), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_4), .A2(n_369), .B(n_526), .C(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g960 ( .A(n_4), .Y(n_960) );
INVx1_ASAP7_75t_L g887 ( .A(n_5), .Y(n_887) );
INVx1_ASAP7_75t_L g1264 ( .A(n_6), .Y(n_1264) );
INVx1_ASAP7_75t_L g818 ( .A(n_7), .Y(n_818) );
INVx1_ASAP7_75t_L g259 ( .A(n_8), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_8), .B(n_269), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_9), .A2(n_215), .B1(n_499), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_9), .A2(n_49), .B1(n_465), .B2(n_479), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g1239 ( .A1(n_10), .A2(n_368), .B(n_575), .C(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1248 ( .A(n_10), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1321 ( .A1(n_11), .A2(n_194), .B1(n_261), .B2(n_850), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_11), .A2(n_194), .B1(n_989), .B2(n_1245), .Y(n_1329) );
INVx1_ASAP7_75t_L g631 ( .A(n_12), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g753 ( .A1(n_13), .A2(n_196), .B1(n_380), .B2(n_387), .C1(n_754), .C2(n_755), .Y(n_753) );
OAI222xp33_ASAP7_75t_L g786 ( .A1(n_13), .A2(n_134), .B1(n_196), .B2(n_787), .C1(n_788), .C2(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g965 ( .A(n_14), .Y(n_965) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_15), .B(n_1051), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_15), .B(n_97), .Y(n_1053) );
INVx2_ASAP7_75t_L g1057 ( .A(n_15), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g910 ( .A1(n_16), .A2(n_239), .B1(n_582), .B2(n_901), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_16), .A2(n_21), .B1(n_916), .B2(n_919), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_17), .A2(n_141), .B1(n_1234), .B2(n_1236), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_17), .A2(n_141), .B1(n_445), .B2(n_663), .Y(n_1249) );
OAI22xp5_ASAP7_75t_SL g655 ( .A1(n_18), .A2(n_133), .B1(n_656), .B2(n_657), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_18), .A2(n_133), .B1(n_662), .B2(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g934 ( .A(n_19), .Y(n_934) );
AO22x2_ASAP7_75t_L g532 ( .A1(n_20), .A2(n_533), .B1(n_598), .B2(n_599), .Y(n_532) );
INVx1_ASAP7_75t_L g598 ( .A(n_20), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_21), .A2(n_163), .B1(n_499), .B2(n_905), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_22), .A2(n_204), .B1(n_405), .B2(n_446), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_22), .A2(n_243), .B1(n_386), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g884 ( .A(n_23), .Y(n_884) );
INVx1_ASAP7_75t_L g611 ( .A(n_24), .Y(n_611) );
INVx1_ASAP7_75t_L g767 ( .A(n_25), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_25), .A2(n_215), .B1(n_479), .B2(n_802), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_26), .A2(n_167), .B1(n_1058), .B2(n_1068), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_27), .A2(n_157), .B1(n_1052), .B2(n_1058), .Y(n_1091) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_28), .A2(n_36), .B1(n_261), .B2(n_750), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_28), .A2(n_36), .B1(n_989), .B2(n_1245), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_29), .A2(n_155), .B1(n_261), .B2(n_395), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_29), .A2(n_155), .B1(n_406), .B2(n_938), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_30), .A2(n_184), .B1(n_1048), .B2(n_1055), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_31), .A2(n_129), .B1(n_386), .B2(n_850), .Y(n_863) );
OAI22xp33_ASAP7_75t_SL g865 ( .A1(n_31), .A2(n_129), .B1(n_405), .B2(n_590), .Y(n_865) );
INVx1_ASAP7_75t_L g540 ( .A(n_32), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_33), .A2(n_186), .B1(n_386), .B2(n_388), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_33), .A2(n_91), .B1(n_405), .B2(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g1263 ( .A(n_34), .Y(n_1263) );
INVx1_ASAP7_75t_L g1015 ( .A(n_35), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_37), .A2(n_154), .B1(n_261), .B2(n_395), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_37), .A2(n_154), .B1(n_673), .B2(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g716 ( .A(n_38), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_39), .A2(n_102), .B1(n_1048), .B2(n_1055), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_40), .A2(n_115), .B1(n_585), .B2(n_848), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_40), .A2(n_51), .B1(n_406), .B2(n_427), .Y(n_961) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_41), .B(n_897), .Y(n_896) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_42), .B(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_42), .A2(n_94), .B1(n_1048), .B2(n_1055), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_43), .A2(n_193), .B1(n_1048), .B2(n_1058), .Y(n_1080) );
INVx1_ASAP7_75t_L g930 ( .A(n_44), .Y(n_930) );
INVx1_ASAP7_75t_L g861 ( .A(n_45), .Y(n_861) );
INVx1_ASAP7_75t_L g1260 ( .A(n_46), .Y(n_1260) );
INVx1_ASAP7_75t_L g294 ( .A(n_47), .Y(n_294) );
INVx1_ASAP7_75t_L g301 ( .A(n_47), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_48), .A2(n_124), .B1(n_675), .B2(n_989), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_48), .A2(n_124), .B1(n_261), .B2(n_395), .Y(n_1010) );
INVx1_ASAP7_75t_L g770 ( .A(n_49), .Y(n_770) );
XOR2xp5_ASAP7_75t_L g804 ( .A(n_50), .B(n_805), .Y(n_804) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_51), .A2(n_191), .B1(n_386), .B2(n_850), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_52), .A2(n_99), .B1(n_585), .B2(n_586), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_52), .A2(n_99), .B1(n_426), .B2(n_427), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g1294 ( .A(n_53), .B(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1303 ( .A(n_54), .Y(n_1303) );
INVx1_ASAP7_75t_L g1309 ( .A(n_55), .Y(n_1309) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_56), .A2(n_368), .B(n_369), .C(n_375), .Y(n_367) );
INVx1_ASAP7_75t_L g424 ( .A(n_56), .Y(n_424) );
INVx1_ASAP7_75t_L g253 ( .A(n_57), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_58), .A2(n_183), .B1(n_462), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_58), .A2(n_192), .B1(n_502), .B2(n_506), .Y(n_508) );
INVx2_ASAP7_75t_L g287 ( .A(n_59), .Y(n_287) );
INVx1_ASAP7_75t_L g619 ( .A(n_60), .Y(n_619) );
INVx1_ASAP7_75t_L g810 ( .A(n_61), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_62), .A2(n_79), .B1(n_1055), .B2(n_1068), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_63), .A2(n_210), .B1(n_520), .B2(n_657), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_63), .A2(n_210), .B1(n_683), .B2(n_997), .Y(n_1333) );
INVx1_ASAP7_75t_L g953 ( .A(n_64), .Y(n_953) );
INVx1_ASAP7_75t_L g1270 ( .A(n_65), .Y(n_1270) );
OAI222xp33_ASAP7_75t_L g448 ( .A1(n_66), .A2(n_100), .B1(n_221), .B2(n_449), .C1(n_451), .C2(n_453), .Y(n_448) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_66), .A2(n_100), .B1(n_221), .B2(n_524), .C1(n_526), .C2(n_528), .Y(n_523) );
INVx1_ASAP7_75t_L g968 ( .A(n_67), .Y(n_968) );
INVx1_ASAP7_75t_L g723 ( .A(n_68), .Y(n_723) );
INVx1_ASAP7_75t_L g1304 ( .A(n_69), .Y(n_1304) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_70), .A2(n_91), .B1(n_392), .B2(n_395), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_70), .A2(n_186), .B1(n_426), .B2(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g879 ( .A(n_71), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_72), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_73), .A2(n_246), .B1(n_471), .B2(n_473), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_73), .A2(n_122), .B1(n_513), .B2(n_514), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_74), .A2(n_122), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_74), .A2(n_246), .B1(n_502), .B2(n_506), .Y(n_501) );
XOR2xp5_ASAP7_75t_L g746 ( .A(n_75), .B(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_75), .A2(n_117), .B1(n_1048), .B2(n_1055), .Y(n_1076) );
INVx1_ASAP7_75t_L g860 ( .A(n_76), .Y(n_860) );
INVx1_ASAP7_75t_L g1242 ( .A(n_77), .Y(n_1242) );
OAI211xp5_ASAP7_75t_L g1246 ( .A1(n_77), .A2(n_451), .B(n_592), .C(n_1247), .Y(n_1246) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_78), .A2(n_200), .B1(n_499), .B2(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_78), .A2(n_80), .B1(n_563), .B2(n_922), .Y(n_921) );
XOR2x2_ASAP7_75t_L g1230 ( .A(n_79), .B(n_1231), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_79), .A2(n_1291), .B1(n_1293), .B2(n_1334), .Y(n_1290) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_80), .A2(n_152), .B1(n_582), .B2(n_901), .Y(n_900) );
XOR2x2_ASAP7_75t_L g854 ( .A(n_81), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g1300 ( .A(n_82), .Y(n_1300) );
OAI211xp5_ASAP7_75t_L g1322 ( .A1(n_83), .A2(n_647), .B(n_1323), .C(n_1326), .Y(n_1322) );
INVx1_ASAP7_75t_L g1332 ( .A(n_83), .Y(n_1332) );
INVx1_ASAP7_75t_L g624 ( .A(n_84), .Y(n_624) );
INVx1_ASAP7_75t_L g276 ( .A(n_85), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_85), .A2(n_116), .B1(n_1048), .B2(n_1055), .Y(n_1085) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_86), .A2(n_243), .B1(n_406), .B2(n_426), .C(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g846 ( .A(n_86), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_87), .A2(n_153), .B1(n_585), .B2(n_848), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_87), .A2(n_153), .B1(n_426), .B2(n_427), .Y(n_872) );
INVx1_ASAP7_75t_L g1020 ( .A(n_88), .Y(n_1020) );
AOI22xp5_ASAP7_75t_SL g1084 ( .A1(n_89), .A2(n_234), .B1(n_1058), .B2(n_1068), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_90), .Y(n_255) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_90), .B(n_253), .Y(n_1049) );
OAI211xp5_ASAP7_75t_L g749 ( .A1(n_92), .A2(n_750), .B(n_751), .C(n_759), .Y(n_749) );
INVx1_ASAP7_75t_L g792 ( .A(n_92), .Y(n_792) );
INVx1_ASAP7_75t_L g812 ( .A(n_93), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g1064 ( .A1(n_95), .A2(n_104), .B1(n_1052), .B2(n_1058), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_96), .A2(n_158), .B1(n_663), .B2(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_96), .A2(n_158), .B1(n_520), .B2(n_657), .Y(n_699) );
INVx1_ASAP7_75t_L g1051 ( .A(n_97), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_97), .B(n_1057), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_98), .A2(n_244), .B1(n_1048), .B2(n_1052), .Y(n_1047) );
INVx1_ASAP7_75t_L g813 ( .A(n_101), .Y(n_813) );
INVx1_ASAP7_75t_L g557 ( .A(n_103), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_105), .A2(n_213), .B1(n_445), .B2(n_446), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_105), .A2(n_213), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g286 ( .A(n_106), .Y(n_286) );
INVx1_ASAP7_75t_L g334 ( .A(n_106), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_107), .Y(n_295) );
INVx1_ASAP7_75t_L g689 ( .A(n_108), .Y(n_689) );
INVx1_ASAP7_75t_L g971 ( .A(n_109), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_110), .A2(n_220), .B1(n_1048), .B2(n_1055), .Y(n_1069) );
INVx1_ASAP7_75t_L g877 ( .A(n_111), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_112), .Y(n_310) );
INVx1_ASAP7_75t_L g652 ( .A(n_113), .Y(n_652) );
INVx1_ASAP7_75t_L g439 ( .A(n_114), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g956 ( .A1(n_115), .A2(n_191), .B1(n_405), .B2(n_426), .Y(n_956) );
INVx1_ASAP7_75t_L g1028 ( .A(n_118), .Y(n_1028) );
INVx1_ASAP7_75t_L g974 ( .A(n_119), .Y(n_974) );
INVx1_ASAP7_75t_L g578 ( .A(n_120), .Y(n_578) );
INVx1_ASAP7_75t_L g886 ( .A(n_121), .Y(n_886) );
INVx1_ASAP7_75t_L g708 ( .A(n_123), .Y(n_708) );
XOR2xp5_ASAP7_75t_L g435 ( .A(n_125), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g714 ( .A(n_126), .Y(n_714) );
INVx1_ASAP7_75t_L g1269 ( .A(n_127), .Y(n_1269) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_128), .A2(n_229), .B1(n_1058), .B2(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g758 ( .A(n_130), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_130), .A2(n_209), .B1(n_426), .B2(n_427), .Y(n_790) );
INVx1_ASAP7_75t_L g972 ( .A(n_131), .Y(n_972) );
INVx1_ASAP7_75t_L g555 ( .A(n_132), .Y(n_555) );
INVx1_ASAP7_75t_L g752 ( .A(n_134), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_135), .Y(n_772) );
BUFx3_ASAP7_75t_L g292 ( .A(n_136), .Y(n_292) );
INVx1_ASAP7_75t_L g966 ( .A(n_137), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_138), .Y(n_327) );
INVx1_ASAP7_75t_L g1014 ( .A(n_139), .Y(n_1014) );
INVx1_ASAP7_75t_L g1301 ( .A(n_140), .Y(n_1301) );
INVx1_ASAP7_75t_L g654 ( .A(n_142), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_142), .A2(n_592), .B(n_665), .C(n_667), .Y(n_664) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_143), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_144), .A2(n_192), .B1(n_462), .B2(n_468), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_144), .A2(n_183), .B1(n_494), .B2(n_498), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_145), .A2(n_189), .B1(n_673), .B2(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_145), .A2(n_189), .B1(n_386), .B2(n_395), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_146), .Y(n_765) );
INVx1_ASAP7_75t_L g835 ( .A(n_147), .Y(n_835) );
INVx1_ASAP7_75t_L g552 ( .A(n_148), .Y(n_552) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_149), .B(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1018 ( .A(n_150), .Y(n_1018) );
INVx1_ASAP7_75t_L g543 ( .A(n_151), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_152), .A2(n_200), .B1(n_913), .B2(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g994 ( .A(n_156), .Y(n_994) );
INVx1_ASAP7_75t_L g1307 ( .A(n_159), .Y(n_1307) );
OA22x2_ASAP7_75t_L g679 ( .A1(n_160), .A2(n_680), .B1(n_738), .B2(n_739), .Y(n_679) );
INVxp67_ASAP7_75t_L g739 ( .A(n_160), .Y(n_739) );
INVx1_ASAP7_75t_L g1253 ( .A(n_162), .Y(n_1253) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_163), .A2(n_239), .B1(n_916), .B2(n_919), .Y(n_915) );
INVx1_ASAP7_75t_L g821 ( .A(n_164), .Y(n_821) );
INVx1_ASAP7_75t_L g1241 ( .A(n_165), .Y(n_1241) );
INVx1_ASAP7_75t_L g932 ( .A(n_166), .Y(n_932) );
INVx1_ASAP7_75t_L g763 ( .A(n_168), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_168), .B(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_169), .A2(n_177), .B1(n_1052), .B2(n_1058), .Y(n_1112) );
INVx1_ASAP7_75t_L g629 ( .A(n_170), .Y(n_629) );
INVx1_ASAP7_75t_L g976 ( .A(n_171), .Y(n_976) );
INVx1_ASAP7_75t_L g705 ( .A(n_172), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_173), .B(n_420), .Y(n_834) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_173), .Y(n_841) );
INVx1_ASAP7_75t_L g580 ( .A(n_174), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_175), .A2(n_413), .B(n_685), .C(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g697 ( .A(n_175), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g991 ( .A1(n_176), .A2(n_592), .B(n_992), .C(n_993), .Y(n_991) );
INVx1_ASAP7_75t_L g1006 ( .A(n_176), .Y(n_1006) );
INVx1_ASAP7_75t_L g1256 ( .A(n_178), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_179), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_180), .A2(n_237), .B1(n_683), .B2(n_997), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_180), .A2(n_237), .B1(n_656), .B2(n_1008), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
INVx1_ASAP7_75t_L g933 ( .A(n_182), .Y(n_933) );
INVx1_ASAP7_75t_L g626 ( .A(n_185), .Y(n_626) );
INVx1_ASAP7_75t_L g544 ( .A(n_187), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_188), .Y(n_289) );
INVx1_ASAP7_75t_L g952 ( .A(n_190), .Y(n_952) );
INVx1_ASAP7_75t_L g816 ( .A(n_195), .Y(n_816) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_197), .A2(n_647), .B(n_650), .C(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_197), .Y(n_670) );
INVx1_ASAP7_75t_L g883 ( .A(n_198), .Y(n_883) );
INVx1_ASAP7_75t_L g537 ( .A(n_199), .Y(n_537) );
INVx1_ASAP7_75t_L g1325 ( .A(n_201), .Y(n_1325) );
OAI211xp5_ASAP7_75t_L g1330 ( .A1(n_201), .A2(n_592), .B(n_992), .C(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g969 ( .A(n_202), .Y(n_969) );
INVx1_ASAP7_75t_L g550 ( .A(n_203), .Y(n_550) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_204), .Y(n_843) );
INVx1_ASAP7_75t_L g929 ( .A(n_205), .Y(n_929) );
INVx1_ASAP7_75t_L g722 ( .A(n_206), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_207), .Y(n_378) );
INVx1_ASAP7_75t_L g880 ( .A(n_208), .Y(n_880) );
INVx1_ASAP7_75t_L g760 ( .A(n_209), .Y(n_760) );
BUFx3_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
INVx1_ASAP7_75t_L g394 ( .A(n_211), .Y(n_394) );
INVx1_ASAP7_75t_L g1324 ( .A(n_212), .Y(n_1324) );
XOR2x2_ASAP7_75t_L g985 ( .A(n_214), .B(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g809 ( .A(n_216), .Y(n_809) );
INVx1_ASAP7_75t_L g1261 ( .A(n_217), .Y(n_1261) );
INVx1_ASAP7_75t_L g717 ( .A(n_218), .Y(n_717) );
INVx1_ASAP7_75t_L g712 ( .A(n_219), .Y(n_712) );
INVx1_ASAP7_75t_L g876 ( .A(n_222), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_223), .Y(n_320) );
INVx1_ASAP7_75t_L g583 ( .A(n_224), .Y(n_583) );
INVx1_ASAP7_75t_L g1025 ( .A(n_225), .Y(n_1025) );
OAI211xp5_ASAP7_75t_L g857 ( .A1(n_226), .A2(n_369), .B(n_858), .C(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g868 ( .A(n_226), .Y(n_868) );
INVx1_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
INVx2_ASAP7_75t_L g332 ( .A(n_227), .Y(n_332) );
INVx1_ASAP7_75t_L g488 ( .A(n_227), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_228), .A2(n_230), .B1(n_1055), .B2(n_1058), .Y(n_1054) );
INVx1_ASAP7_75t_L g820 ( .A(n_231), .Y(n_820) );
INVx1_ASAP7_75t_L g609 ( .A(n_232), .Y(n_609) );
INVx1_ASAP7_75t_L g1310 ( .A(n_233), .Y(n_1310) );
INVx1_ASAP7_75t_L g615 ( .A(n_235), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_236), .A2(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g795 ( .A(n_236), .Y(n_795) );
INVx1_ASAP7_75t_L g1027 ( .A(n_238), .Y(n_1027) );
INVx1_ASAP7_75t_L g995 ( .A(n_240), .Y(n_995) );
OAI211xp5_ASAP7_75t_L g1000 ( .A1(n_240), .A2(n_650), .B(n_1001), .C(n_1004), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_241), .Y(n_329) );
INVx1_ASAP7_75t_L g441 ( .A(n_242), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_245), .Y(n_756) );
INVx1_ASAP7_75t_L g1306 ( .A(n_247), .Y(n_1306) );
INVx1_ASAP7_75t_L g384 ( .A(n_248), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_248), .A2(n_410), .B(n_413), .C(n_417), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1041), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1289 ( .A(n_251), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_252), .B(n_255), .Y(n_1292) );
INVx1_ASAP7_75t_L g1335 ( .A(n_252), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_255), .B(n_1335), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g400 ( .A(n_258), .B(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_SL g748 ( .A1(n_258), .A2(n_749), .B(n_761), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_258), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g365 ( .A(n_259), .B(n_269), .Y(n_365) );
AND2x4_ASAP7_75t_L g778 ( .A(n_259), .B(n_268), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_260), .A2(n_396), .B1(n_439), .B2(n_441), .Y(n_517) );
AND2x4_ASAP7_75t_SL g1287 ( .A(n_260), .B(n_1288), .Y(n_1287) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
OR2x6_ASAP7_75t_L g392 ( .A(n_262), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g585 ( .A(n_262), .B(n_393), .Y(n_585) );
BUFx4f_ASAP7_75t_L g764 ( .A(n_262), .Y(n_764) );
INVx1_ASAP7_75t_L g895 ( .A(n_262), .Y(n_895) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_263), .Y(n_342) );
INVx3_ASAP7_75t_L g387 ( .A(n_263), .Y(n_387) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
INVx2_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
NAND2x1_ASAP7_75t_L g357 ( .A(n_265), .B(n_266), .Y(n_357) );
AND2x2_ASAP7_75t_L g374 ( .A(n_265), .B(n_266), .Y(n_374) );
INVx1_ASAP7_75t_L g383 ( .A(n_265), .Y(n_383) );
AND2x2_ASAP7_75t_L g397 ( .A(n_265), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_266), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g352 ( .A(n_266), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g377 ( .A(n_266), .Y(n_377) );
INVx2_ASAP7_75t_L g398 ( .A(n_266), .Y(n_398) );
INVx1_ASAP7_75t_L g497 ( .A(n_266), .Y(n_497) );
AND2x2_ASAP7_75t_L g500 ( .A(n_266), .B(n_348), .Y(n_500) );
OR2x6_ASAP7_75t_L g386 ( .A(n_267), .B(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_267), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g371 ( .A(n_268), .Y(n_371) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g381 ( .A(n_269), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g390 ( .A(n_269), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_741), .B2(n_742), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AO22x1_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_433), .B2(n_740), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
XNOR2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND3x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_366), .C(n_403), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_336), .Y(n_278) );
OAI33xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_288), .A3(n_303), .B1(n_315), .B2(n_324), .B3(n_330), .Y(n_279) );
OAI33xp33_ASAP7_75t_L g874 ( .A1(n_280), .A2(n_330), .A3(n_875), .B1(n_878), .B2(n_881), .B3(n_885), .Y(n_874) );
OAI33xp33_ASAP7_75t_L g977 ( .A1(n_280), .A2(n_330), .A3(n_978), .B1(n_979), .B2(n_981), .B3(n_983), .Y(n_977) );
BUFx4f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g559 ( .A(n_281), .Y(n_559) );
BUFx4f_ASAP7_75t_L g1272 ( .A(n_281), .Y(n_1272) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_282), .B(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_282), .Y(n_432) );
INVx1_ASAP7_75t_L g511 ( .A(n_282), .Y(n_511) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g402 ( .A(n_283), .Y(n_402) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_287), .Y(n_285) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_286), .Y(n_430) );
AND3x4_ASAP7_75t_L g459 ( .A(n_286), .B(n_420), .C(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
BUFx3_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B1(n_295), .B2(n_296), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_289), .A2(n_327), .B1(n_341), .B2(n_343), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_290), .A2(n_296), .B1(n_543), .B2(n_555), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_290), .A2(n_328), .B1(n_544), .B2(n_557), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_290), .A2(n_787), .B1(n_809), .B2(n_810), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_290), .A2(n_687), .B1(n_820), .B2(n_821), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_290), .A2(n_687), .B1(n_876), .B2(n_877), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_290), .A2(n_328), .B1(n_886), .B2(n_887), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_290), .A2(n_966), .B1(n_972), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1275 ( .A(n_290), .Y(n_1275) );
BUFx4f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
OR2x4_ASAP7_75t_L g405 ( .A(n_291), .B(n_335), .Y(n_405) );
OR2x4_ASAP7_75t_L g426 ( .A(n_291), .B(n_408), .Y(n_426) );
BUFx3_ASAP7_75t_L g634 ( .A(n_291), .Y(n_634) );
BUFx3_ASAP7_75t_L g728 ( .A(n_291), .Y(n_728) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_292), .Y(n_302) );
INVx2_ASAP7_75t_L g309 ( .A(n_292), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_292), .B(n_301), .Y(n_314) );
AND2x4_ASAP7_75t_L g415 ( .A(n_292), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g467 ( .A(n_293), .Y(n_467) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_295), .A2(n_329), .B1(n_359), .B2(n_360), .Y(n_358) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g1016 ( .A(n_297), .Y(n_1016) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g452 ( .A(n_298), .Y(n_452) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_298), .Y(n_635) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_298), .Y(n_687) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
BUFx2_ASAP7_75t_L g412 ( .A(n_299), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
BUFx2_ASAP7_75t_L g423 ( .A(n_300), .Y(n_423) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g416 ( .A(n_301), .Y(n_416) );
BUFx2_ASAP7_75t_L g421 ( .A(n_302), .Y(n_421) );
AND2x4_ASAP7_75t_L g475 ( .A(n_302), .B(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_310), .B2(n_311), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_304), .A2(n_316), .B1(n_350), .B2(n_354), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_305), .A2(n_969), .B1(n_976), .B2(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g407 ( .A(n_306), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g442 ( .A(n_306), .B(n_408), .Y(n_442) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_306), .Y(n_638) );
INVx2_ASAP7_75t_L g641 ( .A(n_306), .Y(n_641) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_306), .Y(n_732) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_307), .Y(n_563) );
BUFx8_ASAP7_75t_L g566 ( .A(n_307), .Y(n_566) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x4_ASAP7_75t_L g466 ( .A(n_309), .B(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_310), .A2(n_320), .B1(n_341), .B2(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_311), .A2(n_968), .B1(n_974), .B2(n_980), .Y(n_979) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
CKINVDCx8_ASAP7_75t_R g733 ( .A(n_312), .Y(n_733) );
INVx3_ASAP7_75t_L g817 ( .A(n_312), .Y(n_817) );
INVx3_ASAP7_75t_L g982 ( .A(n_312), .Y(n_982) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g569 ( .A(n_313), .Y(n_569) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g323 ( .A(n_314), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_320), .B2(n_321), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g735 ( .A(n_318), .Y(n_735) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g472 ( .A(n_319), .Y(n_472) );
INVx1_ASAP7_75t_L g481 ( .A(n_319), .Y(n_481) );
BUFx2_ASAP7_75t_L g800 ( .A(n_319), .Y(n_800) );
OAI22xp33_ASAP7_75t_SL g561 ( .A1(n_321), .A2(n_537), .B1(n_550), .B2(n_562), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_321), .A2(n_565), .B1(n_879), .B2(n_880), .Y(n_878) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g427 ( .A(n_323), .B(n_335), .Y(n_427) );
BUFx3_ASAP7_75t_L g639 ( .A(n_323), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_328), .B2(n_329), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_325), .A2(n_328), .B1(n_965), .B2(n_971), .Y(n_978) );
INVx2_ASAP7_75t_SL g1284 ( .A(n_325), .Y(n_1284) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g1277 ( .A(n_328), .Y(n_1277) );
BUFx6f_ASAP7_75t_L g1285 ( .A(n_328), .Y(n_1285) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
AND2x4_ASAP7_75t_L g338 ( .A(n_331), .B(n_339), .Y(n_338) );
OR2x6_ASAP7_75t_L g570 ( .A(n_331), .B(n_333), .Y(n_570) );
INVx1_ASAP7_75t_L g782 ( .A(n_331), .Y(n_782) );
BUFx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g460 ( .A(n_332), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND3x1_ASAP7_75t_L g486 ( .A(n_334), .B(n_335), .C(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g408 ( .A(n_335), .Y(n_408) );
AND2x4_ASAP7_75t_L g414 ( .A(n_335), .B(n_415), .Y(n_414) );
OAI33xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .A3(n_349), .B1(n_358), .B2(n_361), .B3(n_363), .Y(n_336) );
OAI33xp33_ASAP7_75t_L g822 ( .A1(n_337), .A2(n_823), .A3(n_824), .B1(n_826), .B2(n_827), .B3(n_829), .Y(n_822) );
OAI33xp33_ASAP7_75t_L g888 ( .A1(n_337), .A2(n_829), .A3(n_889), .B1(n_891), .B2(n_892), .B3(n_893), .Y(n_888) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g492 ( .A(n_338), .Y(n_492) );
INVx4_ASAP7_75t_L g548 ( .A(n_338), .Y(n_548) );
INVx2_ASAP7_75t_L g710 ( .A(n_338), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_341), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_341), .A2(n_876), .B1(n_886), .B2(n_890), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_341), .A2(n_343), .B1(n_965), .B2(n_966), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_341), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
INVx4_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_342), .Y(n_707) );
INVx3_ASAP7_75t_L g1033 ( .A(n_342), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_343), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_343), .A2(n_813), .B1(n_818), .B2(n_828), .Y(n_827) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
INVx1_ASAP7_75t_L g545 ( .A(n_345), .Y(n_545) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_345), .Y(n_613) );
INVx1_ASAP7_75t_L g890 ( .A(n_345), .Y(n_890) );
INVx2_ASAP7_75t_SL g975 ( .A(n_345), .Y(n_975) );
INVx8_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g389 ( .A(n_346), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g848 ( .A(n_346), .B(n_371), .Y(n_848) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_350), .A2(n_541), .B1(n_968), .B2(n_969), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_350), .A2(n_556), .B1(n_971), .B2(n_972), .Y(n_970) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g623 ( .A(n_351), .Y(n_623) );
BUFx2_ASAP7_75t_L g769 ( .A(n_351), .Y(n_769) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g359 ( .A(n_352), .Y(n_359) );
INVx1_ASAP7_75t_L g539 ( .A(n_352), .Y(n_539) );
BUFx3_ASAP7_75t_L g554 ( .A(n_352), .Y(n_554) );
BUFx2_ASAP7_75t_L g618 ( .A(n_352), .Y(n_618) );
AND2x2_ASAP7_75t_L g496 ( .A(n_353), .B(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_354), .A2(n_538), .B1(n_879), .B2(n_883), .Y(n_891) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_355), .Y(n_368) );
INVx1_ASAP7_75t_L g695 ( .A(n_355), .Y(n_695) );
INVx2_ASAP7_75t_L g1035 ( .A(n_355), .Y(n_1035) );
INVx4_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_356), .Y(n_541) );
BUFx4f_ASAP7_75t_L g556 ( .A(n_356), .Y(n_556) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_356), .Y(n_649) );
BUFx4f_ASAP7_75t_L g773 ( .A(n_356), .Y(n_773) );
BUFx4f_ASAP7_75t_L g825 ( .A(n_356), .Y(n_825) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g360 ( .A(n_357), .Y(n_360) );
INVx2_ASAP7_75t_SL g527 ( .A(n_360), .Y(n_527) );
BUFx2_ASAP7_75t_SL g625 ( .A(n_360), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_360), .A2(n_538), .B1(n_877), .B2(n_887), .Y(n_892) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_360), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_360), .A2(n_623), .B1(n_1303), .B2(n_1304), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_362), .A2(n_551), .B1(n_809), .B2(n_820), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_362), .A2(n_880), .B1(n_884), .B2(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g1258 ( .A(n_362), .Y(n_1258) );
OAI33xp33_ASAP7_75t_L g535 ( .A1(n_363), .A2(n_536), .A3(n_542), .B1(n_546), .B2(n_549), .B3(n_553), .Y(n_535) );
OAI33xp33_ASAP7_75t_L g963 ( .A1(n_363), .A2(n_492), .A3(n_964), .B1(n_967), .B2(n_970), .B3(n_973), .Y(n_963) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g829 ( .A(n_364), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_364), .B(n_908), .C(n_910), .Y(n_907) );
AND2x4_ASAP7_75t_L g509 ( .A(n_365), .B(n_510), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_365), .A2(n_695), .B1(n_767), .B2(n_768), .C(n_770), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_365), .B(n_510), .Y(n_1267) );
OAI31xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_385), .A3(n_391), .B(n_399), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_368), .A2(n_768), .B1(n_1015), .B2(n_1028), .Y(n_1036) );
NAND3xp33_ASAP7_75t_SL g839 ( .A(n_369), .B(n_840), .C(n_842), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g927 ( .A(n_369), .B(n_928), .C(n_931), .Y(n_927) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x2_ASAP7_75t_L g376 ( .A(n_371), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g529 ( .A(n_371), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g507 ( .A(n_373), .Y(n_507) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_374), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_379), .B2(n_384), .Y(n_375) );
INVx1_ASAP7_75t_L g754 ( .A(n_376), .Y(n_754) );
AND2x4_ASAP7_75t_L g525 ( .A(n_377), .B(n_390), .Y(n_525) );
AND2x2_ASAP7_75t_L g577 ( .A(n_377), .B(n_390), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_378), .A2(n_418), .B1(n_422), .B2(n_424), .Y(n_417) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g528 ( .A(n_381), .Y(n_528) );
BUFx3_ASAP7_75t_L g579 ( .A(n_381), .Y(n_579) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g551 ( .A(n_387), .Y(n_551) );
BUFx3_ASAP7_75t_L g610 ( .A(n_387), .Y(n_610) );
INVx2_ASAP7_75t_SL g721 ( .A(n_387), .Y(n_721) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_387), .Y(n_828) );
INVx2_ASAP7_75t_SL g1009 ( .A(n_388), .Y(n_1009) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g522 ( .A(n_389), .Y(n_522) );
INVx2_ASAP7_75t_L g587 ( .A(n_389), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_390), .A2(n_582), .B(n_752), .C(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g757 ( .A(n_390), .Y(n_757) );
AND2x2_ASAP7_75t_L g844 ( .A(n_390), .B(n_845), .Y(n_844) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_392), .Y(n_520) );
BUFx2_ASAP7_75t_L g656 ( .A(n_392), .Y(n_656) );
INVx1_ASAP7_75t_L g1235 ( .A(n_392), .Y(n_1235) );
AND2x4_ASAP7_75t_L g396 ( .A(n_393), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_SL g750 ( .A(n_396), .Y(n_750) );
INVx4_ASAP7_75t_L g850 ( .A(n_396), .Y(n_850) );
INVx2_ASAP7_75t_L g505 ( .A(n_397), .Y(n_505) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_397), .Y(n_776) );
BUFx3_ASAP7_75t_L g903 ( .A(n_397), .Y(n_903) );
OAI31xp33_ASAP7_75t_L g572 ( .A1(n_399), .A2(n_573), .A3(n_574), .B(n_584), .Y(n_572) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g531 ( .A(n_400), .Y(n_531) );
BUFx3_ASAP7_75t_L g659 ( .A(n_400), .Y(n_659) );
BUFx2_ASAP7_75t_SL g701 ( .A(n_400), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_400), .A2(n_839), .B(n_849), .Y(n_838) );
OAI31xp33_ASAP7_75t_L g948 ( .A1(n_400), .A2(n_949), .A3(n_950), .B(n_954), .Y(n_948) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI31xp33_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_409), .A3(n_425), .B(n_428), .Y(n_403) );
INVx2_ASAP7_75t_SL g440 ( .A(n_405), .Y(n_440) );
INVx1_ASAP7_75t_L g674 ( .A(n_405), .Y(n_674) );
INVx2_ASAP7_75t_SL g990 ( .A(n_405), .Y(n_990) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_407), .A2(n_674), .B1(n_756), .B2(n_792), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_410), .A2(n_634), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1319 ( .A1(n_410), .A2(n_1301), .B1(n_1307), .B2(n_1313), .Y(n_1319) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g644 ( .A(n_412), .Y(n_644) );
INVx1_ASAP7_75t_L g666 ( .A(n_412), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_413), .B(n_867), .C(n_869), .Y(n_866) );
NAND3xp33_ASAP7_75t_SL g957 ( .A(n_413), .B(n_958), .C(n_959), .Y(n_957) );
CKINVDCx8_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_414), .B(n_444), .C(n_448), .Y(n_443) );
CKINVDCx8_ASAP7_75t_R g592 ( .A(n_414), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_414), .B(n_786), .C(n_790), .Y(n_785) );
INVx2_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
BUFx2_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
BUFx2_ASAP7_75t_L g595 ( .A(n_415), .Y(n_595) );
BUFx2_ASAP7_75t_L g833 ( .A(n_415), .Y(n_833) );
BUFx3_ASAP7_75t_L g871 ( .A(n_415), .Y(n_871) );
BUFx2_ASAP7_75t_L g941 ( .A(n_415), .Y(n_941) );
INVx1_ASAP7_75t_L g476 ( .A(n_416), .Y(n_476) );
INVx1_ASAP7_75t_L g788 ( .A(n_418), .Y(n_788) );
AOI222xp33_ASAP7_75t_L g832 ( .A1(n_418), .A2(n_422), .B1(n_833), .B2(n_834), .C1(n_835), .C2(n_836), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_418), .A2(n_422), .B1(n_952), .B2(n_960), .Y(n_959) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_419), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g450 ( .A(n_419), .B(n_421), .Y(n_450) );
AND2x4_ASAP7_75t_L g454 ( .A(n_419), .B(n_423), .Y(n_454) );
AND2x2_ASAP7_75t_L g669 ( .A(n_419), .B(n_421), .Y(n_669) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g789 ( .A(n_422), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_422), .A2(n_450), .B1(n_860), .B2(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g445 ( .A(n_426), .Y(n_445) );
BUFx2_ASAP7_75t_L g662 ( .A(n_426), .Y(n_662) );
BUFx3_ASAP7_75t_L g683 ( .A(n_426), .Y(n_683) );
INVx2_ASAP7_75t_SL g944 ( .A(n_426), .Y(n_944) );
INVx2_ASAP7_75t_L g447 ( .A(n_427), .Y(n_447) );
BUFx3_ASAP7_75t_L g663 ( .A(n_427), .Y(n_663) );
INVx1_ASAP7_75t_L g998 ( .A(n_427), .Y(n_998) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_428), .A2(n_831), .B(n_837), .Y(n_830) );
OAI31xp33_ASAP7_75t_L g864 ( .A1(n_428), .A2(n_865), .A3(n_866), .B(n_872), .Y(n_864) );
OAI21xp5_ASAP7_75t_L g936 ( .A1(n_428), .A2(n_937), .B(n_939), .Y(n_936) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x4_ASAP7_75t_L g456 ( .A(n_429), .B(n_431), .Y(n_456) );
AND2x2_ASAP7_75t_L g597 ( .A(n_429), .B(n_431), .Y(n_597) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_429), .B(n_431), .Y(n_677) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g740 ( .A(n_433), .Y(n_740) );
XNOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_602), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_532), .B1(n_600), .B2(n_601), .Y(n_434) );
INVx1_ASAP7_75t_L g601 ( .A(n_435), .Y(n_601) );
NAND4xp25_ASAP7_75t_SL g436 ( .A(n_437), .B(n_457), .C(n_489), .D(n_516), .Y(n_436) );
AO21x1_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_443), .B(n_455), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx2_ASAP7_75t_SL g938 ( .A(n_440), .Y(n_938) );
INVx1_ASAP7_75t_L g590 ( .A(n_442), .Y(n_590) );
INVx2_ASAP7_75t_L g675 ( .A(n_442), .Y(n_675) );
INVx1_ASAP7_75t_L g692 ( .A(n_442), .Y(n_692) );
INVx1_ASAP7_75t_L g1245 ( .A(n_442), .Y(n_1245) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_447), .A2(n_929), .B1(n_930), .B2(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_450), .A2(n_454), .B1(n_578), .B2(n_583), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_450), .A2(n_454), .B1(n_689), .B2(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g787 ( .A(n_452), .Y(n_787) );
INVx1_ASAP7_75t_L g984 ( .A(n_452), .Y(n_984) );
INVx2_ASAP7_75t_L g992 ( .A(n_452), .Y(n_992) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_454), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g940 ( .A1(n_454), .A2(n_932), .B1(n_933), .B2(n_934), .C1(n_941), .C2(n_942), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_455), .A2(n_531), .B1(n_1232), .B2(n_1243), .C(n_1250), .Y(n_1231) );
CKINVDCx14_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
OAI31xp33_ASAP7_75t_L g681 ( .A1(n_456), .A2(n_682), .A3(n_684), .B(n_691), .Y(n_681) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .A3(n_470), .B1(n_477), .B2(n_480), .B3(n_483), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g911 ( .A(n_459), .B(n_912), .C(n_915), .Y(n_911) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx8_ASAP7_75t_L g803 ( .A(n_466), .Y(n_803) );
BUFx3_ASAP7_75t_L g918 ( .A(n_466), .Y(n_918) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g919 ( .A(n_469), .Y(n_919) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g482 ( .A(n_474), .Y(n_482) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g798 ( .A(n_475), .Y(n_798) );
BUFx3_ASAP7_75t_L g914 ( .A(n_475), .Y(n_914) );
BUFx12f_ASAP7_75t_L g922 ( .A(n_475), .Y(n_922) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g1279 ( .A(n_481), .Y(n_1279) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_484), .A2(n_559), .A3(n_633), .B1(n_636), .B2(n_640), .B3(n_642), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_484), .A2(n_559), .B1(n_794), .B2(n_799), .Y(n_793) );
OAI33xp33_ASAP7_75t_L g1012 ( .A1(n_484), .A2(n_559), .A3(n_1013), .B1(n_1017), .B2(n_1021), .B3(n_1026), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g736 ( .A(n_485), .Y(n_736) );
INVx2_ASAP7_75t_L g1318 ( .A(n_485), .Y(n_1318) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g924 ( .A(n_486), .Y(n_924) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI33xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .A3(n_501), .B1(n_508), .B2(n_509), .B3(n_512), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_491), .A2(n_608), .A3(n_614), .B1(n_620), .B2(n_627), .B3(n_628), .Y(n_607) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g513 ( .A(n_495), .Y(n_513) );
INVx2_ASAP7_75t_L g780 ( .A(n_495), .Y(n_780) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_496), .Y(n_845) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g515 ( .A(n_500), .Y(n_515) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g627 ( .A(n_509), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_509), .Y(n_718) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AO21x1_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_531), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .C(n_529), .Y(n_518) );
INVx2_ASAP7_75t_L g1237 ( .A(n_521), .Y(n_1237) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_522), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g653 ( .A(n_525), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_525), .A2(n_579), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI222xp33_ASAP7_75t_L g931 ( .A1(n_525), .A2(n_579), .B1(n_582), .B2(n_932), .C1(n_933), .C2(n_934), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_525), .A2(n_579), .B1(n_952), .B2(n_953), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_526), .A2(n_615), .B1(n_616), .B2(n_619), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_526), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g1262 ( .A1(n_526), .A2(n_623), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
INVx5_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g698 ( .A(n_528), .Y(n_698) );
INVx2_ASAP7_75t_L g1005 ( .A(n_528), .Y(n_1005) );
INVx3_ASAP7_75t_L g575 ( .A(n_529), .Y(n_575) );
INVx1_ASAP7_75t_L g650 ( .A(n_529), .Y(n_650) );
INVx1_ASAP7_75t_L g1326 ( .A(n_529), .Y(n_1326) );
BUFx3_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
INVx3_ASAP7_75t_SL g600 ( .A(n_532), .Y(n_600) );
INVx1_ASAP7_75t_L g599 ( .A(n_533), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_572), .C(n_588), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_558), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B1(n_540), .B2(n_541), .Y(n_536) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g713 ( .A(n_539), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_540), .A2(n_552), .B1(n_565), .B2(n_567), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_541), .A2(n_713), .B1(n_810), .B2(n_821), .Y(n_826) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_541), .Y(n_858) );
BUFx3_ASAP7_75t_L g630 ( .A(n_545), .Y(n_630) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_547), .B(n_900), .C(n_904), .Y(n_899) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g1255 ( .A(n_551), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_554), .A2(n_812), .B1(n_816), .B2(n_825), .Y(n_824) );
OAI33xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .A3(n_561), .B1(n_564), .B2(n_570), .B3(n_571), .Y(n_558) );
OAI33xp33_ASAP7_75t_L g724 ( .A1(n_559), .A2(n_725), .A3(n_730), .B1(n_734), .B2(n_736), .B3(n_737), .Y(n_724) );
OAI33xp33_ASAP7_75t_L g807 ( .A1(n_559), .A2(n_570), .A3(n_808), .B1(n_811), .B2(n_815), .B3(n_819), .Y(n_807) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_562), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_562), .A2(n_733), .B1(n_1303), .B2(n_1309), .Y(n_1315) );
INVx5_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_563), .Y(n_913) );
INVx3_ASAP7_75t_L g980 ( .A(n_563), .Y(n_980) );
INVx2_ASAP7_75t_SL g1317 ( .A(n_563), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_565), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g882 ( .A(n_566), .Y(n_882) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g814 ( .A(n_569), .Y(n_814) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .C(n_581), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_577), .A2(n_689), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI222xp33_ASAP7_75t_L g840 ( .A1(n_577), .A2(n_579), .B1(n_582), .B2(n_835), .C1(n_836), .C2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_577), .A2(n_994), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_579), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_579), .A2(n_653), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_580), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g657 ( .A(n_587), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_587), .A2(n_844), .B1(n_929), .B2(n_930), .Y(n_928) );
OAI31xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .A3(n_596), .B(n_597), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .C(n_594), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_592), .B(n_940), .C(n_943), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_595), .B(n_953), .Y(n_958) );
OAI31xp33_ASAP7_75t_SL g955 ( .A1(n_597), .A2(n_956), .A3(n_957), .B(n_961), .Y(n_955) );
OA22x2_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_678), .B2(n_679), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_645), .C(n_660), .Y(n_605) );
NOR2xp33_ASAP7_75t_SL g606 ( .A(n_607), .B(n_632), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_609), .A2(n_624), .B1(n_634), .B2(n_635), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_610), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_610), .A2(n_612), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_611), .A2(n_626), .B1(n_634), .B2(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_612), .A2(n_1014), .B1(n_1027), .B2(n_1031), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_612), .A2(n_1020), .B1(n_1025), .B2(n_1031), .Y(n_1037) );
OAI22xp5_ASAP7_75t_SL g1299 ( .A1(n_612), .A2(n_1033), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
INVx6_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx5_ASAP7_75t_L g709 ( .A(n_613), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_615), .A2(n_629), .B1(n_637), .B2(n_639), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_616), .A2(n_625), .B1(n_1306), .B2(n_1307), .Y(n_1305) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx4_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_619), .A2(n_631), .B1(n_639), .B2(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_623), .A2(n_825), .B1(n_1260), .B2(n_1261), .Y(n_1259) );
OAI33xp33_ASAP7_75t_L g1298 ( .A1(n_627), .A2(n_710), .A3(n_1299), .B1(n_1302), .B2(n_1305), .B3(n_1308), .Y(n_1298) );
OAI22xp33_ASAP7_75t_L g1013 ( .A1(n_634), .A2(n_1014), .B1(n_1015), .B2(n_1016), .Y(n_1013) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_639), .A2(n_714), .B1(n_723), .B2(n_735), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_639), .A2(n_1022), .B1(n_1024), .B2(n_1025), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_639), .A2(n_1304), .B1(n_1310), .B2(n_1317), .Y(n_1316) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_655), .A3(n_658), .B(n_659), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_649), .A2(n_713), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_652), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_653), .A2(n_1005), .B1(n_1324), .B2(n_1325), .Y(n_1323) );
OAI31xp33_ASAP7_75t_L g999 ( .A1(n_659), .A2(n_1000), .A3(n_1007), .B(n_1010), .Y(n_999) );
OAI31xp33_ASAP7_75t_L g1320 ( .A1(n_659), .A2(n_1321), .A3(n_1322), .B(n_1327), .Y(n_1320) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .A3(n_672), .B(n_676), .Y(n_660) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g729 ( .A(n_666), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_668), .A2(n_671), .B1(n_994), .B2(n_995), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_668), .A2(n_671), .B1(n_1324), .B2(n_1332), .Y(n_1331) );
BUFx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g942 ( .A(n_669), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_671), .A2(n_942), .B1(n_1241), .B2(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI31xp33_ASAP7_75t_L g987 ( .A1(n_676), .A2(n_988), .A3(n_991), .B(n_996), .Y(n_987) );
OAI31xp33_ASAP7_75t_L g1328 ( .A1(n_676), .A2(n_1329), .A3(n_1330), .B(n_1333), .Y(n_1328) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_677), .A2(n_784), .B(n_793), .Y(n_783) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g738 ( .A(n_680), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_693), .C(n_702), .Y(n_680) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_687), .A2(n_708), .B1(n_717), .B2(n_726), .Y(n_737) );
OAI31xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .A3(n_700), .B(n_701), .Y(n_693) );
OAI31xp33_ASAP7_75t_SL g856 ( .A1(n_701), .A2(n_857), .A3(n_862), .B(n_863), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_701), .A2(n_927), .B(n_935), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_724), .Y(n_702) );
OAI33xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_710), .A3(n_711), .B1(n_715), .B2(n_718), .B3(n_719), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_708), .B2(n_709), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_705), .A2(n_716), .B1(n_726), .B2(n_729), .Y(n_725) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_709), .A2(n_720), .B1(n_722), .B2(n_723), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_709), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
OAI33xp33_ASAP7_75t_L g1029 ( .A1(n_710), .A2(n_718), .A3(n_1030), .B1(n_1034), .B2(n_1036), .B3(n_1037), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1251 ( .A1(n_710), .A2(n_1252), .A3(n_1259), .B1(n_1262), .B2(n_1265), .B3(n_1268), .Y(n_1251) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_712), .A2(n_722), .B1(n_731), .B2(n_733), .Y(n_730) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_728), .Y(n_1314) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_731), .A2(n_795), .B(n_796), .C(n_797), .Y(n_794) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_733), .A2(n_765), .B1(n_772), .B2(n_800), .C(n_801), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_733), .A2(n_1018), .B1(n_1019), .B2(n_1020), .Y(n_1017) );
OAI33xp33_ASAP7_75t_L g1271 ( .A1(n_736), .A2(n_1272), .A3(n_1273), .B1(n_1278), .B2(n_1280), .B3(n_1282), .Y(n_1271) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_851), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
XOR2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_804), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_781), .B(n_783), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_766), .B(n_771), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_768), .A2(n_1018), .B1(n_1024), .B2(n_1035), .Y(n_1034) );
INVx4_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI211xp5_ASAP7_75t_SL g771 ( .A1(n_772), .A2(n_773), .B(n_774), .C(n_779), .Y(n_771) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_785), .B(n_791), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_800), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_830), .C(n_838), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_822), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_814), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g1278 ( .A1(n_817), .A2(n_1260), .B1(n_1269), .B2(n_1279), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_846), .B2(n_847), .Y(n_842) );
INVx3_ASAP7_75t_L g906 ( .A(n_845), .Y(n_906) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_845), .Y(n_909) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_945), .B2(n_1040), .Y(n_851) );
INVx2_ASAP7_75t_SL g852 ( .A(n_853), .Y(n_852) );
XNOR2x1_ASAP7_75t_L g853 ( .A(n_854), .B(n_896), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_864), .C(n_873), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_861), .B(n_870), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_888), .Y(n_873) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_926), .C(n_936), .Y(n_897) );
AND4x1_ASAP7_75t_L g898 ( .A(n_899), .B(n_907), .C(n_911), .D(n_920), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g1281 ( .A(n_913), .Y(n_1281) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_923), .C(n_925), .Y(n_920) );
BUFx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1040 ( .A(n_945), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_985), .B1(n_1038), .B2(n_1039), .Y(n_945) );
INVx1_ASAP7_75t_L g1038 ( .A(n_946), .Y(n_1038) );
NAND3xp33_ASAP7_75t_SL g947 ( .A(n_948), .B(n_955), .C(n_962), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_977), .Y(n_962) );
INVx2_ASAP7_75t_L g1023 ( .A(n_980), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_982), .A2(n_1261), .B1(n_1270), .B2(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1039 ( .A(n_985), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_999), .C(n_1011), .Y(n_986) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1029), .Y(n_1011) );
INVx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_1033), .Y(n_1032) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1226), .B1(n_1230), .B2(n_1286), .C(n_1290), .Y(n_1041) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1165), .C(n_1202), .Y(n_1042) );
AOI32xp33_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1131), .A3(n_1150), .B1(n_1154), .B2(n_1164), .Y(n_1043) );
AOI211xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1060), .B(n_1095), .C(n_1119), .Y(n_1044) );
OAI311xp33_ASAP7_75t_L g1095 ( .A1(n_1045), .A2(n_1096), .A3(n_1101), .B1(n_1102), .C1(n_1114), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1045), .B(n_1066), .Y(n_1163) );
AOI21xp33_ASAP7_75t_L g1198 ( .A1(n_1045), .A2(n_1199), .B(n_1201), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1045), .B(n_1062), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1045), .B(n_1089), .Y(n_1224) );
INVx3_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1046), .B(n_1104), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1046), .B(n_1066), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1046), .B(n_1134), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1046), .B(n_1100), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1046), .B(n_1115), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1046), .B(n_1130), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1046), .B(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1046), .B(n_1164), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1046), .B(n_1066), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1046), .B(n_1086), .Y(n_1215) );
AND2x4_ASAP7_75t_SL g1046 ( .A(n_1047), .B(n_1054), .Y(n_1046) );
AND2x6_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1049), .B(n_1053), .Y(n_1052) );
AND2x4_ASAP7_75t_L g1055 ( .A(n_1049), .B(n_1056), .Y(n_1055) );
AND2x6_ASAP7_75t_L g1058 ( .A(n_1049), .B(n_1059), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1049), .B(n_1053), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1049), .B(n_1053), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1051), .B(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1052), .Y(n_1229) );
OAI21xp5_ASAP7_75t_L g1334 ( .A1(n_1053), .A2(n_1335), .B(n_1336), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1070), .B1(n_1086), .B2(n_1088), .Y(n_1060) );
A2O1A1Ixp33_ASAP7_75t_L g1146 ( .A1(n_1061), .A2(n_1089), .B(n_1147), .C(n_1148), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1061), .B(n_1121), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1061), .B(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1066), .Y(n_1062) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1063), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1063), .B(n_1066), .Y(n_1100) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1063), .Y(n_1105) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1063), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_1066), .B(n_1105), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1066), .B(n_1158), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1069), .Y(n_1066) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1067), .B(n_1069), .Y(n_1122) );
AOI31xp33_ASAP7_75t_L g1172 ( .A1(n_1070), .A2(n_1168), .A3(n_1170), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1179 ( .A1(n_1071), .A2(n_1180), .B(n_1182), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1077), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1072), .B(n_1117), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1072), .B(n_1094), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1072), .B(n_1141), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1072), .B(n_1149), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1072), .B(n_1171), .Y(n_1170) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_1073), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1073), .B(n_1094), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1073), .B(n_1079), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1073), .B(n_1078), .Y(n_1109) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_1073), .B(n_1089), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1073), .B(n_1149), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1073), .B(n_1089), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1076), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1074), .B(n_1076), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1077), .B(n_1098), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1077), .B(n_1135), .Y(n_1160) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1077), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1082), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1079), .B(n_1082), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1079), .B(n_1082), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1079), .B(n_1083), .Y(n_1149) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1079), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .Y(n_1079) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1082), .Y(n_1094) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1083), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1086), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1086), .B(n_1190), .Y(n_1200) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1092), .Y(n_1088) );
INVx3_ASAP7_75t_L g1099 ( .A(n_1089), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1089), .B(n_1105), .Y(n_1104) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1089), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .Y(n_1089) );
OAI332xp33_ASAP7_75t_L g1217 ( .A1(n_1092), .A2(n_1133), .A3(n_1196), .B1(n_1218), .B2(n_1221), .B3(n_1222), .C1(n_1223), .C2(n_1225), .Y(n_1217) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1093), .B(n_1098), .Y(n_1181) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1100), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1098), .B(n_1128), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1098), .B(n_1106), .Y(n_1204) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1099), .B(n_1118), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1099), .B(n_1129), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1099), .B(n_1160), .Y(n_1216) );
CKINVDCx14_ASAP7_75t_R g1125 ( .A(n_1100), .Y(n_1125) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1101), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_1103), .A2(n_1106), .B1(n_1107), .B2(n_1109), .C(n_1110), .Y(n_1102) );
CKINVDCx14_ASAP7_75t_R g1184 ( .A(n_1104), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1105), .B(n_1122), .Y(n_1194) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1192 ( .A1(n_1108), .A2(n_1120), .B1(n_1193), .B2(n_1196), .C(n_1197), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1109), .B(n_1121), .Y(n_1120) );
CKINVDCx14_ASAP7_75t_R g1225 ( .A(n_1109), .Y(n_1225) );
OAI31xp33_ASAP7_75t_L g1166 ( .A1(n_1110), .A2(n_1167), .A3(n_1172), .B(n_1175), .Y(n_1166) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1111), .Y(n_1164) );
AOI21xp33_ASAP7_75t_SL g1212 ( .A1(n_1111), .A2(n_1213), .B(n_1214), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1115), .Y(n_1128) );
A2O1A1Ixp33_ASAP7_75t_SL g1154 ( .A1(n_1115), .A2(n_1155), .B(n_1157), .C(n_1163), .Y(n_1154) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1116), .Y(n_1201) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1118), .Y(n_1141) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1122), .B1(n_1123), .B2(n_1125), .C(n_1126), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1121), .B(n_1153), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_1121), .A2(n_1158), .B1(n_1159), .B2(n_1161), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1121), .Y(n_1158) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1122), .Y(n_1130) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI21xp33_ASAP7_75t_L g1167 ( .A1(n_1125), .A2(n_1168), .B(n_1170), .Y(n_1167) );
A2O1A1Ixp33_ASAP7_75t_L g1188 ( .A1(n_1125), .A2(n_1177), .B(n_1189), .C(n_1191), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1129), .C(n_1130), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1128), .B(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1129), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1129), .B(n_1156), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1129), .B(n_1169), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_1132), .A2(n_1135), .B1(n_1136), .B2(n_1137), .C(n_1138), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx2_ASAP7_75t_SL g1186 ( .A(n_1134), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1135), .B(n_1143), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1136), .B(n_1140), .Y(n_1191) );
AOI321xp33_ASAP7_75t_L g1211 ( .A1(n_1137), .A2(n_1158), .A3(n_1207), .B1(n_1212), .B2(n_1216), .C(n_1217), .Y(n_1211) );
A2O1A1Ixp33_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1142), .B(n_1144), .C(n_1146), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1141), .B(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1141), .B(n_1169), .Y(n_1168) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1142), .A2(n_1203), .B(n_1205), .C(n_1211), .Y(n_1202) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1148), .Y(n_1153) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1149), .Y(n_1220) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_1158), .B(n_1194), .C(n_1195), .Y(n_1193) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI21xp5_ASAP7_75t_L g1197 ( .A1(n_1160), .A2(n_1180), .B(n_1186), .Y(n_1197) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
OAI21xp33_ASAP7_75t_L g1183 ( .A1(n_1162), .A2(n_1184), .B(n_1185), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1187), .Y(n_1165) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
OAI211xp5_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1177), .B(n_1179), .C(n_1183), .Y(n_1175) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
NOR3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1192), .C(n_1198), .Y(n_1187) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1194), .Y(n_1213) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1195), .Y(n_1222) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
CKINVDCx14_ASAP7_75t_R g1203 ( .A(n_1204), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .B(n_1209), .Y(n_1205) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1220), .Y(n_1218) );
CKINVDCx20_ASAP7_75t_R g1226 ( .A(n_1227), .Y(n_1226) );
CKINVDCx20_ASAP7_75t_R g1227 ( .A(n_1228), .Y(n_1227) );
INVx4_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
NOR3xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1238), .C(n_1239), .Y(n_1232) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1246), .C(n_1249), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1271), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1254), .B1(n_1256), .B2(n_1257), .Y(n_1252) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_1253), .A2(n_1263), .B1(n_1274), .B2(n_1276), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_1254), .A2(n_1257), .B1(n_1269), .B2(n_1270), .Y(n_1268) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OAI22xp33_ASAP7_75t_L g1282 ( .A1(n_1256), .A2(n_1264), .B1(n_1283), .B2(n_1285), .Y(n_1282) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
OAI33xp33_ASAP7_75t_L g1311 ( .A1(n_1272), .A2(n_1312), .A3(n_1315), .B1(n_1316), .B2(n_1318), .B3(n_1319), .Y(n_1311) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
OAI22xp33_ASAP7_75t_L g1312 ( .A1(n_1276), .A2(n_1300), .B1(n_1306), .B2(n_1313), .Y(n_1312) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1286 ( .A(n_1287), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVxp33_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
NAND3xp33_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1320), .C(n_1328), .Y(n_1296) );
NOR2xp33_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1311), .Y(n_1297) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
endmodule