module fake_netlist_1_12553_n_740 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_740);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_740;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_88), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_84), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_26), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_95), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_29), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_90), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_79), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_27), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_20), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_30), .B(n_18), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_33), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_15), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_100), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_87), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_54), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_85), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_94), .B(n_16), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_42), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_35), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_7), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_19), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_52), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_6), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_28), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_7), .Y(n_131) );
BUFx10_ASAP7_75t_L g132 ( .A(n_2), .Y(n_132) );
INVxp67_ASAP7_75t_SL g133 ( .A(n_73), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_70), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_19), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_68), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_96), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_2), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_49), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_66), .Y(n_140) );
INVx6_ASAP7_75t_L g141 ( .A(n_140), .Y(n_141) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_101), .A2(n_46), .B(n_98), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_128), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_101), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_128), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_119), .B(n_0), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_117), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_102), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_103), .B(n_1), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_102), .B(n_4), .Y(n_150) );
OAI22x1_ASAP7_75t_SL g151 ( .A1(n_127), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_140), .B(n_5), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_104), .B(n_8), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g156 ( .A(n_132), .Y(n_156) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_115), .B(n_50), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_108), .B(n_8), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_131), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_141), .B(n_105), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_149), .A2(n_157), .B1(n_159), .B2(n_148), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_141), .B(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_156), .B(n_120), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_156), .B(n_107), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_141), .B(n_109), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_141), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_141), .B(n_109), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_144), .B(n_121), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_144), .B(n_148), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_159), .B(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_157), .B(n_115), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_154), .A2(n_129), .B1(n_104), .B2(n_135), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_189), .B(n_146), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_184), .A2(n_149), .B1(n_158), .B2(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_189), .B(n_149), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_166), .B(n_158), .C(n_150), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_165), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_174), .B(n_155), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_176), .B(n_149), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_169), .B(n_155), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_179), .B(n_132), .Y(n_201) );
INVxp67_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NOR2x2_ASAP7_75t_L g203 ( .A(n_184), .B(n_151), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_184), .B(n_132), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_183), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g208 ( .A1(n_178), .A2(n_116), .B1(n_106), .B2(n_132), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_169), .B(n_134), .Y(n_210) );
AND2x6_ASAP7_75t_SL g211 ( .A(n_171), .B(n_151), .Y(n_211) );
AND2x6_ASAP7_75t_SL g212 ( .A(n_173), .B(n_147), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_177), .B(n_152), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_181), .B(n_152), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_172), .B(n_137), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_187), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_167), .B(n_152), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_172), .B(n_111), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_163), .B(n_153), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_168), .B(n_126), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_186), .B(n_142), .C(n_153), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_178), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_170), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_185), .B(n_153), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_188), .B(n_110), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_188), .B(n_126), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_190), .B(n_178), .Y(n_230) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_222), .A2(n_182), .B(n_180), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_198), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_199), .A2(n_186), .B(n_142), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_138), .B(n_186), .C(n_147), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_194), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_202), .B(n_178), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_222), .A2(n_186), .B(n_142), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_198), .Y(n_239) );
BUFx6f_ASAP7_75t_SL g240 ( .A(n_194), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_206), .A2(n_142), .B(n_161), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_204), .B(n_160), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_190), .B(n_160), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_197), .B(n_186), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_195), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_196), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_197), .B(n_186), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_192), .B(n_129), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_214), .A2(n_182), .B(n_180), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_223), .B(n_111), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_191), .A2(n_193), .B1(n_192), .B2(n_228), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_193), .B(n_112), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_226), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_230), .B(n_208), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_258), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_240), .B(n_204), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_249), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_233), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_246), .B(n_201), .Y(n_268) );
AND2x6_ASAP7_75t_L g269 ( .A(n_258), .B(n_226), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_214), .B(n_219), .C(n_210), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_217), .B(n_227), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_233), .Y(n_273) );
CKINVDCx11_ASAP7_75t_R g274 ( .A(n_244), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_231), .A2(n_229), .B(n_206), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_255), .A2(n_217), .B(n_213), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_260), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_234), .A2(n_218), .B(n_227), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_246), .B(n_201), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_260), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_SL g281 ( .A1(n_259), .A2(n_225), .B(n_215), .C(n_112), .Y(n_281) );
AOI21x1_ASAP7_75t_L g282 ( .A1(n_238), .A2(n_164), .B(n_162), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g283 ( .A1(n_257), .A2(n_220), .B(n_228), .C(n_135), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_230), .B(n_212), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_240), .Y(n_285) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_282), .A2(n_238), .B(n_231), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_268), .B(n_251), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_270), .A2(n_257), .B(n_253), .Y(n_288) );
OAI21x1_ASAP7_75t_SL g289 ( .A1(n_264), .A2(n_260), .B(n_262), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_284), .A2(n_244), .B1(n_261), .B2(n_251), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_283), .A2(n_272), .B(n_277), .C(n_280), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_272), .B(n_244), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_277), .A2(n_280), .B1(n_264), .B2(n_285), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_269), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_275), .A2(n_243), .B(n_262), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_263), .A2(n_254), .B(n_244), .C(n_261), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_274), .A2(n_228), .B1(n_254), .B2(n_262), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_280), .A2(n_232), .B(n_239), .C(n_247), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g300 ( .A1(n_265), .A2(n_216), .B1(n_220), .B2(n_138), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_282), .A2(n_243), .B(n_122), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_269), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_269), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_275), .A2(n_232), .B(n_241), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_278), .A2(n_122), .B(n_136), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_276), .A2(n_271), .B(n_113), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_293), .B(n_269), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_306), .A2(n_281), .B(n_125), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_297), .A2(n_279), .B1(n_266), .B2(n_256), .C(n_228), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_292), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_303), .B(n_305), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g315 ( .A1(n_290), .A2(n_203), .B(n_103), .C(n_114), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g316 ( .A1(n_300), .A2(n_265), .B(n_266), .C(n_237), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
OR2x6_ASAP7_75t_L g319 ( .A(n_294), .B(n_267), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_287), .B(n_269), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_293), .B(n_285), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_297), .A2(n_114), .B1(n_212), .B2(n_239), .C(n_241), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_293), .B(n_273), .Y(n_325) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_286), .A2(n_113), .B(n_118), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_303), .B(n_269), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_287), .B(n_247), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_290), .A2(n_220), .B1(n_240), .B2(n_233), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_306), .A2(n_118), .B(n_123), .Y(n_330) );
BUFx2_ASAP7_75t_R g331 ( .A(n_306), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_305), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_273), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_295), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_318), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_333), .B(n_306), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g341 ( .A(n_318), .B(n_305), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_319), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_333), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_333), .B(n_306), .Y(n_345) );
AOI31xp33_ASAP7_75t_L g346 ( .A1(n_316), .A2(n_295), .A3(n_300), .B(n_298), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_310), .B(n_288), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_310), .B(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_313), .B(n_288), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_321), .B(n_288), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_321), .B(n_328), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_313), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_332), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_315), .A2(n_298), .B1(n_302), .B2(n_288), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_308), .B(n_307), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_319), .Y(n_363) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_330), .A2(n_301), .B(n_286), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_336), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_308), .B(n_307), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_337), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_337), .B(n_307), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_314), .B(n_307), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_314), .B(n_307), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_312), .A2(n_291), .B1(n_307), .B2(n_220), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_328), .B(n_291), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_319), .B(n_302), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_314), .B(n_296), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_314), .B(n_296), .Y(n_381) );
INVx5_ASAP7_75t_SL g382 ( .A(n_327), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_296), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_327), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_325), .B(n_296), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_335), .B(n_299), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_320), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_334), .B(n_301), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_338), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_376), .B(n_309), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_343), .B(n_327), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_357), .B(n_309), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_369), .B(n_331), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_324), .B1(n_316), .B2(n_326), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_380), .B(n_327), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_343), .B(n_330), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_380), .B(n_326), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_380), .B(n_326), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_343), .B(n_311), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_381), .B(n_326), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_385), .B(n_296), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_355), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_354), .B(n_329), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_344), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_351), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_354), .B(n_311), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_344), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_381), .B(n_123), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_349), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_343), .B(n_311), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_349), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_385), .B(n_9), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_344), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_346), .B(n_267), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_381), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_342), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_361), .B(n_236), .Y(n_424) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_361), .B(n_124), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_358), .B(n_124), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_390), .B(n_10), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_383), .B(n_125), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_342), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_383), .B(n_11), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_347), .B(n_301), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_356), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_356), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_347), .B(n_301), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_347), .B(n_301), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_359), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_360), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_359), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_339), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_371), .B(n_130), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_383), .B(n_374), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_371), .B(n_130), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_339), .Y(n_443) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_363), .B(n_240), .Y(n_444) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_391), .A2(n_136), .B(n_133), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_12), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_367), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_370), .B(n_13), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_370), .B(n_13), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_372), .B(n_14), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_379), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_363), .B(n_220), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_378), .B(n_211), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_378), .B(n_211), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_375), .B(n_170), .Y(n_455) );
INVxp67_ASAP7_75t_R g456 ( .A(n_372), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_384), .B(n_24), .Y(n_457) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_391), .B(n_14), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_374), .B(n_15), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_386), .B(n_16), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_367), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_339), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_372), .B(n_17), .Y(n_463) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_389), .B(n_170), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_362), .B(n_17), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_384), .B(n_65), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_388), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_386), .B(n_18), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_362), .B(n_20), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_360), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_420), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_419), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_457), .B(n_375), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_402), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_428), .B(n_362), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_456), .B(n_384), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_392), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_422), .B(n_340), .Y(n_478) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_444), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_453), .B(n_345), .C(n_340), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_403), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_400), .B(n_340), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_414), .B(n_366), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_465), .B(n_366), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_457), .B(n_341), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_407), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_469), .B(n_366), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_454), .B(n_353), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_464), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_411), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_409), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_406), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_458), .B(n_341), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_415), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_441), .B(n_388), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_409), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_401), .B(n_405), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_430), .B(n_353), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_425), .B(n_389), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_413), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_446), .B(n_345), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_398), .B(n_345), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_462), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_439), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_413), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_417), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_393), .B(n_348), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_395), .B(n_384), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_431), .B(n_352), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_434), .B(n_352), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_448), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_432), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_462), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_435), .B(n_352), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_449), .B(n_368), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g520 ( .A1(n_396), .A2(n_348), .B(n_389), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_437), .B(n_368), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_460), .B(n_379), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_437), .B(n_368), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_396), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_418), .B(n_360), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_436), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_450), .B(n_382), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_438), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_389), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_429), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_463), .B(n_365), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_408), .B(n_365), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_461), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_427), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_439), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_425), .A2(n_389), .B(n_365), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_399), .B(n_364), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_443), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_429), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_416), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_468), .B(n_364), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_443), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_440), .B(n_364), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_399), .B(n_364), .Y(n_546) );
AOI21xp33_ASAP7_75t_SL g547 ( .A1(n_442), .A2(n_21), .B(n_22), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_423), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_445), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_442), .B(n_379), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_440), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_399), .B(n_377), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_423), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_445), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_451), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_440), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_394), .B(n_387), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_459), .B(n_22), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_412), .B(n_382), .Y(n_559) );
AND3x2_ASAP7_75t_L g560 ( .A(n_457), .B(n_387), .C(n_377), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_397), .A2(n_387), .B(n_377), .C(n_373), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_500), .B(n_416), .Y(n_562) );
OAI21xp33_ASAP7_75t_SL g563 ( .A1(n_502), .A2(n_455), .B(n_452), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_495), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g565 ( .A(n_491), .B(n_455), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_524), .B(n_426), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_502), .A2(n_444), .B(n_397), .Y(n_567) );
AOI31xp33_ASAP7_75t_L g568 ( .A1(n_479), .A2(n_421), .A3(n_424), .B(n_416), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_490), .B(n_480), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g570 ( .A(n_491), .B(n_404), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_500), .B(n_394), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_474), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_494), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_490), .B(n_445), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_483), .B(n_404), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_477), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_473), .A2(n_452), .B1(n_421), .B2(n_424), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_514), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_487), .B(n_426), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_512), .B(n_452), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_482), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_493), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_505), .B(n_394), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_512), .B(n_373), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_488), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_473), .A2(n_466), .B1(n_382), .B2(n_373), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_513), .B(n_382), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g589 ( .A(n_506), .B(n_466), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_547), .A2(n_466), .B(n_175), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_492), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_505), .B(n_382), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_558), .A2(n_162), .B(n_164), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_497), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_513), .B(n_517), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_509), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_483), .B(n_510), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_499), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_531), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_555), .B(n_382), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_515), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_517), .B(n_23), .Y(n_603) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_491), .B(n_252), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_478), .B(n_23), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_536), .B(n_161), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_561), .A2(n_175), .B1(n_250), .B2(n_242), .C(n_252), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_478), .B(n_25), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_511), .B(n_31), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g610 ( .A(n_538), .B(n_252), .C(n_250), .D(n_242), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_548), .B(n_32), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_34), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_498), .B(n_36), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_501), .B(n_37), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_553), .B(n_38), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_472), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_533), .B(n_39), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_558), .B(n_250), .C(n_242), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_557), .B(n_40), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_541), .B(n_41), .Y(n_620) );
NAND2xp5_ASAP7_75t_R g621 ( .A(n_539), .B(n_43), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_519), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_526), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_516), .B(n_236), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_245), .B(n_229), .C(n_224), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_529), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_476), .B(n_44), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_518), .B(n_45), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_539), .B(n_47), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_496), .B(n_245), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_535), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_471), .B(n_48), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_534), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_551), .B(n_245), .C(n_229), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_521), .B(n_51), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_534), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_598), .B(n_504), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_562), .B(n_546), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_564), .Y(n_639) );
AOI211xp5_ASAP7_75t_SL g640 ( .A1(n_568), .A2(n_520), .B(n_550), .C(n_556), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_600), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_600), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_563), .A2(n_479), .B(n_550), .C(n_516), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_564), .B(n_542), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_573), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_574), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_579), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_589), .A2(n_569), .A3(n_618), .B1(n_575), .B2(n_571), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_577), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_596), .B(n_540), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_618), .A2(n_522), .B1(n_546), .B2(n_545), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_567), .A2(n_507), .B(n_540), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_570), .B(n_542), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_582), .Y(n_654) );
NAND2xp33_ASAP7_75t_L g655 ( .A(n_589), .B(n_486), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_586), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_591), .A2(n_554), .B(n_549), .C(n_486), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_585), .B(n_532), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_572), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_542), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_565), .A2(n_522), .B(n_527), .C(n_489), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_566), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_594), .A2(n_549), .B1(n_554), .B2(n_485), .C(n_525), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_592), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_566), .A2(n_544), .B(n_537), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_576), .A2(n_559), .B(n_530), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_595), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_578), .A2(n_544), .B(n_537), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_578), .A2(n_530), .B1(n_552), .B2(n_475), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_587), .B(n_552), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_572), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_597), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_602), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_580), .A2(n_552), .B1(n_484), .B2(n_521), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_605), .A2(n_481), .B(n_472), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_587), .B(n_481), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_622), .B(n_523), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_616), .B(n_523), .Y(n_679) );
OAI21xp33_ASAP7_75t_SL g680 ( .A1(n_584), .A2(n_576), .B(n_601), .Y(n_680) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_580), .A2(n_528), .B1(n_508), .B2(n_503), .C1(n_560), .C2(n_58), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_652), .B(n_603), .C(n_629), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_680), .A2(n_581), .B1(n_588), .B2(n_629), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g684 ( .A1(n_643), .A2(n_669), .B1(n_651), .B2(n_662), .C(n_661), .Y(n_684) );
NAND2x1_ASAP7_75t_L g685 ( .A(n_644), .B(n_593), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_638), .B(n_623), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_662), .A2(n_634), .B1(n_608), .B2(n_628), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_640), .A2(n_631), .B1(n_626), .B2(n_624), .C(n_613), .Y(n_688) );
OAI222xp33_ASAP7_75t_L g689 ( .A1(n_647), .A2(n_624), .B1(n_614), .B2(n_609), .C1(n_612), .C2(n_619), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_639), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_639), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_641), .Y(n_692) );
OAI322xp33_ASAP7_75t_L g693 ( .A1(n_675), .A2(n_636), .A3(n_633), .B1(n_606), .B2(n_635), .C1(n_617), .C2(n_599), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_668), .A2(n_604), .B(n_630), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_645), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_679), .B(n_590), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_655), .A2(n_627), .A3(n_599), .B1(n_590), .B2(n_583), .C1(n_634), .C2(n_615), .Y(n_697) );
OAI222xp33_ASAP7_75t_L g698 ( .A1(n_670), .A2(n_625), .B1(n_620), .B2(n_611), .C1(n_607), .C2(n_583), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_642), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_678), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_651), .A2(n_632), .B1(n_528), .B2(n_508), .C(n_503), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_676), .A2(n_621), .B1(n_610), .B2(n_604), .C(n_57), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_665), .B(n_53), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_646), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_666), .A2(n_224), .B1(n_221), .B2(n_206), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_649), .B(n_55), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_684), .A2(n_663), .B1(n_677), .B2(n_681), .C(n_657), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_688), .A2(n_663), .B1(n_657), .B2(n_674), .C(n_664), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_695), .A2(n_648), .B1(n_693), .B2(n_701), .C(n_682), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_698), .A2(n_694), .B(n_697), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_702), .B(n_653), .C(n_650), .D(n_660), .Y(n_711) );
AOI211xp5_ASAP7_75t_L g712 ( .A1(n_698), .A2(n_653), .B(n_674), .C(n_672), .Y(n_712) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_683), .A2(n_673), .B(n_654), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_685), .A2(n_637), .B1(n_658), .B2(n_667), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_700), .B(n_656), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_690), .A2(n_671), .B1(n_659), .B2(n_224), .C(n_221), .Y(n_716) );
OAI321xp33_ASAP7_75t_L g717 ( .A1(n_687), .A2(n_56), .A3(n_59), .B1(n_61), .B2(n_62), .C(n_63), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_689), .B(n_64), .Y(n_718) );
OAI22x1_ASAP7_75t_L g719 ( .A1(n_691), .A2(n_67), .B1(n_69), .B2(n_71), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_708), .B(n_704), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_710), .B(n_703), .C(n_689), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g722 ( .A(n_718), .B(n_706), .C(n_699), .D(n_692), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g723 ( .A1(n_712), .A2(n_687), .B(n_705), .C(n_696), .Y(n_723) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_707), .A2(n_686), .B(n_74), .C(n_76), .Y(n_724) );
NAND3xp33_ASAP7_75t_SL g725 ( .A(n_709), .B(n_72), .C(n_77), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_720), .Y(n_726) );
NAND4xp75_ASAP7_75t_L g727 ( .A(n_725), .B(n_716), .C(n_715), .D(n_711), .Y(n_727) );
NOR4xp25_ASAP7_75t_L g728 ( .A(n_723), .B(n_713), .C(n_717), .D(n_714), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_721), .B(n_719), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_729), .B(n_724), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_729), .Y(n_731) );
OR4x2_ASAP7_75t_L g732 ( .A(n_728), .B(n_722), .C(n_81), .D(n_82), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_731), .Y(n_733) );
AO22x2_ASAP7_75t_L g734 ( .A1(n_730), .A2(n_726), .B1(n_727), .B2(n_86), .Y(n_734) );
AOI22x1_ASAP7_75t_L g735 ( .A1(n_734), .A2(n_732), .B1(n_83), .B2(n_89), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_733), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_735), .A2(n_734), .B1(n_221), .B2(n_92), .Y(n_737) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_737), .B(n_736), .Y(n_738) );
AOI21xp33_ASAP7_75t_SL g739 ( .A1(n_738), .A2(n_80), .B(n_91), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_739), .A2(n_93), .B1(n_97), .B2(n_99), .Y(n_740) );
endmodule