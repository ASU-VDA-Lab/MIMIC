module fake_jpeg_16816_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_32),
.B1(n_19),
.B2(n_21),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_55),
.B1(n_57),
.B2(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_18),
.C(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_0),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_31),
.B1(n_30),
.B2(n_20),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_34),
.B(n_42),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_67),
.B(n_68),
.Y(n_109)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_18),
.CON(n_72),
.SN(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_35),
.B1(n_20),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_81),
.B1(n_43),
.B2(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_30),
.B1(n_31),
.B2(n_2),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_40),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_70),
.B1(n_69),
.B2(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_91),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_0),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_99),
.B(n_87),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_34),
.A3(n_40),
.B1(n_33),
.B2(n_22),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_103),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_100),
.B1(n_94),
.B2(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_103),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_13),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_42),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_115),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_62),
.B1(n_61),
.B2(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_62),
.B1(n_61),
.B2(n_64),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_71),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_33),
.B(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_74),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_64),
.B1(n_74),
.B2(n_77),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_64),
.B1(n_50),
.B2(n_53),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_23),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_54),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_129),
.C(n_113),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_136),
.C(n_138),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_87),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_102),
.B(n_101),
.C(n_88),
.D(n_93),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_150),
.B(n_154),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_108),
.C(n_95),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_41),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_41),
.C(n_104),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_3),
.B(n_5),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_133),
.B(n_132),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_92),
.B(n_0),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_54),
.C(n_96),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_3),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_119),
.B(n_111),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_170),
.B(n_7),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_116),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_126),
.B1(n_118),
.B2(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_169),
.B1(n_178),
.B2(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_145),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_117),
.B1(n_114),
.B2(n_125),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_155),
.B1(n_159),
.B2(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_177),
.B(n_144),
.Y(n_195)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_180),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_7),
.C(n_9),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_148),
.B(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_143),
.B1(n_141),
.B2(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_154),
.B(n_137),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_189),
.B(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_166),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_136),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_162),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_144),
.B(n_9),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_178),
.B(n_165),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_165),
.B(n_176),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_210),
.B(n_196),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_177),
.Y(n_200)
);

XNOR2x2_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_168),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_211),
.B1(n_208),
.B2(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_186),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_215),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_217),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_221),
.C(n_210),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_219),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_191),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_189),
.B(n_188),
.C(n_192),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_182),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_187),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_185),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_192),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_190),
.B(n_197),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_180),
.B1(n_219),
.B2(n_163),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_234),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_172),
.B1(n_171),
.B2(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_225),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_230),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_241),
.B(n_234),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_242),
.A2(n_10),
.B(n_14),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_10),
.A3(n_11),
.B1(n_14),
.B2(n_15),
.C1(n_233),
.C2(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_SL g245 ( 
.A(n_244),
.B(n_237),
.C(n_14),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_10),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_15),
.Y(n_249)
);


endmodule