module fake_jpeg_12204_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_89),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_28),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_19),
.B1(n_38),
.B2(n_36),
.Y(n_125)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_65),
.Y(n_149)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_101),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_9),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_11),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_93),
.B(n_30),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_11),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_105),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_35),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_35),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_46),
.B1(n_47),
.B2(n_21),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_114),
.A2(n_136),
.B1(n_138),
.B2(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_123),
.B(n_132),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_131),
.B1(n_36),
.B2(n_48),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_59),
.A2(n_19),
.B1(n_47),
.B2(n_35),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_25),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_134),
.B(n_137),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_47),
.B1(n_51),
.B2(n_21),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_53),
.B(n_25),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_76),
.A2(n_47),
.B1(n_51),
.B2(n_21),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_82),
.A2(n_104),
.B1(n_100),
.B2(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_25),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_156),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_36),
.B1(n_31),
.B2(n_48),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_96),
.B(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_168),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_71),
.B(n_30),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_174),
.A2(n_228),
.B1(n_70),
.B2(n_74),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_77),
.C(n_64),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_176),
.B(n_198),
.C(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_141),
.A2(n_41),
.B1(n_24),
.B2(n_51),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_180),
.A2(n_193),
.B1(n_203),
.B2(n_215),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_120),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_48),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_197),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_142),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_149),
.A3(n_152),
.B1(n_142),
.B2(n_164),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_196),
.A2(n_52),
.B(n_143),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_34),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_39),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_200),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_136),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_204),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_24),
.B1(n_42),
.B2(n_34),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_206),
.Y(n_262)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_207),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_208),
.B(n_161),
.Y(n_263)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_209),
.B(n_212),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_151),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_161),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_170),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_213),
.B(n_217),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_16),
.C(n_17),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_113),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_127),
.B(n_39),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_218),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_148),
.A2(n_31),
.B1(n_44),
.B2(n_92),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_219),
.A2(n_223),
.B1(n_226),
.B2(n_232),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_224),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_113),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_230),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_166),
.A2(n_44),
.B1(n_94),
.B2(n_91),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_114),
.A2(n_72),
.B1(n_62),
.B2(n_67),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_166),
.B(n_44),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_231),
.C(n_135),
.Y(n_283)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_110),
.B(n_0),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_182),
.A2(n_174),
.B1(n_221),
.B2(n_228),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_239),
.A2(n_251),
.B1(n_278),
.B2(n_216),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_197),
.B(n_176),
.CI(n_227),
.CON(n_243),
.SN(n_243)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_243),
.B(n_266),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_102),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_271),
.C(n_281),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_252),
.Y(n_305)
);

AO22x1_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_84),
.B1(n_116),
.B2(n_110),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_192),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_175),
.A2(n_16),
.B(n_14),
.C(n_13),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_257),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_116),
.Y(n_257)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_210),
.A2(n_97),
.A3(n_105),
.B1(n_143),
.B2(n_140),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_259),
.A2(n_229),
.B(n_218),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_263),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_208),
.B(n_14),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_157),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_268),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_171),
.A2(n_14),
.B(n_12),
.C(n_17),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_229),
.B(n_211),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_171),
.B(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_157),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_201),
.A2(n_140),
.B1(n_135),
.B2(n_130),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_198),
.B(n_52),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_198),
.B(n_130),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_286),
.B(n_0),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_288),
.A2(n_292),
.B1(n_311),
.B2(n_313),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_214),
.B(n_216),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_289),
.A2(n_306),
.B(n_319),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_334),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_212),
.B1(n_232),
.B2(n_218),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_189),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_293),
.B(n_294),
.C(n_312),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_185),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_257),
.A2(n_223),
.B1(n_215),
.B2(n_173),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_300),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_233),
.A2(n_188),
.B1(n_213),
.B2(n_209),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_233),
.A2(n_272),
.B1(n_266),
.B2(n_243),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_243),
.A2(n_178),
.B1(n_179),
.B2(n_191),
.Y(n_300)
);

BUFx24_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_322),
.C(n_324),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_260),
.A2(n_195),
.B(n_206),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_246),
.A2(n_184),
.B(n_217),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_194),
.B1(n_200),
.B2(n_187),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_307),
.A2(n_270),
.B1(n_279),
.B2(n_280),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_199),
.B(n_224),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_250),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_310),
.B(n_315),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_207),
.B1(n_52),
.B2(n_7),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_245),
.B(n_52),
.C(n_1),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_251),
.A2(n_52),
.B1(n_7),
.B2(n_12),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_277),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_52),
.C(n_1),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_321),
.C(n_330),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_6),
.B1(n_15),
.B2(n_13),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_318),
.A2(n_327),
.B1(n_301),
.B2(n_326),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_283),
.A2(n_6),
.B(n_15),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_0),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_240),
.B(n_13),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_268),
.A2(n_17),
.B(n_12),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_323),
.A2(n_327),
.B(n_329),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_236),
.B(n_7),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_252),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_326),
.A2(n_337),
.B1(n_237),
.B2(n_277),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_328),
.B(n_332),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_286),
.A2(n_0),
.B(n_1),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_248),
.B(n_3),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_236),
.B(n_3),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_252),
.A2(n_5),
.B(n_274),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_235),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_235),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_259),
.A2(n_5),
.B1(n_267),
.B2(n_241),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_241),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_298),
.C(n_294),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_253),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_340),
.B(n_365),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_341),
.B(n_351),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_279),
.B(n_270),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_344),
.A2(n_367),
.B(n_360),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_347),
.A2(n_362),
.B1(n_364),
.B2(n_366),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_359),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_301),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_234),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_369),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_337),
.A2(n_237),
.B1(n_280),
.B2(n_253),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_294),
.B(n_284),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_288),
.A2(n_284),
.B1(n_242),
.B2(n_255),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_334),
.A2(n_242),
.B1(n_262),
.B2(n_285),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_367),
.A2(n_363),
.B1(n_381),
.B2(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_265),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_305),
.A2(n_244),
.B1(n_247),
.B2(n_275),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_307),
.B1(n_304),
.B2(n_292),
.Y(n_384)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_301),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_310),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_295),
.A2(n_247),
.B1(n_244),
.B2(n_258),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_296),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_316),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_358),
.B(n_300),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_383),
.A2(n_407),
.B(n_380),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_384),
.A2(n_386),
.B1(n_389),
.B2(n_400),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_297),
.B1(n_325),
.B2(n_336),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_339),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_387),
.B(n_393),
.C(n_406),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_291),
.B1(n_327),
.B2(n_325),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_345),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_391),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_349),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_289),
.B(n_336),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_348),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_409),
.Y(n_430)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_358),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_366),
.A2(n_290),
.B1(n_309),
.B2(n_331),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_308),
.C(n_298),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_356),
.A2(n_331),
.B(n_291),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_340),
.B(n_308),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_417),
.C(n_375),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_371),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_342),
.A2(n_313),
.B1(n_298),
.B2(n_318),
.Y(n_410)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_357),
.A2(n_306),
.B1(n_312),
.B2(n_321),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_415),
.B1(n_418),
.B2(n_419),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_322),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_413),
.B(n_343),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_303),
.B1(n_332),
.B2(n_312),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_317),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_344),
.A2(n_321),
.B1(n_329),
.B2(n_317),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_324),
.B1(n_323),
.B2(n_319),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_360),
.B(n_368),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_420),
.A2(n_435),
.B(n_438),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_378),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_422),
.B(n_431),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_358),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_424),
.B(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_428),
.B(n_432),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_375),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_359),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_396),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_408),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_443),
.C(n_451),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g435 ( 
.A1(n_382),
.A2(n_400),
.B(n_384),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_396),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_436),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_394),
.C(n_401),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_392),
.A2(n_379),
.B(n_346),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_385),
.B(n_369),
.Y(n_442)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_403),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_344),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_382),
.A2(n_370),
.B1(n_364),
.B2(n_373),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_444),
.A2(n_447),
.B1(n_412),
.B2(n_380),
.Y(n_480)
);

OAI22x1_ASAP7_75t_L g445 ( 
.A1(n_404),
.A2(n_380),
.B1(n_346),
.B2(n_352),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_445),
.A2(n_446),
.B(n_448),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_352),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_386),
.A2(n_343),
.B1(n_372),
.B2(n_355),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_449),
.A2(n_402),
.B1(n_395),
.B2(n_397),
.Y(n_454)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_416),
.Y(n_450)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_450),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_338),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_452),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_338),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_415),
.C(n_389),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_454),
.A2(n_473),
.B1(n_354),
.B2(n_258),
.Y(n_505)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_459),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_460),
.B(n_480),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_441),
.A2(n_411),
.B1(n_418),
.B2(n_398),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_461),
.A2(n_261),
.B1(n_256),
.B2(n_238),
.Y(n_506)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_464),
.B1(n_465),
.B2(n_467),
.Y(n_491)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_R g466 ( 
.A(n_440),
.B(n_403),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_479),
.B(n_420),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_427),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_474),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_394),
.C(n_410),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_477),
.C(n_478),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_435),
.A2(n_419),
.B1(n_405),
.B2(n_416),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_443),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_401),
.C(n_397),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_388),
.C(n_412),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_477),
.A2(n_440),
.B(n_469),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_484),
.B(n_496),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_495),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_423),
.Y(n_487)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_429),
.C(n_437),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_424),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_493),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_448),
.B(n_438),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_490),
.A2(n_503),
.B(n_462),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_451),
.C(n_426),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_498),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_455),
.B(n_453),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_463),
.B(n_470),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_445),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_441),
.B1(n_439),
.B2(n_435),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_421),
.C(n_442),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_461),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_501),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_449),
.C(n_423),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_459),
.A2(n_423),
.B(n_377),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_450),
.C(n_354),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_482),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_505),
.A2(n_500),
.B1(n_497),
.B2(n_479),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_487),
.A2(n_481),
.B(n_465),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_508),
.A2(n_509),
.B(n_517),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_502),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_512),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_467),
.Y(n_513)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g515 ( 
.A(n_498),
.B(n_481),
.CI(n_476),
.CON(n_515),
.SN(n_515)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_525),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_501),
.B(n_500),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_505),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_522),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_506),
.Y(n_541)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_521),
.B(n_456),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_538),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_507),
.B(n_456),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_533),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_523),
.B(n_485),
.C(n_488),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_520),
.B(n_485),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_537),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_499),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_524),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_508),
.A2(n_504),
.B(n_495),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_518),
.B(n_509),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_492),
.C(n_489),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_540),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_483),
.C(n_493),
.Y(n_540)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_541),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_542),
.B(n_552),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_483),
.C(n_512),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_545),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_536),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_511),
.C(n_513),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_550),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_511),
.C(n_519),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_486),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_527),
.A2(n_522),
.B(n_514),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_553),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_528),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_555),
.A2(n_560),
.B(n_561),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_546),
.A2(n_526),
.B1(n_531),
.B2(n_514),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_541),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_551),
.A2(n_527),
.B(n_529),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_547),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_562),
.A2(n_563),
.B(n_564),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_548),
.C(n_542),
.Y(n_563)
);

AOI21xp33_ASAP7_75t_L g564 ( 
.A1(n_556),
.A2(n_529),
.B(n_553),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_565),
.B(n_558),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_567),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_565),
.A2(n_554),
.B(n_516),
.Y(n_568)
);

AOI321xp33_ASAP7_75t_L g570 ( 
.A1(n_568),
.A2(n_554),
.A3(n_515),
.B1(n_552),
.B2(n_525),
.C(n_457),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_570),
.B(n_566),
.Y(n_571)
);

BUFx24_ASAP7_75t_SL g572 ( 
.A(n_571),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_569),
.B(n_515),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_482),
.B(n_256),
.Y(n_574)
);


endmodule