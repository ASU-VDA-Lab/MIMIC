module real_aes_8610_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g421 ( .A(n_0), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_1), .A2(n_119), .B(n_131), .C(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g238 ( .A(n_2), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_3), .A2(n_146), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_4), .B(n_142), .Y(n_479) );
AOI21xp33_ASAP7_75t_L g145 ( .A1(n_5), .A2(n_146), .B(n_147), .Y(n_145) );
AND2x6_ASAP7_75t_L g119 ( .A(n_6), .B(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_7), .A2(n_214), .B(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_8), .B(n_41), .Y(n_422) );
INVx1_ASAP7_75t_L g450 ( .A(n_9), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_10), .B(n_152), .Y(n_438) );
INVx1_ASAP7_75t_L g154 ( .A(n_11), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_12), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g220 ( .A(n_14), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_15), .A2(n_155), .B(n_221), .C(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_16), .B(n_142), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_17), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_18), .B(n_165), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_19), .B(n_146), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_20), .B(n_492), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_21), .A2(n_122), .B(n_206), .C(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_22), .B(n_142), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_23), .B(n_152), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_24), .A2(n_218), .B(n_219), .C(n_221), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_25), .B(n_152), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_26), .Y(n_509) );
INVx1_ASAP7_75t_L g499 ( .A(n_27), .Y(n_499) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_28), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_29), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_30), .B(n_152), .Y(n_239) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_31), .A2(n_101), .B1(n_704), .B2(n_713), .C1(n_723), .C2(n_729), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_31), .A2(n_64), .B1(n_718), .B2(n_719), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_31), .Y(n_719) );
INVx1_ASAP7_75t_L g488 ( .A(n_32), .Y(n_488) );
INVx1_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
INVx2_ASAP7_75t_L g124 ( .A(n_34), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_35), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_36), .A2(n_156), .B(n_206), .C(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g489 ( .A(n_37), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_38), .A2(n_119), .B(n_131), .C(n_176), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g475 ( .A(n_39), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_40), .A2(n_131), .B(n_498), .C(n_502), .Y(n_497) );
INVx1_ASAP7_75t_L g128 ( .A(n_42), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_43), .A2(n_151), .B(n_181), .C(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_44), .B(n_152), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_45), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_46), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_47), .A2(n_103), .B1(n_694), .B2(n_697), .C1(n_698), .C2(n_700), .Y(n_102) );
INVx1_ASAP7_75t_L g465 ( .A(n_48), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_49), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_50), .B(n_146), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_51), .A2(n_122), .B1(n_125), .B2(n_131), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_52), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_53), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_54), .A2(n_151), .B(n_153), .C(n_156), .Y(n_150) );
CKINVDCx14_ASAP7_75t_R g447 ( .A(n_55), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_56), .Y(n_195) );
INVx1_ASAP7_75t_L g148 ( .A(n_57), .Y(n_148) );
INVx1_ASAP7_75t_L g120 ( .A(n_58), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_59), .A2(n_77), .B1(n_695), .B2(n_696), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_59), .Y(n_696) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_SL g478 ( .A(n_61), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_62), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_63), .B(n_142), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_64), .Y(n_718) );
INVx1_ASAP7_75t_L g512 ( .A(n_65), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_SL g164 ( .A1(n_66), .A2(n_156), .B(n_165), .C(n_166), .Y(n_164) );
INVxp67_ASAP7_75t_L g167 ( .A(n_67), .Y(n_167) );
INVx1_ASAP7_75t_L g708 ( .A(n_68), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_69), .A2(n_146), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_70), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_71), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_72), .A2(n_146), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g188 ( .A(n_73), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_74), .A2(n_214), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g457 ( .A(n_75), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_76), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_77), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_78), .A2(n_119), .B(n_131), .C(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_79), .A2(n_146), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g460 ( .A(n_80), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_81), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
INVx1_ASAP7_75t_L g436 ( .A(n_83), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_84), .B(n_165), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_85), .A2(n_119), .B(n_131), .C(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g419 ( .A(n_86), .Y(n_419) );
OR2x2_ASAP7_75t_L g693 ( .A(n_86), .B(n_420), .Y(n_693) );
OR2x2_ASAP7_75t_L g712 ( .A(n_86), .B(n_703), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_87), .A2(n_131), .B(n_511), .C(n_514), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_88), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_89), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_90), .A2(n_119), .B(n_131), .C(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_91), .Y(n_210) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_93), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_94), .B(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_95), .B(n_144), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_96), .B(n_144), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_97), .A2(n_146), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g468 ( .A(n_98), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_99), .B(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_416), .B1(n_423), .B2(n_691), .Y(n_103) );
INVx1_ASAP7_75t_L g699 ( .A(n_104), .Y(n_699) );
AND3x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_341), .C(n_390), .Y(n_104) );
NOR3xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_248), .C(n_286), .Y(n_105) );
OAI222xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_169), .B1(n_223), .B2(n_229), .C1(n_243), .C2(n_246), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_140), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_108), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_108), .B(n_291), .Y(n_382) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g259 ( .A(n_109), .B(n_160), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_109), .B(n_141), .Y(n_267) );
AND2x2_ASAP7_75t_L g302 ( .A(n_109), .B(n_279), .Y(n_302) );
OR2x2_ASAP7_75t_L g326 ( .A(n_109), .B(n_141), .Y(n_326) );
OR2x2_ASAP7_75t_L g334 ( .A(n_109), .B(n_233), .Y(n_334) );
AND2x2_ASAP7_75t_L g337 ( .A(n_109), .B(n_160), .Y(n_337) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g231 ( .A(n_110), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g245 ( .A(n_110), .B(n_160), .Y(n_245) );
AND2x2_ASAP7_75t_L g295 ( .A(n_110), .B(n_233), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_110), .B(n_141), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_110), .B(n_394), .Y(n_415) );
AO21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_117), .B(n_138), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_111), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g183 ( .A(n_111), .Y(n_183) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_111), .A2(n_234), .B(n_241), .Y(n_233) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_113), .B(n_114), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OAI22xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B1(n_134), .B2(n_135), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_118), .A2(n_148), .B(n_149), .C(n_150), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_118), .A2(n_149), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_118), .A2(n_149), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_118), .A2(n_149), .B(n_447), .C(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_118), .A2(n_149), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_118), .A2(n_149), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_118), .A2(n_149), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_118), .A2(n_149), .B(n_485), .C(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g514 ( .A(n_118), .Y(n_514) );
INVx4_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_119), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g146 ( .A(n_119), .B(n_136), .Y(n_146) );
BUFx3_ASAP7_75t_L g502 ( .A(n_119), .Y(n_502) );
INVx2_ASAP7_75t_L g240 ( .A(n_122), .Y(n_240) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_125) );
INVx2_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
INVx4_ASAP7_75t_L g218 ( .A(n_126), .Y(n_218) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
AND2x2_ASAP7_75t_L g136 ( .A(n_127), .B(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
INVx2_ASAP7_75t_L g437 ( .A(n_129), .Y(n_437) );
INVx5_ASAP7_75t_L g149 ( .A(n_131), .Y(n_149) );
AND2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
BUFx3_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_135), .A2(n_188), .B(n_189), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_135), .A2(n_235), .B(n_236), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_135), .A2(n_433), .B(n_434), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_135), .A2(n_159), .B(n_496), .C(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_135), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g490 ( .A(n_137), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_140), .A2(n_334), .B(n_335), .C(n_338), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_140), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_140), .B(n_278), .Y(n_400) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_160), .Y(n_140) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_141), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g258 ( .A(n_141), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_141), .B(n_279), .Y(n_285) );
INVx1_ASAP7_75t_SL g293 ( .A(n_141), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_141), .B(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g394 ( .A(n_141), .Y(n_394) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_158), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g184 ( .A(n_143), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_143), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_143), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_143), .A2(n_508), .B(n_515), .Y(n_507) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_144), .A2(n_161), .B(n_168), .Y(n_160) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_144), .Y(n_454) );
BUFx2_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_155), .B(n_167), .Y(n_166) );
INVx5_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_155), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_213), .B(n_222), .Y(n_212) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_159), .A2(n_445), .B(n_451), .Y(n_444) );
BUFx2_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g292 ( .A(n_160), .Y(n_292) );
INVx3_ASAP7_75t_L g317 ( .A(n_160), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_169), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_197), .Y(n_169) );
INVx1_ASAP7_75t_L g313 ( .A(n_170), .Y(n_313) );
OAI32xp33_ASAP7_75t_L g319 ( .A1(n_170), .A2(n_258), .A3(n_320), .B1(n_321), .B2(n_322), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_170), .A2(n_324), .B1(n_327), .B2(n_332), .Y(n_323) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g261 ( .A(n_171), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g339 ( .A(n_171), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g409 ( .A(n_171), .B(n_355), .Y(n_409) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_186), .Y(n_171) );
AND2x2_ASAP7_75t_L g224 ( .A(n_172), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
INVx1_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
OR2x2_ASAP7_75t_L g281 ( .A(n_172), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_172), .B(n_262), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_172), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_172), .B(n_227), .Y(n_309) );
INVx3_ASAP7_75t_L g331 ( .A(n_172), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_172), .B(n_228), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_172), .B(n_321), .Y(n_404) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_184), .Y(n_172) );
AOI21xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_183), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_180), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_178), .A2(n_238), .B(n_239), .C(n_240), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_178), .A2(n_218), .B1(n_488), .B2(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_178), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_180), .A2(n_191), .B(n_192), .Y(n_190) );
O2A1O1Ixp5_ASAP7_75t_L g435 ( .A1(n_180), .A2(n_436), .B(n_437), .C(n_438), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_180), .A2(n_437), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
INVx1_ASAP7_75t_L g193 ( .A(n_183), .Y(n_193) );
INVx2_ASAP7_75t_L g228 ( .A(n_186), .Y(n_228) );
AND2x2_ASAP7_75t_L g360 ( .A(n_186), .B(n_198), .Y(n_360) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_186) );
INVx1_ASAP7_75t_L g482 ( .A(n_193), .Y(n_482) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_193), .A2(n_535), .B(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_196), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_196), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_196), .A2(n_432), .B(n_439), .Y(n_431) );
INVx2_ASAP7_75t_L g402 ( .A(n_197), .Y(n_402) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_211), .Y(n_197) );
INVx1_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
AND2x2_ASAP7_75t_L g274 ( .A(n_198), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_198), .B(n_228), .Y(n_282) );
AND2x2_ASAP7_75t_L g340 ( .A(n_198), .B(n_263), .Y(n_340) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g226 ( .A(n_199), .Y(n_226) );
AND2x2_ASAP7_75t_L g253 ( .A(n_199), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_199), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_199), .B(n_228), .Y(n_328) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_209), .Y(n_199) );
INVx1_ASAP7_75t_L g492 ( .A(n_200), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_200), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_208), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_206), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_211), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_211), .B(n_228), .Y(n_321) );
AND2x2_ASAP7_75t_L g330 ( .A(n_211), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g355 ( .A(n_211), .Y(n_355) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g227 ( .A(n_212), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_218), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_218), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_218), .B(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_223), .A2(n_233), .B1(n_392), .B2(n_395), .Y(n_391) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_225), .A2(n_336), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_226), .B(n_331), .Y(n_348) );
INVx1_ASAP7_75t_L g373 ( .A(n_226), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_227), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g300 ( .A(n_227), .B(n_253), .Y(n_300) );
INVx2_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_229), .A2(n_381), .B1(n_398), .B2(n_401), .C(n_403), .Y(n_397) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_230), .B(n_279), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_231), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_268), .Y(n_322) );
INVx3_ASAP7_75t_SL g363 ( .A(n_231), .Y(n_363) );
AND2x2_ASAP7_75t_L g307 ( .A(n_232), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_232), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_232), .B(n_245), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_232), .B(n_291), .Y(n_377) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
OAI322xp33_ASAP7_75t_L g374 ( .A1(n_233), .A2(n_305), .A3(n_327), .B1(n_375), .B2(n_377), .C1(n_378), .C2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_244), .A2(n_247), .B(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_SL g324 ( .A(n_245), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g346 ( .A(n_245), .B(n_258), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_245), .B(n_285), .Y(n_361) );
INVxp67_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_247), .A2(n_319), .B(n_323), .C(n_333), .Y(n_318) );
OAI221xp5_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_257), .B1(n_260), .B2(n_264), .C(n_269), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g272 ( .A(n_256), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g389 ( .A(n_256), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_257), .A2(n_406), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_405) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_258), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g305 ( .A(n_258), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_258), .B(n_336), .Y(n_343) );
AND2x2_ASAP7_75t_L g385 ( .A(n_258), .B(n_363), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_259), .B(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_259), .A2(n_271), .B1(n_381), .B2(n_382), .Y(n_380) );
OR2x2_ASAP7_75t_L g411 ( .A(n_259), .B(n_279), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g388 ( .A(n_262), .Y(n_388) );
AND2x2_ASAP7_75t_L g413 ( .A(n_262), .B(n_356), .Y(n_413) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g277 ( .A(n_267), .B(n_278), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_276), .B1(n_280), .B2(n_283), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_272), .B(n_312), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g303 ( .A1(n_274), .A2(n_304), .A3(n_306), .B1(n_307), .B2(n_309), .C1(n_310), .C2(n_314), .Y(n_303) );
INVxp67_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_277), .A2(n_282), .B1(n_299), .B2(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_278), .B(n_291), .Y(n_378) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_279), .B(n_317), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_279), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g375 ( .A(n_281), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_303), .C(n_318), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_294), .B2(n_296), .C(n_298), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_290), .B(n_295), .Y(n_294) );
INVx3_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_295), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_297), .Y(n_376) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_302), .B(n_316), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_305), .B(n_363), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_306), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g381 ( .A(n_309), .Y(n_381) );
AND2x2_ASAP7_75t_L g396 ( .A(n_309), .B(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_320), .A2(n_391), .B(n_397), .C(n_405), .Y(n_390) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_360), .Y(n_359) );
NAND2x1_ASAP7_75t_SL g401 ( .A(n_331), .B(n_402), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g371 ( .A(n_334), .Y(n_371) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g366 ( .A(n_340), .Y(n_366) );
AND2x2_ASAP7_75t_L g370 ( .A(n_340), .B(n_356), .Y(n_370) );
NOR5xp2_ASAP7_75t_L g341 ( .A(n_342), .B(n_357), .C(n_374), .D(n_380), .E(n_383), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_345), .B2(n_347), .C(n_349), .Y(n_342) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_346), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g372 ( .A(n_356), .B(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B1(n_362), .B2(n_364), .C(n_367), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_371), .B2(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AOI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_388), .C(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g698 ( .A1(n_416), .A2(n_424), .B1(n_693), .B2(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
NOR2x2_ASAP7_75t_L g702 ( .A(n_419), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_420), .Y(n_703) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_423), .A2(n_424), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_646), .Y(n_424) );
NAND5xp2_ASAP7_75t_L g425 ( .A(n_426), .B(n_558), .C(n_596), .D(n_617), .E(n_634), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_530), .C(n_551), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_470), .B1(n_493), .B2(n_517), .C(n_521), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_441), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_430), .B(n_519), .Y(n_538) );
OR2x2_ASAP7_75t_L g565 ( .A(n_430), .B(n_453), .Y(n_565) );
AND2x2_ASAP7_75t_L g579 ( .A(n_430), .B(n_453), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_430), .B(n_444), .Y(n_593) );
AND2x2_ASAP7_75t_L g631 ( .A(n_430), .B(n_595), .Y(n_631) );
AND2x2_ASAP7_75t_L g660 ( .A(n_430), .B(n_570), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_430), .B(n_542), .Y(n_677) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g557 ( .A(n_431), .B(n_452), .Y(n_557) );
BUFx3_ASAP7_75t_L g582 ( .A(n_431), .Y(n_582) );
AND2x2_ASAP7_75t_L g611 ( .A(n_431), .B(n_453), .Y(n_611) );
AND3x2_ASAP7_75t_L g624 ( .A(n_431), .B(n_625), .C(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g547 ( .A(n_441), .Y(n_547) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .Y(n_441) );
AOI32xp33_ASAP7_75t_L g602 ( .A1(n_442), .A2(n_554), .A3(n_603), .B1(n_606), .B2(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g529 ( .A(n_443), .B(n_452), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_443), .B(n_557), .Y(n_600) );
AND2x2_ASAP7_75t_L g607 ( .A(n_443), .B(n_579), .Y(n_607) );
OR2x2_ASAP7_75t_L g613 ( .A(n_443), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_443), .B(n_568), .Y(n_638) );
OR2x2_ASAP7_75t_L g656 ( .A(n_443), .B(n_481), .Y(n_656) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g520 ( .A(n_444), .B(n_462), .Y(n_520) );
INVx2_ASAP7_75t_L g542 ( .A(n_444), .Y(n_542) );
OR2x2_ASAP7_75t_L g564 ( .A(n_444), .B(n_462), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_444), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_444), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_444), .B(n_519), .Y(n_625) );
INVx1_ASAP7_75t_SL g676 ( .A(n_452), .Y(n_676) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
INVx1_ASAP7_75t_SL g519 ( .A(n_453), .Y(n_519) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_453), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_453), .B(n_605), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_453), .B(n_542), .C(n_660), .Y(n_671) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_461), .Y(n_453) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_454), .A2(n_463), .B(n_469), .Y(n_462) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_454), .A2(n_473), .B(n_479), .Y(n_472) );
INVx2_ASAP7_75t_L g570 ( .A(n_462), .Y(n_570) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_462), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
INVx1_ASAP7_75t_L g606 ( .A(n_471), .Y(n_606) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g524 ( .A(n_472), .B(n_506), .Y(n_524) );
INVx2_ASAP7_75t_L g541 ( .A(n_472), .Y(n_541) );
AND2x2_ASAP7_75t_L g546 ( .A(n_472), .B(n_507), .Y(n_546) );
AND2x2_ASAP7_75t_L g561 ( .A(n_472), .B(n_494), .Y(n_561) );
AND2x2_ASAP7_75t_L g573 ( .A(n_472), .B(n_545), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_480), .B(n_589), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_480), .B(n_546), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_480), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_480), .B(n_540), .Y(n_668) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g505 ( .A(n_481), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_481), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g550 ( .A(n_481), .B(n_494), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_481), .B(n_506), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_481), .B(n_616), .Y(n_615) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_491), .Y(n_481) );
INVx1_ASAP7_75t_L g535 ( .A(n_483), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx2_ASAP7_75t_L g501 ( .A(n_490), .Y(n_501) );
INVx1_ASAP7_75t_L g536 ( .A(n_491), .Y(n_536) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_494), .B(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g540 ( .A(n_494), .B(n_541), .Y(n_540) );
INVx3_ASAP7_75t_SL g545 ( .A(n_494), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_494), .B(n_532), .Y(n_598) );
OR2x2_ASAP7_75t_L g608 ( .A(n_494), .B(n_534), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_494), .B(n_576), .Y(n_636) );
OR2x2_ASAP7_75t_L g666 ( .A(n_494), .B(n_506), .Y(n_666) );
AND2x2_ASAP7_75t_L g670 ( .A(n_494), .B(n_507), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_494), .B(n_546), .Y(n_683) );
AND2x2_ASAP7_75t_L g690 ( .A(n_494), .B(n_572), .Y(n_690) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx1_ASAP7_75t_SL g633 ( .A(n_505), .Y(n_633) );
AND2x2_ASAP7_75t_L g572 ( .A(n_506), .B(n_534), .Y(n_572) );
AND2x2_ASAP7_75t_L g586 ( .A(n_506), .B(n_541), .Y(n_586) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_545), .Y(n_589) );
INVx1_ASAP7_75t_L g616 ( .A(n_506), .Y(n_616) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_518), .A2(n_564), .B(n_688), .C(n_689), .Y(n_687) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g594 ( .A(n_519), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_520), .B(n_537), .Y(n_552) );
AND2x2_ASAP7_75t_L g578 ( .A(n_520), .B(n_579), .Y(n_578) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_525), .B(n_529), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_523), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g549 ( .A(n_524), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_524), .B(n_545), .Y(n_590) );
AND2x2_ASAP7_75t_L g681 ( .A(n_524), .B(n_532), .Y(n_681) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g554 ( .A(n_528), .B(n_541), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_528), .B(n_539), .Y(n_555) );
OAI322xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_538), .A3(n_539), .B1(n_542), .B2(n_543), .C1(n_547), .C2(n_548), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
AND2x2_ASAP7_75t_L g642 ( .A(n_532), .B(n_554), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_532), .B(n_606), .Y(n_688) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g585 ( .A(n_534), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_564), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_539), .B(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_540), .B(n_572), .Y(n_629) );
AND2x2_ASAP7_75t_L g575 ( .A(n_541), .B(n_545), .Y(n_575) );
AND2x2_ASAP7_75t_L g583 ( .A(n_542), .B(n_584), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_542), .A2(n_621), .B(n_681), .C(n_682), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_543), .A2(n_556), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_545), .B(n_572), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_545), .B(n_586), .Y(n_618) );
AND2x2_ASAP7_75t_L g652 ( .A(n_545), .B(n_554), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_546), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g662 ( .A(n_546), .Y(n_662) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_550), .A2(n_578), .B1(n_580), .B2(n_585), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_552), .A2(n_588), .B1(n_590), .B2(n_591), .Y(n_587) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_557), .A2(n_659), .B1(n_661), .B2(n_663), .C(n_667), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_566), .C(n_587), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OR2x2_ASAP7_75t_L g628 ( .A(n_564), .B(n_581), .Y(n_628) );
INVx1_ASAP7_75t_L g679 ( .A(n_564), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_565), .A2(n_567), .B1(n_571), .B2(n_574), .C(n_577), .Y(n_566) );
INVx2_ASAP7_75t_SL g621 ( .A(n_565), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g686 ( .A(n_568), .Y(n_686) );
AND2x2_ASAP7_75t_L g610 ( .A(n_569), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g595 ( .A(n_570), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g657 ( .A(n_573), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_581), .B(n_683), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g626 ( .A(n_584), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_585), .A2(n_597), .B(n_599), .C(n_601), .Y(n_596) );
INVx1_ASAP7_75t_L g674 ( .A(n_588), .Y(n_674) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_592), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g605 ( .A(n_595), .Y(n_605) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI222xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_608), .B1(n_609), .B2(n_612), .C1(n_613), .C2(n_615), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g641 ( .A(n_605), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_608), .B(n_662), .Y(n_661) );
NAND2xp33_ASAP7_75t_SL g639 ( .A(n_609), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g614 ( .A(n_611), .Y(n_614) );
AND2x2_ASAP7_75t_L g678 ( .A(n_611), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g644 ( .A(n_614), .B(n_641), .Y(n_644) );
INVx1_ASAP7_75t_L g673 ( .A(n_615), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B(n_622), .C(n_627), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_621), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AOI322xp5_ASAP7_75t_L g672 ( .A1(n_624), .A2(n_652), .A3(n_657), .B1(n_673), .B2(n_674), .C1(n_675), .C2(n_678), .Y(n_672) );
AND2x2_ASAP7_75t_L g659 ( .A(n_625), .B(n_660), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_630), .B2(n_632), .Y(n_627) );
INVxp33_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_639), .B2(n_642), .C(n_643), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_647), .B(n_658), .C(n_672), .D(n_680), .E(n_684), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_652), .B(n_653), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_660), .A2(n_685), .B(n_686), .C(n_687), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g667 ( .A1(n_662), .A2(n_668), .A3(n_669), .B(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g685 ( .A(n_683), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
CKINVDCx14_ASAP7_75t_R g697 ( .A(n_694), .Y(n_697) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx3_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
NOR2xp33_ASAP7_75t_SL g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g728 ( .A(n_707), .Y(n_728) );
INVx1_ASAP7_75t_L g727 ( .A(n_709), .Y(n_727) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_709), .A2(n_728), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g714 ( .A(n_712), .Y(n_714) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_712), .Y(n_722) );
BUFx2_ASAP7_75t_L g731 ( .A(n_712), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_720), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
endmodule