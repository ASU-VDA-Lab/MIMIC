module real_aes_18016_n_13 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_13);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_13;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_19;
wire n_25;
wire n_30;
wire n_14;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
AOI322xp5_ASAP7_75t_R g13 ( .A1(n_0), .A2(n_4), .A3(n_8), .B1(n_14), .B2(n_16), .C1(n_23), .C2(n_27), .Y(n_13) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_1), .B(n_7), .C(n_19), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_2), .B(n_15), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_2), .B(n_5), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_2), .Y(n_30) );
NOR5xp2_ASAP7_75t_SL g16 ( .A(n_3), .B(n_10), .C(n_17), .D(n_21), .E(n_22), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_5), .B(n_30), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_6), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_9), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_11), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_12), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_16), .Y(n_26) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_20), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_24), .B(n_26), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_25), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_26), .B(n_28), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_29), .Y(n_28) );
endmodule