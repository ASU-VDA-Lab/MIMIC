module fake_jpeg_24535_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_25),
.Y(n_49)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_48),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_26),
.B1(n_14),
.B2(n_60),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_35),
.B(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_18),
.B1(n_16),
.B2(n_27),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_14),
.B1(n_18),
.B2(n_16),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_41),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_67),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_51),
.B1(n_62),
.B2(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_72),
.B1(n_62),
.B2(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_39),
.B1(n_45),
.B2(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_45),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_78),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_23),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_67),
.B1(n_75),
.B2(n_77),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_68),
.B(n_66),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_0),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_43),
.B(n_2),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_80),
.B(n_74),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_106),
.B1(n_89),
.B2(n_87),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_73),
.C(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_102),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_86),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_114),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_85),
.C(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_115),
.C(n_5),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_86),
.B1(n_82),
.B2(n_93),
.Y(n_112)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_96),
.A3(n_103),
.B1(n_105),
.B2(n_100),
.C(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_92),
.C(n_24),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_112),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_123),
.B(n_114),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_2),
.CI(n_3),
.CON(n_119),
.SN(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_115),
.C(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_5),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.C(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_109),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_120),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_117),
.B(n_119),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_131),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_10),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_129),
.C(n_11),
.Y(n_138)
);

AOI321xp33_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_6),
.A3(n_12),
.B1(n_136),
.B2(n_92),
.C(n_126),
.Y(n_139)
);


endmodule