module fake_aes_2897_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx4_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVxp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_10), .B(n_6), .Y(n_16) );
BUFx2_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_2), .B(n_9), .Y(n_18) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_17), .B(n_0), .C(n_1), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_13), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_19), .B1(n_13), .B2(n_15), .C(n_18), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_25), .B(n_16), .C(n_2), .Y(n_26) );
OR4x1_ASAP7_75t_L g27 ( .A(n_26), .B(n_1), .C(n_3), .D(n_4), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_16), .B1(n_4), .B2(n_3), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_7), .B(n_12), .Y(n_29) );
endmodule