module fake_jpeg_31340_n_127 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_127);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_25),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_14),
.B1(n_18),
.B2(n_24),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_14),
.B1(n_18),
.B2(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_35),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_43),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_31),
.B1(n_35),
.B2(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_79),
.B1(n_32),
.B2(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_15),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_28),
.B(n_47),
.C(n_32),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_55),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_36),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_93),
.B(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_79),
.B(n_70),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_79),
.B(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_106),
.B1(n_109),
.B2(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_74),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_73),
.A3(n_52),
.B1(n_53),
.B2(n_78),
.C1(n_6),
.C2(n_0),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_100),
.C(n_98),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_114),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_112),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_117),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_102),
.B1(n_16),
.B2(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_48),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

AOI31xp33_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_115),
.A3(n_6),
.B(n_7),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_1),
.B(n_29),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_122),
.B(n_119),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_1),
.Y(n_127)
);


endmodule