module fake_jpeg_793_n_39 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_22),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_15),
.C(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_15),
.B1(n_16),
.B2(n_24),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_26),
.B1(n_16),
.B2(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_17),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_0),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.A3(n_17),
.B1(n_7),
.B2(n_6),
.C1(n_3),
.C2(n_0),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_4),
.B(n_5),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_4),
.Y(n_39)
);


endmodule