module fake_jpeg_21008_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

OAI32xp33_ASAP7_75t_L g12 ( 
.A1(n_10),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_8),
.B1(n_7),
.B2(n_9),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.C(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_11),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_6),
.B(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_8),
.B1(n_7),
.B2(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_8),
.B1(n_9),
.B2(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_12),
.Y(n_30)
);

NOR2xp67_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_27),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B(n_2),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_24),
.C(n_4),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g35 ( 
.A(n_34),
.Y(n_35)
);


endmodule