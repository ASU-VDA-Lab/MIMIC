module fake_aes_3393_n_48 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_30;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_7), .B(n_1), .Y(n_16) );
AND2x6_ASAP7_75t_L g17 ( .A(n_8), .B(n_9), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_3), .B(n_10), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_4), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_5), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_15), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_22), .B(n_0), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_20), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_17), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_19), .Y(n_29) );
BUFx4f_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
OR2x6_ASAP7_75t_L g31 ( .A(n_29), .B(n_16), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_27), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_27), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_31), .B(n_26), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_33), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_35), .B(n_32), .Y(n_37) );
INVx1_ASAP7_75t_SL g38 ( .A(n_34), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
NAND4xp25_ASAP7_75t_L g40 ( .A(n_36), .B(n_23), .C(n_21), .D(n_18), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
OAI21xp33_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_38), .B(n_28), .Y(n_42) );
INVx3_ASAP7_75t_L g43 ( .A(n_41), .Y(n_43) );
NOR4xp75_ASAP7_75t_L g44 ( .A(n_42), .B(n_6), .C(n_13), .D(n_24), .Y(n_44) );
BUFx6f_ASAP7_75t_L g45 ( .A(n_43), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_43), .Y(n_46) );
XOR2xp5_ASAP7_75t_L g47 ( .A(n_45), .B(n_44), .Y(n_47) );
AOI22xp5_ASAP7_75t_SL g48 ( .A1(n_47), .A2(n_45), .B1(n_46), .B2(n_44), .Y(n_48) );
endmodule