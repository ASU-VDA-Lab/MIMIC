module fake_jpeg_20690_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_37),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_70),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_64),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_22),
.B1(n_13),
.B2(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_13),
.B(n_32),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_22),
.B1(n_14),
.B2(n_13),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_22),
.B1(n_47),
.B2(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_82),
.B1(n_55),
.B2(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_47),
.B1(n_20),
.B2(n_22),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_95),
.B1(n_52),
.B2(n_20),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_83),
.Y(n_113)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_70),
.Y(n_98)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_63),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_56),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_103),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_19),
.B(n_90),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_90),
.B1(n_76),
.B2(n_77),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_91),
.B1(n_92),
.B2(n_14),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_65),
.C(n_66),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_115),
.C(n_71),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_69),
.B1(n_68),
.B2(n_63),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_82),
.B1(n_79),
.B2(n_90),
.Y(n_121)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_85),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_64),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_14),
.B1(n_20),
.B2(n_61),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_86),
.B1(n_88),
.B2(n_94),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_92),
.B1(n_111),
.B2(n_85),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_89),
.B(n_86),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_127),
.B(n_129),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_88),
.C(n_80),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_131),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_135),
.B(n_15),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_76),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_99),
.B(n_85),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_141),
.B1(n_142),
.B2(n_20),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_84),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_76),
.C(n_71),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_140),
.C(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_26),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_71),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_115),
.C(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_92),
.B1(n_14),
.B2(n_24),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_106),
.C(n_112),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_154),
.Y(n_171)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_101),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_101),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_111),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_165),
.B1(n_137),
.B2(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_23),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_25),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_61),
.C(n_29),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_131),
.C(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_21),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_191),
.C(n_146),
.Y(n_203)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_177),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_176),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_193),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_161),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_137),
.B(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_158),
.B1(n_167),
.B2(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_142),
.Y(n_191)
);

INVxp33_ASAP7_75t_SL g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_189),
.B(n_175),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_201),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_169),
.B(n_161),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_199),
.B(n_204),
.C(n_173),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_183),
.B(n_174),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_173),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_177),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_162),
.B1(n_153),
.B2(n_149),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_207),
.B1(n_180),
.B2(n_178),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_129),
.B1(n_127),
.B2(n_21),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_19),
.Y(n_208)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_0),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_176),
.C(n_191),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_221),
.C(n_228),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_220),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_198),
.B(n_204),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_171),
.B1(n_21),
.B2(n_17),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_196),
.B1(n_197),
.B2(n_18),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_16),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_207),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_230),
.B1(n_227),
.B2(n_194),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_17),
.C(n_18),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_243),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_198),
.B1(n_204),
.B2(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_241),
.B1(n_27),
.B2(n_18),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_244),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_220),
.C(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_232),
.C(n_236),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_199),
.B(n_17),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_219),
.B1(n_223),
.B2(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_219),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_232),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_251),
.B1(n_0),
.B2(n_2),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_27),
.B1(n_10),
.B2(n_16),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_10),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_265),
.C(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_16),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_252),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_263),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_15),
.C(n_4),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_245),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_3),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_254),
.B1(n_246),
.B2(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_272),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_271),
.Y(n_278)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_3),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_259),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_281),
.B(n_276),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_282),
.B(n_278),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_275),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_278),
.B(n_273),
.C(n_6),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_6),
.B(n_276),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_6),
.Y(n_289)
);


endmodule