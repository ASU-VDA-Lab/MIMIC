module real_aes_978_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_577;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_528;
wire n_578;
wire n_495;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_559;
wire n_636;
wire n_872;
wire n_466;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_817;
wire n_443;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_737;
wire n_1017;
wire n_936;
wire n_610;
wire n_581;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_967;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_0), .A2(n_45), .B1(n_698), .B2(n_764), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_1), .A2(n_230), .B1(n_547), .B2(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_2), .A2(n_313), .B1(n_492), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_3), .A2(n_79), .B1(n_448), .B2(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_4), .A2(n_139), .B1(n_741), .B2(n_742), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_5), .A2(n_18), .B1(n_575), .B2(n_710), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_6), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_7), .A2(n_250), .B1(n_458), .B2(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_8), .A2(n_86), .B1(n_436), .B2(n_482), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_9), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_10), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_11), .A2(n_351), .B1(n_484), .B2(n_597), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_12), .A2(n_77), .B1(n_709), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_13), .A2(n_25), .B1(n_507), .B2(n_510), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_14), .A2(n_213), .B1(n_507), .B2(n_552), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_15), .A2(n_205), .B1(n_611), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_16), .A2(n_252), .B1(n_512), .B2(n_515), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_17), .A2(n_259), .B1(n_675), .B2(n_784), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_19), .A2(n_324), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_20), .A2(n_305), .B1(n_504), .B2(n_861), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_21), .A2(n_93), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_22), .A2(n_195), .B1(n_458), .B2(n_522), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_23), .A2(n_337), .B1(n_408), .B2(n_424), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_24), .A2(n_201), .B1(n_764), .B2(n_863), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_26), .A2(n_256), .B1(n_408), .B2(n_424), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_27), .B(n_960), .Y(n_959) );
AOI22x1_ASAP7_75t_L g900 ( .A1(n_28), .A2(n_901), .B1(n_902), .B2(n_916), .Y(n_900) );
INVx1_ASAP7_75t_L g916 ( .A(n_28), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_29), .A2(n_298), .B1(n_530), .B2(n_532), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_30), .A2(n_257), .B1(n_486), .B2(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_31), .B(n_943), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_32), .A2(n_478), .B1(n_523), .B2(n_524), .Y(n_477) );
INVx1_ASAP7_75t_L g523 ( .A(n_32), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_33), .A2(n_285), .B1(n_510), .B2(n_519), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_34), .A2(n_151), .B1(n_481), .B2(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g419 ( .A(n_35), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_35), .B(n_54), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_36), .A2(n_39), .B1(n_458), .B2(n_465), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_37), .A2(n_128), .B1(n_781), .B2(n_844), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_38), .A2(n_272), .B1(n_542), .B2(n_996), .Y(n_995) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_40), .A2(n_316), .B1(n_354), .B2(n_428), .C1(n_680), .C2(n_682), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_41), .B(n_569), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_42), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_43), .A2(n_350), .B1(n_549), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_44), .A2(n_94), .B1(n_636), .B2(n_670), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_46), .A2(n_140), .B1(n_448), .B2(n_675), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_47), .A2(n_239), .B1(n_611), .B2(n_639), .Y(n_638) );
XNOR2x1_ASAP7_75t_SL g564 ( .A(n_48), .B(n_565), .Y(n_564) );
AOI22xp5_ASAP7_75t_SL g614 ( .A1(n_48), .A2(n_565), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_48), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_49), .A2(n_265), .B1(n_531), .B2(n_710), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_50), .A2(n_119), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_51), .A2(n_114), .B1(n_641), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_52), .A2(n_254), .B1(n_580), .B2(n_1020), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_53), .A2(n_383), .B1(n_391), .B2(n_975), .C(n_985), .Y(n_382) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_54), .A2(n_359), .B1(n_411), .B2(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_55), .A2(n_271), .B1(n_490), .B2(n_492), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_56), .A2(n_120), .B1(n_610), .B2(n_611), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_57), .A2(n_200), .B1(n_639), .B2(n_865), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_58), .A2(n_210), .B1(n_436), .B2(n_735), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_59), .A2(n_106), .B1(n_471), .B2(n_472), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_60), .A2(n_279), .B1(n_501), .B2(n_607), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_61), .A2(n_125), .B1(n_555), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_62), .A2(n_284), .B1(n_592), .B2(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g420 ( .A(n_63), .Y(n_420) );
AO222x2_ASAP7_75t_SL g921 ( .A1(n_64), .A2(n_214), .B1(n_292), .B2(n_408), .C1(n_424), .C2(n_429), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_65), .A2(n_352), .B1(n_714), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_66), .A2(n_215), .B1(n_482), .B2(n_734), .Y(n_904) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_67), .A2(n_202), .B1(n_346), .B2(n_495), .C1(n_536), .C2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_68), .A2(n_248), .B1(n_469), .B2(n_791), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_69), .A2(n_130), .B1(n_575), .B2(n_576), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_70), .A2(n_238), .B1(n_610), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_71), .A2(n_109), .B1(n_741), .B2(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_72), .A2(n_330), .B1(n_471), .B2(n_472), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_73), .A2(n_112), .B1(n_507), .B2(n_547), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_74), .A2(n_301), .B1(n_468), .B2(n_469), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_75), .A2(n_150), .B1(n_870), .B2(n_872), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_76), .A2(n_297), .B1(n_436), .B2(n_542), .Y(n_541) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_78), .A2(n_207), .B1(n_411), .B2(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_80), .A2(n_329), .B1(n_519), .B2(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_81), .B(n_534), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_82), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_83), .A2(n_169), .B1(n_469), .B2(n_791), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_84), .A2(n_283), .B1(n_675), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_85), .A2(n_194), .B1(n_484), .B2(n_597), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_87), .A2(n_339), .B1(n_436), .B2(n_542), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_88), .A2(n_176), .B1(n_490), .B2(n_492), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_89), .A2(n_172), .B1(n_606), .B2(n_607), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_90), .A2(n_334), .B1(n_464), .B2(n_465), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_91), .A2(n_266), .B1(n_458), .B2(n_553), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_92), .B(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_95), .A2(n_249), .B1(n_515), .B2(n_555), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_96), .A2(n_278), .B1(n_464), .B2(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_97), .A2(n_288), .B1(n_504), .B2(n_993), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_98), .A2(n_379), .B1(n_490), .B2(n_731), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_99), .A2(n_229), .B1(n_492), .B2(n_537), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_100), .A2(n_247), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_101), .A2(n_126), .B1(n_522), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_102), .A2(n_209), .B1(n_596), .B2(n_597), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_103), .A2(n_303), .B1(n_490), .B2(n_492), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_104), .B(n_534), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_105), .A2(n_179), .B1(n_582), .B2(n_912), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_107), .A2(n_148), .B1(n_458), .B2(n_462), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_108), .A2(n_281), .B1(n_592), .B2(n_960), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_110), .A2(n_221), .B1(n_512), .B2(n_515), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_111), .A2(n_235), .B1(n_507), .B2(n_552), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g808 ( .A1(n_113), .A2(n_318), .B1(n_781), .B2(n_782), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_115), .A2(n_242), .B1(n_817), .B2(n_818), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_116), .A2(n_340), .B1(n_448), .B2(n_453), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_117), .A2(n_302), .B1(n_604), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_118), .A2(n_341), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_121), .A2(n_987), .B1(n_988), .B2(n_1004), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_121), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_122), .A2(n_152), .B1(n_436), .B2(n_735), .Y(n_885) );
OAI22x1_ASAP7_75t_L g955 ( .A1(n_123), .A2(n_956), .B1(n_957), .B2(n_971), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_123), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_124), .A2(n_253), .B1(n_515), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_127), .A2(n_196), .B1(n_521), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_129), .A2(n_332), .B1(n_500), .B2(n_582), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_131), .A2(n_325), .B1(n_482), .B2(n_734), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_132), .A2(n_342), .B1(n_547), .B2(n_659), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_133), .A2(n_307), .B1(n_641), .B2(n_706), .Y(n_765) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_134), .A2(n_289), .B1(n_411), .B2(n_412), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_135), .A2(n_212), .B1(n_519), .B2(n_949), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_136), .A2(n_158), .B1(n_604), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_137), .A2(n_217), .B1(n_610), .B2(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_138), .A2(n_320), .B1(n_500), .B2(n_504), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_141), .A2(n_270), .B1(n_504), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_142), .A2(n_159), .B1(n_531), .B2(n_576), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_143), .A2(n_168), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_144), .A2(n_365), .B1(n_670), .B2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_145), .A2(n_311), .B1(n_636), .B2(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_146), .A2(n_335), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_147), .A2(n_355), .B1(n_613), .B2(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_149), .B(n_534), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_153), .A2(n_322), .B1(n_408), .B2(n_682), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_154), .A2(n_299), .B1(n_468), .B2(n_469), .Y(n_848) );
XOR2x2_ASAP7_75t_L g621 ( .A(n_155), .B(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_156), .A2(n_251), .B1(n_490), .B2(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_157), .A2(n_368), .B1(n_868), .B2(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_160), .A2(n_323), .B1(n_469), .B2(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_161), .A2(n_315), .B1(n_484), .B2(n_597), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_162), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_163), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_164), .A2(n_185), .B1(n_530), .B2(n_532), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_165), .A2(n_234), .B1(n_761), .B2(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_166), .B(n_495), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_167), .A2(n_273), .B1(n_519), .B2(n_547), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_170), .A2(n_268), .B1(n_606), .B2(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_171), .A2(n_227), .B1(n_471), .B2(n_472), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_173), .A2(n_189), .B1(n_817), .B2(n_818), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_174), .A2(n_274), .B1(n_606), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_175), .A2(n_360), .B1(n_781), .B2(n_782), .Y(n_780) );
OA22x2_ASAP7_75t_L g882 ( .A1(n_177), .A2(n_883), .B1(n_896), .B2(n_897), .Y(n_882) );
INVx1_ASAP7_75t_L g896 ( .A(n_177), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_178), .A2(n_218), .B1(n_515), .B2(n_555), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_180), .A2(n_262), .B1(n_604), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_181), .A2(n_367), .B1(n_436), .B2(n_482), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_182), .A2(n_236), .B1(n_505), .B2(n_606), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_183), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_184), .A2(n_243), .B1(n_641), .B2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_186), .A2(n_290), .B1(n_603), .B2(n_667), .Y(n_666) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_187), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_188), .A2(n_357), .B1(n_464), .B2(n_465), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_190), .A2(n_222), .B1(n_471), .B2(n_472), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_191), .Y(n_451) );
AOI22x1_ASAP7_75t_SL g750 ( .A1(n_192), .A2(n_751), .B1(n_752), .B2(n_766), .Y(n_750) );
INVx1_ASAP7_75t_L g766 ( .A(n_192), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_193), .A2(n_244), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_197), .A2(n_233), .B1(n_507), .B2(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_198), .B(n_495), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_199), .A2(n_246), .B1(n_555), .B2(n_793), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_203), .A2(n_333), .B1(n_670), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_204), .A2(n_294), .B1(n_537), .B2(n_731), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_206), .A2(n_374), .B1(n_471), .B2(n_472), .Y(n_927) );
INVx1_ASAP7_75t_L g983 ( .A(n_207), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_208), .A2(n_269), .B1(n_453), .B2(n_784), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_211), .A2(n_364), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_216), .A2(n_370), .B1(n_550), .B2(n_582), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_219), .A2(n_377), .B1(n_611), .B2(n_636), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_220), .A2(n_375), .B1(n_408), .B2(n_424), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_223), .A2(n_240), .B1(n_492), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_224), .A2(n_381), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g390 ( .A(n_225), .Y(n_390) );
XOR2x2_ASAP7_75t_L g526 ( .A(n_226), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_228), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_231), .A2(n_255), .B1(n_464), .B2(n_465), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_232), .A2(n_349), .B1(n_481), .B2(n_599), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_237), .A2(n_312), .B1(n_469), .B2(n_791), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_241), .A2(n_336), .B1(n_453), .B2(n_784), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_245), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_258), .A2(n_280), .B1(n_519), .B2(n_521), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_260), .A2(n_267), .B1(n_500), .B2(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_261), .A2(n_1009), .B1(n_1010), .B2(n_1026), .Y(n_1008) );
INVx1_ASAP7_75t_L g1026 ( .A(n_261), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_263), .B(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_264), .A2(n_356), .B1(n_462), .B2(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_275), .A2(n_328), .B1(n_536), .B2(n_538), .Y(n_535) );
OA22x2_ASAP7_75t_L g661 ( .A1(n_276), .A2(n_662), .B1(n_663), .B2(n_683), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_276), .Y(n_662) );
AO21x2_ASAP7_75t_L g686 ( .A1(n_276), .A2(n_663), .B(n_687), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g800 ( .A(n_277), .B(n_801), .Y(n_800) );
XNOR2x1_ASAP7_75t_L g588 ( .A(n_282), .B(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_286), .A2(n_291), .B1(n_531), .B2(n_542), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_287), .A2(n_348), .B1(n_700), .B2(n_701), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_289), .B(n_982), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_293), .A2(n_317), .B1(n_458), .B2(n_465), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_295), .B(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_296), .A2(n_371), .B1(n_781), .B2(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_300), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_304), .A2(n_319), .B1(n_522), .B2(n_641), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_306), .A2(n_376), .B1(n_703), .B2(n_967), .Y(n_966) );
OA22x2_ASAP7_75t_L g402 ( .A1(n_308), .A2(n_403), .B1(n_404), .B2(n_474), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_308), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_309), .A2(n_327), .B1(n_582), .B2(n_761), .Y(n_893) );
INVx3_ASAP7_75t_L g411 ( .A(n_310), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_314), .A2(n_353), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_321), .A2(n_331), .B1(n_492), .B2(n_592), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_326), .A2(n_372), .B1(n_599), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_338), .A2(n_380), .B1(n_481), .B2(n_868), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_343), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_344), .B(n_569), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_345), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_347), .B(n_569), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_358), .B(n_569), .Y(n_600) );
OAI22x1_ASAP7_75t_L g935 ( .A1(n_361), .A2(n_936), .B1(n_937), .B2(n_954), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_361), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_362), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_363), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g979 ( .A(n_363), .Y(n_979) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
AND2x2_ASAP7_75t_R g1006 ( .A(n_366), .B(n_979), .Y(n_1006) );
INVxp67_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
XNOR2xp5_ASAP7_75t_L g855 ( .A(n_373), .B(n_856), .Y(n_855) );
XOR2x2_ASAP7_75t_L g725 ( .A(n_378), .B(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_385), .B(n_387), .Y(n_1030) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_386), .B(n_979), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_770), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g975 ( .A1(n_392), .A2(n_770), .B(n_976), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_618), .B2(n_769), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_561), .B2(n_617), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_525), .B1(n_558), .B2(n_559), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_475), .Y(n_398) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_399), .A2(n_475), .B(n_556), .Y(n_558) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_400), .A2(n_694), .B1(n_718), .B2(n_719), .Y(n_693) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g557 ( .A(n_402), .Y(n_557) );
INVx1_ASAP7_75t_L g474 ( .A(n_404), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_455), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_433), .C(n_445), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_427), .Y(n_406) );
INVx1_ASAP7_75t_SL g681 ( .A(n_408), .Y(n_681) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_416), .Y(n_408) );
AND2x2_ASAP7_75t_L g448 ( .A(n_409), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g462 ( .A(n_409), .B(n_461), .Y(n_462) );
AND2x4_ASAP7_75t_L g485 ( .A(n_409), .B(n_449), .Y(n_485) );
AND2x2_ASAP7_75t_L g491 ( .A(n_409), .B(n_416), .Y(n_491) );
AND2x2_ASAP7_75t_L g784 ( .A(n_409), .B(n_449), .Y(n_784) );
AND2x2_ASAP7_75t_L g818 ( .A(n_409), .B(n_461), .Y(n_818) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
AND2x2_ASAP7_75t_L g426 ( .A(n_410), .B(n_414), .Y(n_426) );
INVx1_ASAP7_75t_L g432 ( .A(n_410), .Y(n_432) );
INVx1_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
INVx2_ASAP7_75t_L g412 ( .A(n_411), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_411), .Y(n_415) );
OAI22x1_ASAP7_75t_L g417 ( .A1(n_411), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_411), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
AND2x4_ASAP7_75t_L g431 ( .A(n_413), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_414), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g437 ( .A(n_416), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g468 ( .A(n_416), .B(n_431), .Y(n_468) );
AND2x4_ASAP7_75t_L g509 ( .A(n_416), .B(n_431), .Y(n_509) );
AND2x4_ASAP7_75t_L g781 ( .A(n_416), .B(n_438), .Y(n_781) );
AND2x2_ASAP7_75t_L g791 ( .A(n_416), .B(n_431), .Y(n_791) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_421), .Y(n_416) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_417), .Y(n_425) );
AND2x2_ASAP7_75t_L g430 ( .A(n_417), .B(n_422), .Y(n_430) );
INVx2_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
AND2x4_ASAP7_75t_L g461 ( .A(n_421), .B(n_450), .Y(n_461) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g449 ( .A(n_422), .B(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g473 ( .A(n_422), .Y(n_473) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x2_ASAP7_75t_L g493 ( .A(n_425), .B(n_426), .Y(n_493) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_425), .B(n_426), .Y(n_682) );
AND2x4_ASAP7_75t_L g469 ( .A(n_426), .B(n_461), .Y(n_469) );
AND2x4_ASAP7_75t_L g472 ( .A(n_426), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g505 ( .A(n_426), .B(n_473), .Y(n_505) );
AND2x4_ASAP7_75t_L g522 ( .A(n_426), .B(n_461), .Y(n_522) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g804 ( .A(n_429), .Y(n_804) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AND2x4_ASAP7_75t_L g442 ( .A(n_430), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g453 ( .A(n_430), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g488 ( .A(n_430), .B(n_454), .Y(n_488) );
AND2x2_ASAP7_75t_L g497 ( .A(n_430), .B(n_431), .Y(n_497) );
AND2x2_ASAP7_75t_L g675 ( .A(n_430), .B(n_454), .Y(n_675) );
AND2x2_ASAP7_75t_L g782 ( .A(n_430), .B(n_443), .Y(n_782) );
AND2x2_ASAP7_75t_L g844 ( .A(n_430), .B(n_443), .Y(n_844) );
AND2x4_ASAP7_75t_L g460 ( .A(n_431), .B(n_461), .Y(n_460) );
AND2x6_ASAP7_75t_L g464 ( .A(n_431), .B(n_449), .Y(n_464) );
AND2x2_ASAP7_75t_L g514 ( .A(n_431), .B(n_449), .Y(n_514) );
AND2x2_ASAP7_75t_L g817 ( .A(n_431), .B(n_461), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_440), .B2(n_441), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_SL g709 ( .A(n_436), .Y(n_709) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
INVx3_ASAP7_75t_L g678 ( .A(n_437), .Y(n_678) );
AND2x6_ASAP7_75t_L g465 ( .A(n_438), .B(n_461), .Y(n_465) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_438), .B(n_449), .Y(n_471) );
AND2x2_ASAP7_75t_L g503 ( .A(n_438), .B(n_449), .Y(n_503) );
AND2x4_ASAP7_75t_L g517 ( .A(n_438), .B(n_461), .Y(n_517) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_439), .Y(n_444) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx4f_ASAP7_75t_L g482 ( .A(n_442), .Y(n_482) );
INVx2_ASAP7_75t_L g544 ( .A(n_442), .Y(n_544) );
BUFx3_ASAP7_75t_L g599 ( .A(n_442), .Y(n_599) );
BUFx6f_ASAP7_75t_SL g735 ( .A(n_442), .Y(n_735) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_451), .B2(n_452), .Y(n_445) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_463), .Y(n_456) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx4_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
INVx2_ASAP7_75t_SL g636 ( .A(n_459), .Y(n_636) );
INVx2_ASAP7_75t_L g700 ( .A(n_459), .Y(n_700) );
INVx3_ASAP7_75t_SL g863 ( .A(n_459), .Y(n_863) );
INVx2_ASAP7_75t_SL g947 ( .A(n_459), .Y(n_947) );
INVx8_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx3_ASAP7_75t_L g510 ( .A(n_462), .Y(n_510) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_462), .Y(n_553) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_462), .Y(n_611) );
INVx2_ASAP7_75t_L g671 ( .A(n_462), .Y(n_671) );
INVx1_ASAP7_75t_L g829 ( .A(n_464), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_477), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
NOR2xp67_ASAP7_75t_L g478 ( .A(n_479), .B(n_498), .Y(n_478) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .C(n_489), .D(n_494), .Y(n_479) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
BUFx3_ASAP7_75t_L g596 ( .A(n_485), .Y(n_596) );
BUFx2_ASAP7_75t_L g940 ( .A(n_485), .Y(n_940) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g532 ( .A(n_487), .Y(n_532) );
INVx2_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
INVx2_ASAP7_75t_L g597 ( .A(n_487), .Y(n_597) );
INVx2_ASAP7_75t_SL g710 ( .A(n_487), .Y(n_710) );
INVx6_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx5_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g537 ( .A(n_491), .Y(n_537) );
INVx2_ASAP7_75t_L g593 ( .A(n_491), .Y(n_593) );
BUFx3_ASAP7_75t_L g714 ( .A(n_491), .Y(n_714) );
INVx2_ASAP7_75t_L g871 ( .A(n_492), .Y(n_871) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_492), .Y(n_1003) );
BUFx12f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g540 ( .A(n_493), .Y(n_540) );
BUFx2_ASAP7_75t_L g534 ( .A(n_495), .Y(n_534) );
INVx4_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_SL g569 ( .A(n_496), .Y(n_569) );
BUFx2_ASAP7_75t_L g625 ( .A(n_496), .Y(n_625) );
INVx3_ASAP7_75t_SL g889 ( .A(n_496), .Y(n_889) );
INVx3_ASAP7_75t_L g943 ( .A(n_496), .Y(n_943) );
INVx6_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_499), .B(n_506), .C(n_511), .D(n_518), .Y(n_498) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g968 ( .A(n_501), .Y(n_968) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
INVx1_ASAP7_75t_L g761 ( .A(n_502), .Y(n_761) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_503), .Y(n_606) );
BUFx3_ASAP7_75t_L g912 ( .A(n_503), .Y(n_912) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g582 ( .A(n_505), .Y(n_582) );
INVx5_ASAP7_75t_SL g608 ( .A(n_505), .Y(n_608) );
BUFx3_ASAP7_75t_L g825 ( .A(n_505), .Y(n_825) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
INVx3_ASAP7_75t_L g610 ( .A(n_508), .Y(n_610) );
INVx2_ASAP7_75t_L g859 ( .A(n_508), .Y(n_859) );
INVx6_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g641 ( .A(n_509), .Y(n_641) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_SL g555 ( .A(n_513), .Y(n_555) );
INVx3_ASAP7_75t_L g603 ( .A(n_513), .Y(n_603) );
INVx2_ASAP7_75t_L g741 ( .A(n_513), .Y(n_741) );
INVx2_ASAP7_75t_L g914 ( .A(n_513), .Y(n_914) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g639 ( .A(n_514), .Y(n_639) );
BUFx2_ASAP7_75t_L g698 ( .A(n_514), .Y(n_698) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g586 ( .A(n_516), .Y(n_586) );
INVx2_ASAP7_75t_L g604 ( .A(n_516), .Y(n_604) );
INVx2_ASAP7_75t_L g667 ( .A(n_516), .Y(n_667) );
INVx2_ASAP7_75t_L g742 ( .A(n_516), .Y(n_742) );
INVx2_ASAP7_75t_SL g764 ( .A(n_516), .Y(n_764) );
INVx2_ASAP7_75t_L g910 ( .A(n_516), .Y(n_910) );
INVx1_ASAP7_75t_SL g949 ( .A(n_516), .Y(n_949) );
INVx8_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g660 ( .A(n_520), .Y(n_660) );
BUFx2_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_SL g547 ( .A(n_522), .Y(n_547) );
BUFx3_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
BUFx3_ASAP7_75t_L g706 ( .A(n_522), .Y(n_706) );
INVx2_ASAP7_75t_L g746 ( .A(n_522), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_556), .Y(n_525) );
INVx5_ASAP7_75t_L g560 ( .A(n_526), .Y(n_560) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_545), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .C(n_535), .D(n_541), .Y(n_528) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx4f_ASAP7_75t_SL g575 ( .A(n_531), .Y(n_575) );
BUFx6f_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g651 ( .A(n_537), .Y(n_651) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g594 ( .A(n_540), .Y(n_594) );
INVx2_ASAP7_75t_L g731 ( .A(n_540), .Y(n_731) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g868 ( .A(n_544), .Y(n_868) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .C(n_551), .D(n_554), .Y(n_545) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g720 ( .A(n_557), .Y(n_720) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_587), .B1(n_588), .B2(n_614), .Y(n_563) );
INVx1_ASAP7_75t_SL g615 ( .A(n_565), .Y(n_615) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_577), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_572), .Y(n_566) );
OAI21xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_571), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_568), .A2(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_601), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g590 ( .A(n_591), .B(n_595), .C(n_598), .D(n_600), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g628 ( .A(n_593), .Y(n_628) );
BUFx2_ASAP7_75t_L g712 ( .A(n_594), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .C(n_609), .D(n_612), .Y(n_601) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_606), .Y(n_861) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g703 ( .A(n_608), .Y(n_703) );
INVx3_ASAP7_75t_L g762 ( .A(n_608), .Y(n_762) );
INVx2_ASAP7_75t_L g953 ( .A(n_608), .Y(n_953) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_611), .Y(n_865) );
INVx1_ASAP7_75t_L g769 ( .A(n_618), .Y(n_769) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_691), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_642), .B1(n_689), .B2(n_690), .Y(n_619) );
INVx1_ASAP7_75t_L g689 ( .A(n_620), .Y(n_689) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2x1_ASAP7_75t_SL g622 ( .A(n_623), .B(n_632), .Y(n_622) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_629), .Y(n_623) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_627), .Y(n_624) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_628), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_637), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g690 ( .A(n_642), .Y(n_690) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_661), .B1(n_684), .B2(n_685), .Y(n_644) );
INVx1_ASAP7_75t_SL g684 ( .A(n_645), .Y(n_684) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_654), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .C(n_652), .D(n_653), .Y(n_647) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_657), .D(n_658), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22x1_ASAP7_75t_SL g748 ( .A1(n_661), .A2(n_685), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_662), .Y(n_688) );
INVx1_ASAP7_75t_L g683 ( .A(n_663), .Y(n_683) );
NOR2x1_ASAP7_75t_SL g687 ( .A(n_663), .B(n_688), .Y(n_687) );
NAND4xp75_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .C(n_673), .D(n_679), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_670), .Y(n_701) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g793 ( .A(n_671), .Y(n_793) );
INVx1_ASAP7_75t_L g1020 ( .A(n_671), .Y(n_1020) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx2_ASAP7_75t_SL g997 ( .A(n_677), .Y(n_997) );
INVx4_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g734 ( .A(n_678), .Y(n_734) );
INVx1_ASAP7_75t_L g1014 ( .A(n_678), .Y(n_1014) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
XOR2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_721), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g718 ( .A(n_694), .Y(n_718) );
XNOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_717), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_696), .B(n_707), .Y(n_695) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .C(n_702), .D(n_704), .Y(n_696) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .C(n_715), .D(n_716), .Y(n_707) );
INVx1_ASAP7_75t_L g1024 ( .A(n_712), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OA22x2_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_748), .B1(n_767), .B2(n_768), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g767 ( .A(n_724), .Y(n_767) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_737), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_732), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_743), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g951 ( .A(n_746), .Y(n_951) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_748), .Y(n_768) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .Y(n_752) );
NAND4xp25_ASAP7_75t_SL g753 ( .A(n_754), .B(n_755), .C(n_756), .D(n_757), .Y(n_753) );
NAND4xp25_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .C(n_763), .D(n_765), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_876), .B2(n_974), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_795), .Y(n_772) );
XOR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_794), .Y(n_773) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_785), .Y(n_774) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_783), .Y(n_779) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_789), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_854), .B2(n_875), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI22x1_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_819), .B1(n_852), .B2(n_853), .Y(n_797) );
INVx1_ASAP7_75t_L g853 ( .A(n_798), .Y(n_853) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_802), .B(n_810), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_807), .Y(n_802) );
OAI21xp5_ASAP7_75t_SL g803 ( .A1(n_804), .A2(n_805), .B(n_806), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx2_ASAP7_75t_L g852 ( .A(n_819), .Y(n_852) );
AO22x2_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_836), .B1(n_850), .B2(n_851), .Y(n_819) );
INVx1_ASAP7_75t_SL g850 ( .A(n_820), .Y(n_850) );
XNOR2x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
OR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_831), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g823 ( .A(n_824), .B(n_826), .C(n_827), .D(n_830), .Y(n_823) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g892 ( .A(n_829), .Y(n_892) );
NAND4xp25_ASAP7_75t_SL g831 ( .A(n_832), .B(n_833), .C(n_834), .D(n_835), .Y(n_831) );
INVx2_ASAP7_75t_SL g851 ( .A(n_836), .Y(n_851) );
XNOR2x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_839), .B(n_845), .Y(n_838) );
NAND4xp25_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .C(n_842), .D(n_843), .Y(n_839) );
NAND4xp25_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .C(n_848), .D(n_849), .Y(n_845) );
INVx2_ASAP7_75t_SL g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_855), .Y(n_875) );
NOR2xp67_ASAP7_75t_L g856 ( .A(n_857), .B(n_866), .Y(n_856) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .C(n_862), .D(n_864), .Y(n_857) );
NAND4xp25_ASAP7_75t_L g866 ( .A(n_867), .B(n_869), .C(n_873), .D(n_874), .Y(n_866) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g974 ( .A(n_876), .Y(n_974) );
XNOR2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_934), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_898), .B1(n_899), .B2(n_933), .Y(n_880) );
INVx2_ASAP7_75t_L g933 ( .A(n_881), .Y(n_933) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g897 ( .A(n_883), .Y(n_897) );
NOR2x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_890), .Y(n_883) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .C(n_887), .D(n_888), .Y(n_884) );
BUFx6f_ASAP7_75t_L g960 ( .A(n_889), .Y(n_960) );
NAND4xp25_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .C(n_894), .D(n_895), .Y(n_890) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
XNOR2x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_917), .Y(n_899) );
INVx1_ASAP7_75t_SL g901 ( .A(n_902), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_908), .Y(n_902) );
NAND4xp25_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .C(n_906), .D(n_907), .Y(n_903) );
NAND4xp25_ASAP7_75t_L g908 ( .A(n_909), .B(n_911), .C(n_913), .D(n_915), .Y(n_908) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
XOR2x2_ASAP7_75t_L g918 ( .A(n_919), .B(n_932), .Y(n_918) );
NAND2x1_ASAP7_75t_L g919 ( .A(n_920), .B(n_925), .Y(n_919) );
NOR2x1_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
NOR2x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_929), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_955), .B1(n_972), .B2(n_973), .Y(n_934) );
INVx1_ASAP7_75t_L g973 ( .A(n_935), .Y(n_973) );
INVx2_ASAP7_75t_L g954 ( .A(n_937), .Y(n_954) );
OR2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_945), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g938 ( .A(n_939), .B(n_941), .C(n_942), .D(n_944), .Y(n_938) );
NAND4xp25_ASAP7_75t_L g945 ( .A(n_946), .B(n_948), .C(n_950), .D(n_952), .Y(n_945) );
INVx1_ASAP7_75t_L g972 ( .A(n_955), .Y(n_972) );
INVx2_ASAP7_75t_SL g971 ( .A(n_957), .Y(n_971) );
OR2x2_ASAP7_75t_L g957 ( .A(n_958), .B(n_964), .Y(n_957) );
NAND4xp25_ASAP7_75t_SL g958 ( .A(n_959), .B(n_961), .C(n_962), .D(n_963), .Y(n_958) );
NAND4xp25_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .C(n_969), .D(n_970), .Y(n_964) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g993 ( .A(n_968), .Y(n_993) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_978), .B(n_980), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_978), .B(n_981), .Y(n_1029) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_983), .B(n_984), .Y(n_982) );
OAI222xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_1005), .B1(n_1007), .B2(n_1026), .C1(n_1027), .C2(n_1030), .Y(n_985) );
CKINVDCx16_ASAP7_75t_R g987 ( .A(n_988), .Y(n_987) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NAND4xp75_ASAP7_75t_L g989 ( .A(n_990), .B(n_994), .C(n_999), .D(n_1002), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_998), .Y(n_994) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
AND2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
INVx1_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
NOR3xp33_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1016), .C(n_1022), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .Y(n_1011) );
BUFx3_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NAND4xp25_ASAP7_75t_SL g1016 ( .A(n_1017), .B(n_1018), .C(n_1019), .D(n_1021), .Y(n_1016) );
OAI21xp5_ASAP7_75t_SL g1022 ( .A1(n_1023), .A2(n_1024), .B(n_1025), .Y(n_1022) );
INVx1_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
CKINVDCx6p67_ASAP7_75t_R g1028 ( .A(n_1029), .Y(n_1028) );
endmodule