module fake_jpeg_18795_n_218 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_218);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_40),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_23),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_25),
.B1(n_27),
.B2(n_15),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_16),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_16),
.C(n_19),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_13),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_27),
.B1(n_15),
.B2(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_20),
.B1(n_30),
.B2(n_0),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_55),
.B1(n_47),
.B2(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_79),
.B1(n_83),
.B2(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_41),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_14),
.B(n_22),
.C(n_28),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_74),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_13),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_84),
.B(n_20),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_81),
.Y(n_125)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_90),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_19),
.B1(n_26),
.B2(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_34),
.B1(n_19),
.B2(n_26),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_13),
.Y(n_84)
);

INVx2_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_89),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_16),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_17),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_17),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_47),
.B(n_20),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_113),
.B1(n_124),
.B2(n_126),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_80),
.B1(n_67),
.B2(n_66),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_78),
.B1(n_90),
.B2(n_70),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_94),
.B1(n_84),
.B2(n_95),
.Y(n_132)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_96),
.Y(n_136)
);

XOR2x2_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_106),
.B1(n_114),
.B2(n_118),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_140),
.B1(n_124),
.B2(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_71),
.B(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_68),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_68),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_102),
.B1(n_95),
.B2(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_99),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_77),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_165),
.B1(n_131),
.B2(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_164),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_120),
.B1(n_115),
.B2(n_117),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_133),
.B1(n_132),
.B2(n_141),
.Y(n_174)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_129),
.C(n_105),
.D(n_122),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_125),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_127),
.B1(n_120),
.B2(n_117),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_123),
.B1(n_104),
.B2(n_116),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_122),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_141),
.B(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_134),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_130),
.B(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_180),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_131),
.B1(n_116),
.B2(n_97),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_104),
.C(n_82),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_158),
.C(n_162),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_151),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_185),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_164),
.A3(n_154),
.B1(n_165),
.B2(n_101),
.C1(n_162),
.C2(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_154),
.C(n_163),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_194),
.B1(n_188),
.B2(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_177),
.B1(n_180),
.B2(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_174),
.B1(n_175),
.B2(n_179),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_186),
.B1(n_144),
.B2(n_1),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_176),
.B1(n_163),
.B2(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_176),
.B(n_2),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_188),
.B(n_5),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_185),
.B1(n_182),
.B2(n_183),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_206),
.B(n_202),
.Y(n_208)
);

OAI222xp33_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.C1(n_186),
.C2(n_10),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_208),
.B1(n_205),
.B2(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_201),
.B(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_215),
.C(n_8),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_12),
.Y(n_218)
);


endmodule