module fake_jpeg_2633_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_41),
.B(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_62),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_43),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_2),
.C(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_67),
.B1(n_74),
.B2(n_55),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_74),
.B(n_55),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_41),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_101),
.B1(n_104),
.B2(n_78),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_98),
.B(n_78),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_49),
.B(n_46),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_67),
.B1(n_46),
.B2(n_42),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_6),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_8),
.C(n_9),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_79),
.B1(n_82),
.B2(n_76),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_118),
.B1(n_119),
.B2(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_21),
.C(n_37),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_29),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_20),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_15),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_96),
.B1(n_98),
.B2(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_16),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_24),
.B(n_36),
.C(n_35),
.D(n_34),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_31),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_28),
.B(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_14),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_115),
.C(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_38),
.B1(n_122),
.B2(n_132),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_140),
.B1(n_121),
.B2(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_145),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_131),
.B(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_134),
.C(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_132),
.B1(n_142),
.B2(n_127),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_156),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_150),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_138),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_149),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_156),
.C(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_147),
.C(n_144),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_143),
.Y(n_165)
);


endmodule