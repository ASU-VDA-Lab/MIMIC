module fake_netlist_6_3456_n_3111 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_3111);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_3111;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_461;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_3106;
wire n_2630;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2739;
wire n_2480;
wire n_3023;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_423;
wire n_1865;
wire n_586;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_928;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1317;
wire n_1082;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_462;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_2932;
wire n_1767;
wire n_627;
wire n_595;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3037;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_716;
wire n_623;
wire n_1475;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_1048;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_527;
wire n_683;
wire n_1207;
wire n_474;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2581;
wire n_1363;
wire n_2294;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_444;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_3109;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_664;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_1409;
wire n_504;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_3105;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2699;
wire n_2272;
wire n_2200;
wire n_3029;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_972;
wire n_1406;
wire n_456;
wire n_2766;
wire n_2670;
wire n_1332;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_3045;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_799;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_706;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_430;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_2833;
wire n_1113;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_841;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_2969;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1785;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1114;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2743;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_3035;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_2802;
wire n_1085;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_2600;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_3038;
wire n_859;
wire n_570;
wire n_2033;
wire n_3086;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_3095;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_190),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_153),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_140),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_313),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_235),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_174),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_231),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_352),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_184),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_197),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_373),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_293),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_35),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_256),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_115),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_315),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_70),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_23),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_34),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_14),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_189),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_150),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_262),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_391),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_216),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_350),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_296),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_49),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_146),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_4),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_225),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_32),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_242),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_207),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_18),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_142),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_22),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_205),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_385),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_37),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_72),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_263),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_192),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_160),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_232),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_150),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_139),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_59),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_89),
.Y(n_472)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_8),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_348),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_52),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_90),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_257),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_405),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_70),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_321),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_135),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_134),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_58),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_44),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_376),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_33),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_261),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_120),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_105),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_164),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g491 ( 
.A(n_191),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_299),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_198),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_105),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_84),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_140),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_49),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_186),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_319),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_174),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_278),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_404),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_139),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_332),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_270),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_87),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_155),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_308),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_37),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_108),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_294),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_344),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_269),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_289),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_39),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_383),
.Y(n_518)
);

CKINVDCx6p67_ASAP7_75t_R g519 ( 
.A(n_124),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_149),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_103),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_116),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_217),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_239),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_283),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_152),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_172),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_154),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_118),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_378),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_366),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_298),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_417),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_295),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_333),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_181),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_310),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_274),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_309),
.Y(n_540)
);

BUFx5_ASAP7_75t_L g541 ( 
.A(n_55),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_142),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_403),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_73),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_38),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_91),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_14),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_402),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_128),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_178),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_106),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_62),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_264),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_358),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_117),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_397),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_161),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_97),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_32),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_72),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_416),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_22),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_317),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_53),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_185),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_233),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_144),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_190),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_209),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_389),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_355),
.Y(n_571)
);

BUFx2_ASAP7_75t_SL g572 ( 
.A(n_284),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_282),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_271),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_304),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_34),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_59),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_192),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_9),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_137),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_63),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_155),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_224),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_414),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_111),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_11),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_27),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_349),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_52),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_164),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_392),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_351),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_86),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_335),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_212),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_171),
.Y(n_596)
);

BUFx5_ASAP7_75t_L g597 ( 
.A(n_372),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_388),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_85),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_26),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_136),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_149),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_29),
.Y(n_603)
);

CKINVDCx14_ASAP7_75t_R g604 ( 
.A(n_194),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_285),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_124),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_44),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_322),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_83),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_87),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_158),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_81),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_387),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_287),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_211),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_96),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_144),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_381),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_260),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_325),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_290),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_328),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_40),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_395),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_33),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_24),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_30),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_166),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_99),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_110),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_254),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_18),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_177),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_85),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_380),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_363),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_206),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_252),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_251),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_113),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_143),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_16),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_222),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_258),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_77),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_54),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_390),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_147),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_54),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_347),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_367),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_221),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_9),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_168),
.Y(n_654)
);

BUFx5_ASAP7_75t_L g655 ( 
.A(n_101),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_130),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_1),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_243),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_314),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_96),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_93),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_48),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_245),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_368),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_82),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_134),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_167),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_178),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_75),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_318),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_200),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_152),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_326),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_246),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_361),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_250),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_194),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_21),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_39),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_241),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_229),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_419),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_31),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_272),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_266),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_135),
.Y(n_686)
);

CKINVDCx14_ASAP7_75t_R g687 ( 
.A(n_130),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_273),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_28),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_26),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_183),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_329),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_411),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_228),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_277),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_183),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_371),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_8),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_191),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_214),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_303),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_398),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_167),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_182),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_359),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_82),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_301),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_353),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_208),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_5),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_306),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_320),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_384),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_365),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_374),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_400),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_195),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_66),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_141),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_176),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_170),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_408),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_123),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_157),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_57),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_327),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_473),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_473),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_473),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_473),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_473),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_473),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_473),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_425),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_566),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_465),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_432),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_712),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_473),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_491),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_491),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_491),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_625),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_491),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_491),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_465),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_491),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_491),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_478),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_604),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_427),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_531),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_491),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_687),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_677),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_541),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_541),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_541),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_555),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_541),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_543),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_632),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_519),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_519),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_541),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_478),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_486),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_488),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_518),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_494),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_495),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_541),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_541),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_518),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_541),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_655),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_496),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_421),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_497),
.Y(n_781)
);

INVxp33_ASAP7_75t_SL g782 ( 
.A(n_421),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_655),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_584),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_423),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_655),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_655),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_655),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_509),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_426),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_655),
.Y(n_791)
);

CKINVDCx16_ASAP7_75t_R g792 ( 
.A(n_526),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_655),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_550),
.Y(n_794)
);

INVxp33_ASAP7_75t_SL g795 ( 
.A(n_429),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_441),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_441),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_550),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_500),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_622),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_599),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_599),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_633),
.Y(n_803)
);

CKINVDCx16_ASAP7_75t_R g804 ( 
.A(n_525),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_633),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_555),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_658),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_503),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_441),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_536),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_441),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_441),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_581),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_581),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_538),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_581),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_581),
.Y(n_817)
);

CKINVDCx14_ASAP7_75t_R g818 ( 
.A(n_555),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_581),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_438),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_440),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_455),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_458),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_597),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_466),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_597),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_680),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_472),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_475),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_485),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_476),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_597),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_483),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_489),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_490),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_529),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_506),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_507),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_510),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_546),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_560),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_516),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_520),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_536),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_429),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_498),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_521),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_565),
.Y(n_848)
);

INVxp33_ASAP7_75t_SL g849 ( 
.A(n_434),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_498),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_511),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_511),
.Y(n_852)
);

INVxp33_ASAP7_75t_SL g853 ( 
.A(n_434),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_545),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_487),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_545),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_567),
.B(n_0),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_597),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_597),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_582),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_585),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_587),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_436),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_522),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_564),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_493),
.Y(n_866)
);

OAI22x1_ASAP7_75t_SL g867 ( 
.A1(n_763),
.A2(n_452),
.B1(n_482),
.B2(n_442),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_815),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_797),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_747),
.B(n_542),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_750),
.B(n_542),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_751),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_741),
.A2(n_639),
.B(n_445),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_796),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_815),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_815),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_797),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_815),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_743),
.A2(n_645),
.B1(n_656),
.B2(n_484),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_796),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_816),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_815),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_816),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_809),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_741),
.A2(n_639),
.B(n_445),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_811),
.Y(n_886)
);

OA21x2_ASAP7_75t_L g887 ( 
.A1(n_729),
.A2(n_517),
.B(n_437),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_812),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_813),
.B(n_624),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_763),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_737),
.A2(n_439),
.B1(n_443),
.B2(n_436),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_814),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_751),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_817),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_767),
.B(n_624),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_768),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_742),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_729),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_755),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_730),
.B(n_639),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_774),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_774),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_738),
.B(n_502),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_727),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_728),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_739),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_740),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_770),
.B(n_502),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_730),
.B(n_594),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_775),
.B(n_594),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_734),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_736),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_731),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_731),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_732),
.B(n_538),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_732),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_778),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_783),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_733),
.A2(n_517),
.B(n_437),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_733),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_786),
.Y(n_922)
);

NOR2x1_ASAP7_75t_L g923 ( 
.A(n_830),
.B(n_572),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_735),
.A2(n_710),
.B1(n_723),
.B2(n_690),
.Y(n_924)
);

AND2x2_ASAP7_75t_SL g925 ( 
.A(n_857),
.B(n_524),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_768),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_855),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_787),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_755),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_745),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_810),
.B(n_564),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_788),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_866),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_745),
.B(n_708),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_746),
.B(n_708),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_844),
.B(n_601),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_791),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_746),
.Y(n_938)
);

OAI22x1_ASAP7_75t_L g939 ( 
.A1(n_760),
.A2(n_443),
.B1(n_451),
.B2(n_439),
.Y(n_939)
);

OA21x2_ASAP7_75t_L g940 ( 
.A1(n_748),
.A2(n_556),
.B(n_524),
.Y(n_940)
);

OA21x2_ASAP7_75t_L g941 ( 
.A1(n_748),
.A2(n_754),
.B(n_749),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_749),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_793),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_754),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_757),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_757),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_758),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_736),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_758),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_804),
.B(n_556),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_824),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_759),
.Y(n_952)
);

BUFx12f_ASAP7_75t_L g953 ( 
.A(n_764),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_759),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_761),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_766),
.Y(n_957)
);

OA21x2_ASAP7_75t_L g958 ( 
.A1(n_766),
.A2(n_631),
.B(n_621),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_773),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_794),
.B(n_621),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_769),
.B(n_448),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_773),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_798),
.B(n_601),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_776),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_776),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_777),
.Y(n_966)
);

OA21x2_ASAP7_75t_L g967 ( 
.A1(n_777),
.A2(n_832),
.B(n_826),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_832),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_858),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_756),
.A2(n_782),
.B1(n_849),
.B2(n_795),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_859),
.B(n_538),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_801),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_802),
.B(n_631),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_859),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_803),
.B(n_674),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_805),
.B(n_674),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_752),
.Y(n_978)
);

OAI22x1_ASAP7_75t_SL g979 ( 
.A1(n_764),
.A2(n_453),
.B1(n_459),
.B2(n_451),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_782),
.A2(n_459),
.B1(n_460),
.B2(n_453),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_857),
.B(n_684),
.Y(n_981)
);

OAI22x1_ASAP7_75t_SL g982 ( 
.A1(n_765),
.A2(n_463),
.B1(n_464),
.B2(n_460),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_769),
.B(n_684),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_795),
.A2(n_464),
.B1(n_467),
.B2(n_463),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_469),
.B1(n_470),
.B2(n_467),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_846),
.Y(n_986)
);

OA21x2_ASAP7_75t_L g987 ( 
.A1(n_846),
.A2(n_692),
.B(n_685),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_820),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_968),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_967),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_925),
.B(n_771),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_967),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_874),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_967),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_927),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_925),
.B(n_771),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_925),
.B(n_772),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_967),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_899),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_899),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_914),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_961),
.B(n_789),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_914),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_868),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_915),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_915),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_881),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_968),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_921),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_921),
.Y(n_1011)
);

BUFx8_ASAP7_75t_L g1012 ( 
.A(n_872),
.Y(n_1012)
);

XNOR2xp5_ASAP7_75t_L g1013 ( 
.A(n_867),
.B(n_753),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_950),
.B(n_792),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_930),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_868),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_983),
.B(n_853),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_930),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_938),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_868),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_971),
.B(n_806),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_898),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_938),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_947),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_898),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_902),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_902),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_888),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_981),
.B(n_772),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_888),
.Y(n_1031)
);

AND2x2_ASAP7_75t_SL g1032 ( 
.A(n_981),
.B(n_685),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_947),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_939),
.B(n_765),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_931),
.B(n_865),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_981),
.B(n_779),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_931),
.B(n_865),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_889),
.B(n_643),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_936),
.B(n_850),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_889),
.B(n_692),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_889),
.B(n_420),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_949),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_896),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_896),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_949),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_889),
.B(n_424),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_904),
.B(n_744),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_903),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_952),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_954),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_954),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_968),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_903),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_968),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_868),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_968),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_873),
.A2(n_477),
.B(n_450),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_962),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_492),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_962),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_923),
.B(n_779),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_910),
.B(n_499),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_944),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_948),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_955),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_955),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_927),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_957),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_912),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_903),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_944),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_969),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_975),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_870),
.B(n_781),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_944),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_870),
.B(n_781),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_975),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_957),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_970),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_970),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_944),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_964),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_868),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_871),
.B(n_799),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_964),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_880),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_965),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_965),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_913),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_871),
.B(n_799),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_913),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_880),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_917),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_917),
.B(n_808),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_970),
.Y(n_1097)
);

OA21x2_ASAP7_75t_L g1098 ( 
.A1(n_873),
.A2(n_508),
.B(n_505),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_917),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_878),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_942),
.B(n_808),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_948),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_910),
.B(n_934),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_923),
.B(n_837),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_942),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_883),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_942),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_910),
.B(n_837),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_948),
.B(n_853),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_941),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_934),
.B(n_838),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_907),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_883),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_883),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_872),
.B(n_762),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_907),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_908),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_908),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_850),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_941),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_918),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_890),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_893),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_918),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_922),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_922),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_932),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_963),
.B(n_851),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_878),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_944),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_945),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_963),
.B(n_851),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_932),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_943),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_973),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_943),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_945),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_934),
.B(n_838),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_869),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_878),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_869),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_945),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_877),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_945),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_941),
.B(n_538),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_945),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_973),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_946),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_946),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_877),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_946),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_986),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_980),
.A2(n_528),
.B1(n_603),
.B2(n_527),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_980),
.B(n_839),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_946),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_946),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_956),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_984),
.B(n_839),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_934),
.B(n_514),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_990),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1128),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1110),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1032),
.A2(n_941),
.B1(n_935),
.B2(n_920),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1032),
.B(n_935),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_1014),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1128),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1065),
.B(n_1102),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_SL g1168 ( 
.A(n_1032),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_991),
.B(n_897),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1110),
.A2(n_935),
.B1(n_920),
.B2(n_887),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_996),
.A2(n_924),
.B1(n_879),
.B2(n_984),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1103),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1110),
.A2(n_935),
.B1(n_920),
.B2(n_887),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1035),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1065),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1070),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1122),
.B(n_953),
.Y(n_1177)
);

BUFx4f_ASAP7_75t_L g1178 ( 
.A(n_1103),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1132),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1103),
.B(n_956),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1005),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1132),
.Y(n_1182)
);

BUFx8_ASAP7_75t_SL g1183 ( 
.A(n_1012),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1000),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1091),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_995),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1000),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_990),
.Y(n_1188)
);

AND2x2_ASAP7_75t_SL g1189 ( 
.A(n_1103),
.B(n_1018),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1001),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1001),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1065),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1076),
.B(n_900),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1035),
.B(n_818),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1002),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1145),
.B(n_956),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1120),
.A2(n_920),
.B1(n_940),
.B2(n_887),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_992),
.B(n_909),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_992),
.B(n_911),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_994),
.B(n_999),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_997),
.B(n_926),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1102),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1012),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1037),
.B(n_900),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1012),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_994),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1120),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1102),
.B(n_973),
.Y(n_1208)
);

AND2x6_ASAP7_75t_L g1209 ( 
.A(n_1120),
.B(n_538),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_999),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1093),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1145),
.A2(n_885),
.B(n_895),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1037),
.B(n_929),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1012),
.B(n_953),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1002),
.B(n_956),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1005),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1064),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1145),
.A2(n_940),
.B1(n_958),
.B2(n_887),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1078),
.B(n_929),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1139),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1023),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1023),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1004),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1004),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1139),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1086),
.B(n_842),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1135),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1039),
.B(n_1119),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1039),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1119),
.B(n_1092),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1005),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1010),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1038),
.B(n_987),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1010),
.A2(n_940),
.B1(n_958),
.B2(n_901),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1026),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1034),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1109),
.B(n_842),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1030),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1141),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1147),
.B(n_843),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1011),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1011),
.A2(n_940),
.B1(n_958),
.B2(n_901),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1015),
.B(n_956),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1015),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_993),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1036),
.B(n_959),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1141),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1019),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1096),
.B(n_843),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1143),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1038),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_993),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1143),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1019),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1020),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1150),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1026),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1060),
.B(n_988),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1038),
.B(n_959),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1020),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1005),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1024),
.B(n_959),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1108),
.B(n_847),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1150),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1038),
.B(n_959),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1027),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1024),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1025),
.A2(n_958),
.B1(n_901),
.B2(n_987),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1025),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_L g1272 ( 
.A(n_1095),
.B(n_901),
.Y(n_1272)
);

CKINVDCx6p67_ASAP7_75t_R g1273 ( 
.A(n_1068),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_SL g1274 ( 
.A(n_1123),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1033),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1111),
.B(n_847),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1040),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1027),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1005),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1033),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1101),
.B(n_959),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1073),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1028),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1042),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1073),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1042),
.A2(n_901),
.B1(n_987),
.B2(n_609),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1041),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1138),
.B(n_966),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1028),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1005),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1040),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1060),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1045),
.B(n_966),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1045),
.A2(n_800),
.B1(n_807),
.B2(n_784),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1049),
.A2(n_901),
.B1(n_987),
.B2(n_609),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1049),
.Y(n_1296)
);

NOR2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1123),
.B(n_893),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1060),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1022),
.B(n_939),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1047),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1003),
.B(n_864),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1050),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1040),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1040),
.B(n_966),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1062),
.B(n_864),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1050),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1051),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1051),
.B(n_966),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1052),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1153),
.B(n_780),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1052),
.B(n_966),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1059),
.B(n_905),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1060),
.B(n_988),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1041),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1104),
.B(n_1154),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1158),
.B(n_985),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1059),
.B(n_985),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1061),
.A2(n_827),
.B1(n_714),
.B2(n_480),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1061),
.B(n_905),
.Y(n_1319)
);

AND2x6_ASAP7_75t_L g1320 ( 
.A(n_1063),
.B(n_523),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1041),
.B(n_905),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_L g1322 ( 
.A(n_1063),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1095),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_998),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1041),
.Y(n_1325)
);

INVx4_ASAP7_75t_SL g1326 ( 
.A(n_1063),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1099),
.B(n_1105),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1046),
.B(n_905),
.Y(n_1328)
);

NAND3x1_ASAP7_75t_L g1329 ( 
.A(n_1153),
.B(n_924),
.C(n_879),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1099),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1105),
.Y(n_1331)
);

INVx4_ASAP7_75t_SL g1332 ( 
.A(n_1063),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1107),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1046),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1107),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1046),
.B(n_905),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1088),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1072),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1017),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1072),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1088),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1046),
.B(n_906),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1159),
.B(n_845),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1017),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1159),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1094),
.Y(n_1346)
);

NAND2xp33_ASAP7_75t_L g1347 ( 
.A(n_1156),
.B(n_901),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1159),
.B(n_988),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1115),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1268),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1167),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1231),
.B(n_1159),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1294),
.B(n_933),
.C(n_978),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1228),
.B(n_1112),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1240),
.B(n_1112),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1193),
.B(n_1219),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1316),
.B(n_891),
.C(n_863),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1162),
.B(n_1156),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1268),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1253),
.B(n_1116),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1189),
.A2(n_1142),
.B1(n_1144),
.B2(n_1137),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1220),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1316),
.B(n_1201),
.C(n_1169),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1169),
.B(n_933),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1317),
.A2(n_974),
.B(n_976),
.C(n_960),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1162),
.B(n_1156),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1253),
.B(n_1116),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1184),
.B(n_1117),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1310),
.A2(n_657),
.B1(n_661),
.B2(n_606),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1201),
.B(n_979),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1187),
.B(n_1117),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1220),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1162),
.B(n_1151),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1190),
.B(n_1124),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1191),
.B(n_1124),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1204),
.B(n_978),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1210),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1177),
.B(n_1123),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1226),
.B(n_1213),
.Y(n_1379)
);

NOR3xp33_ASAP7_75t_L g1380 ( 
.A(n_1171),
.B(n_724),
.C(n_422),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1225),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_L g1382 ( 
.A(n_1305),
.B(n_1013),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1242),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1195),
.B(n_1223),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1225),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1317),
.B(n_979),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1189),
.A2(n_1142),
.B1(n_1144),
.B2(n_1137),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_L g1388 ( 
.A(n_1315),
.B(n_977),
.C(n_703),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1168),
.A2(n_1151),
.B1(n_1155),
.B2(n_1146),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1211),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1160),
.A2(n_1206),
.B1(n_1188),
.B2(n_1199),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1241),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1168),
.A2(n_1155),
.B1(n_1157),
.B2(n_1146),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1167),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1241),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1224),
.B(n_1126),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1249),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1283),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1283),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1234),
.B(n_1126),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1207),
.B(n_1157),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1249),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1207),
.B(n_1077),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1186),
.B(n_1013),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1315),
.A2(n_1134),
.B1(n_1136),
.B2(n_1133),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1289),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1211),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1273),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1185),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1289),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1243),
.B(n_1133),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1251),
.B(n_982),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1338),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1252),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1167),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1252),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1227),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_L g1418 ( 
.A(n_1209),
.B(n_597),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1255),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1246),
.B(n_1134),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1338),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1227),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1340),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1340),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1261),
.A2(n_1009),
.B(n_989),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1250),
.B(n_1136),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1343),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1255),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1251),
.B(n_982),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1256),
.B(n_1066),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1210),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1174),
.A2(n_629),
.B1(n_657),
.B2(n_606),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1177),
.B(n_1123),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1175),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1257),
.B(n_1066),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1262),
.B(n_1067),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1210),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1239),
.B(n_1067),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1210),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1258),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1258),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1207),
.B(n_1077),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1266),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1266),
.Y(n_1444)
);

INVxp33_ASAP7_75t_L g1445 ( 
.A(n_1194),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1323),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1160),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1178),
.B(n_1172),
.Y(n_1448)
);

BUFx8_ASAP7_75t_L g1449 ( 
.A(n_1274),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1301),
.B(n_1305),
.C(n_1318),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1188),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1206),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1198),
.A2(n_689),
.B1(n_661),
.B2(n_610),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1164),
.A2(n_689),
.B1(n_611),
.B2(n_616),
.Y(n_1454)
);

NOR3xp33_ASAP7_75t_L g1455 ( 
.A(n_1301),
.B(n_822),
.C(n_821),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1269),
.B(n_1069),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1176),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1271),
.B(n_1069),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1221),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1265),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1330),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1300),
.B(n_1080),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1229),
.B(n_785),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1178),
.B(n_1077),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1331),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1172),
.B(n_1083),
.Y(n_1466)
);

INVx8_ASAP7_75t_L g1467 ( 
.A(n_1320),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1221),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1286),
.B(n_1083),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1298),
.Y(n_1470)
);

NAND2xp33_ASAP7_75t_L g1471 ( 
.A(n_1209),
.B(n_597),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1333),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1221),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1276),
.B(n_1080),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1275),
.B(n_1084),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_SL g1476 ( 
.A(n_1203),
.B(n_447),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1165),
.B(n_1161),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1175),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1175),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1175),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1286),
.B(n_1083),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1280),
.B(n_1084),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1284),
.B(n_1087),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1166),
.B(n_790),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1179),
.Y(n_1485)
);

BUFx8_ASAP7_75t_L g1486 ( 
.A(n_1274),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1222),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1335),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1182),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1203),
.B(n_1118),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1205),
.B(n_447),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1238),
.A2(n_470),
.B1(n_471),
.B2(n_469),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1296),
.B(n_1087),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1165),
.B(n_1089),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1165),
.B(n_1089),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1277),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1177),
.B(n_823),
.Y(n_1497)
);

NOR2xp67_ASAP7_75t_L g1498 ( 
.A(n_1205),
.B(n_1118),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1222),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_L g1500 ( 
.A(n_1209),
.B(n_1163),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1238),
.B(n_428),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1447),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1363),
.B(n_1322),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1480),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1379),
.B(n_1364),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1480),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1409),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1457),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1450),
.B(n_1322),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1457),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1379),
.A2(n_1329),
.B1(n_1292),
.B2(n_1208),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1440),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1480),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_SL g1514 ( 
.A(n_1378),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1447),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1351),
.B(n_1394),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1451),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1417),
.B(n_1314),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1364),
.B(n_1299),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1451),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1452),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1438),
.B(n_1474),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1480),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1351),
.B(n_1163),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1417),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1422),
.B(n_1314),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1500),
.A2(n_1173),
.B(n_1170),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1440),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1452),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1422),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1434),
.B(n_1277),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1391),
.A2(n_1173),
.B1(n_1170),
.B2(n_1295),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1470),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1362),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1372),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1444),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1381),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1438),
.B(n_1302),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1386),
.A2(n_1299),
.B1(n_1307),
.B2(n_1306),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1385),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1434),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1474),
.B(n_1309),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1460),
.A2(n_1329),
.B1(n_1208),
.B2(n_1299),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1392),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1391),
.A2(n_1295),
.B1(n_1200),
.B2(n_1196),
.Y(n_1545)
);

AND2x6_ASAP7_75t_L g1546 ( 
.A(n_1377),
.B(n_1431),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1444),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1354),
.B(n_1230),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1390),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1407),
.B(n_1325),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1352),
.B(n_1233),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1384),
.B(n_1260),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1356),
.B(n_1349),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1459),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1459),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1386),
.A2(n_1291),
.B1(n_1303),
.B2(n_1325),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1383),
.B(n_1376),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1462),
.B(n_1260),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1394),
.B(n_1291),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1469),
.A2(n_1235),
.B(n_1236),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1370),
.A2(n_1212),
.B(n_1334),
.C(n_1196),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1395),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1377),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1350),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1462),
.B(n_1260),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1494),
.B(n_1313),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1397),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1470),
.Y(n_1568)
);

AOI22x1_ASAP7_75t_L g1569 ( 
.A1(n_1425),
.A2(n_1341),
.B1(n_1346),
.B2(n_1337),
.Y(n_1569)
);

NOR2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1404),
.B(n_1214),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1494),
.B(n_1313),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1449),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1467),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1402),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1495),
.B(n_1313),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1495),
.B(n_1348),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1355),
.B(n_1348),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1449),
.Y(n_1578)
);

AO22x2_ASAP7_75t_L g1579 ( 
.A1(n_1357),
.A2(n_867),
.B1(n_1248),
.B2(n_623),
.Y(n_1579)
);

CKINVDCx6p67_ASAP7_75t_R g1580 ( 
.A(n_1378),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1408),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1445),
.B(n_1348),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1463),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1414),
.Y(n_1584)
);

INVx5_ASAP7_75t_L g1585 ( 
.A(n_1467),
.Y(n_1585)
);

AND2x6_ASAP7_75t_SL g1586 ( 
.A(n_1412),
.B(n_1183),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1485),
.A2(n_1370),
.B1(n_1489),
.B2(n_1429),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1446),
.B(n_1208),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1427),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1505),
.B(n_1477),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1522),
.B(n_1388),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1553),
.B(n_1477),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1380),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1553),
.B(n_1445),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1557),
.B(n_1382),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1557),
.B(n_1476),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1412),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1587),
.B(n_1583),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_SL g1600 ( 
.A(n_1539),
.B(n_1297),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1587),
.B(n_1491),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1508),
.B(n_1353),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1510),
.B(n_1429),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1565),
.B(n_1501),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1532),
.B(n_1431),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1538),
.B(n_1454),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1556),
.B(n_1490),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1556),
.B(n_1498),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1582),
.B(n_1415),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1539),
.B(n_1461),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1582),
.B(n_1415),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_SL g1614 ( 
.A(n_1545),
.B(n_1439),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1518),
.B(n_1448),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1526),
.B(n_1472),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1542),
.B(n_1439),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1533),
.B(n_1369),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1551),
.B(n_1454),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1507),
.B(n_1389),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1566),
.B(n_1393),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1570),
.B(n_1469),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1514),
.B(n_1479),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1571),
.B(n_1455),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1575),
.B(n_1334),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1576),
.B(n_1365),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1577),
.B(n_1369),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1533),
.B(n_1368),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1511),
.B(n_1432),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1552),
.B(n_1369),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1589),
.B(n_1432),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1568),
.B(n_1453),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1543),
.B(n_1371),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1550),
.B(n_1345),
.Y(n_1637)
);

NAND2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1550),
.B(n_1345),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1530),
.B(n_1345),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1549),
.B(n_1303),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1549),
.B(n_1492),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1598),
.B(n_1591),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1606),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1602),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1561),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1601),
.A2(n_1624),
.B1(n_1632),
.B2(n_1612),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1592),
.B(n_1588),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1594),
.B(n_1503),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1561),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1624),
.A2(n_1579),
.B1(n_1509),
.B2(n_1503),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1596),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1616),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1614),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1619),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1619),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1633),
.B(n_1502),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1616),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1590),
.B(n_1509),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_L g1663 ( 
.A(n_1636),
.B(n_1573),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1611),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1613),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1631),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1607),
.B(n_1527),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1502),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1616),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1635),
.B(n_1521),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1623),
.B(n_1521),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1627),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1593),
.B(n_1568),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1630),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1630),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1625),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1609),
.B(n_1536),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1603),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1599),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1610),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1626),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1605),
.B(n_1536),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1608),
.B(n_1515),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1595),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1604),
.B(n_1584),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1615),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1637),
.B(n_1534),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1597),
.A2(n_1560),
.B(n_1524),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_SL g1691 ( 
.A(n_1622),
.B(n_1453),
.C(n_1405),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1639),
.B(n_1516),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1650),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1658),
.A2(n_1248),
.B(n_1361),
.Y(n_1694)
);

BUFx12f_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1656),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1658),
.A2(n_1569),
.B(n_885),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1661),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1676),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.B(n_1579),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1666),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1689),
.A2(n_1559),
.B(n_1366),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_SL g1703 ( 
.A1(n_1654),
.A2(n_1387),
.B(n_1430),
.Y(n_1703)
);

CKINVDCx11_ASAP7_75t_R g1704 ( 
.A(n_1655),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1650),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1682),
.A2(n_1579),
.B1(n_1642),
.B2(n_1634),
.Y(n_1706)
);

INVx6_ASAP7_75t_SL g1707 ( 
.A(n_1692),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1645),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1648),
.B(n_1535),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1659),
.A2(n_1524),
.B(n_1559),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1657),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1661),
.B(n_1516),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1659),
.A2(n_1464),
.B(n_1281),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1689),
.A2(n_1654),
.B(n_1680),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1645),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1645),
.B(n_1573),
.Y(n_1718)
);

AO21x2_ASAP7_75t_L g1719 ( 
.A1(n_1674),
.A2(n_1464),
.B(n_1281),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1661),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1661),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1644),
.A2(n_1366),
.B(n_1358),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1656),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1644),
.A2(n_1358),
.B(n_1245),
.Y(n_1724)
);

INVx6_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1656),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1647),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1682),
.B(n_1467),
.Y(n_1728)
);

AOI22x1_ASAP7_75t_L g1729 ( 
.A1(n_1682),
.A2(n_1531),
.B1(n_1540),
.B2(n_1537),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1647),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1691),
.A2(n_1448),
.B(n_1288),
.Y(n_1731)
);

AOI22x1_ASAP7_75t_L g1732 ( 
.A1(n_1675),
.A2(n_1531),
.B1(n_1562),
.B2(n_1544),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1675),
.B(n_1676),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1660),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1685),
.Y(n_1735)
);

AO21x2_ASAP7_75t_L g1736 ( 
.A1(n_1649),
.A2(n_1373),
.B(n_1418),
.Y(n_1736)
);

BUFx4_ASAP7_75t_R g1737 ( 
.A(n_1664),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1678),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1676),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1660),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1669),
.B(n_1640),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1669),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1671),
.A2(n_1264),
.B(n_1215),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1669),
.B(n_1573),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1652),
.A2(n_540),
.B1(n_447),
.B2(n_1580),
.Y(n_1745)
);

INVx6_ASAP7_75t_L g1746 ( 
.A(n_1692),
.Y(n_1746)
);

BUFx5_ASAP7_75t_L g1747 ( 
.A(n_1677),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1660),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1669),
.B(n_1573),
.Y(n_1749)
);

BUFx12f_ASAP7_75t_L g1750 ( 
.A(n_1692),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1653),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1692),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1666),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1676),
.Y(n_1754)
);

NAND2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1680),
.B(n_1585),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1653),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1671),
.A2(n_1667),
.B(n_1668),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1677),
.Y(n_1758)
);

AO21x2_ASAP7_75t_L g1759 ( 
.A1(n_1649),
.A2(n_1373),
.B(n_1471),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1677),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1648),
.B(n_1567),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1643),
.B(n_1578),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1664),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1667),
.A2(n_1288),
.B(n_1481),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1690),
.B(n_1617),
.Y(n_1765)
);

AO21x2_ASAP7_75t_L g1766 ( 
.A1(n_1662),
.A2(n_1367),
.B(n_1360),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1673),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1664),
.Y(n_1768)
);

INVx6_ASAP7_75t_L g1769 ( 
.A(n_1670),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1691),
.A2(n_1618),
.B(n_1375),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1679),
.B(n_1585),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1665),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1670),
.B(n_1665),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1665),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1673),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1668),
.A2(n_1308),
.B(n_1293),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1687),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1651),
.B(n_1574),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1706),
.A2(n_1679),
.B1(n_1687),
.B2(n_1686),
.Y(n_1779)
);

BUFx2_ASAP7_75t_R g1780 ( 
.A(n_1696),
.Y(n_1780)
);

BUFx2_ASAP7_75t_SL g1781 ( 
.A(n_1738),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1704),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1767),
.A2(n_1686),
.B1(n_1433),
.B2(n_1378),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1775),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1700),
.B(n_1670),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1707),
.Y(n_1786)
);

INVx6_ASAP7_75t_L g1787 ( 
.A(n_1754),
.Y(n_1787)
);

BUFx12f_ASAP7_75t_L g1788 ( 
.A(n_1695),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1769),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1695),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1700),
.A2(n_1663),
.B1(n_1672),
.B2(n_1681),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1725),
.A2(n_1672),
.B1(n_1681),
.B2(n_540),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1725),
.A2(n_1672),
.B1(n_540),
.B2(n_634),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1725),
.A2(n_665),
.B1(n_666),
.B2(n_589),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1701),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1769),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1735),
.Y(n_1797)
);

INVx6_ASAP7_75t_L g1798 ( 
.A(n_1754),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1762),
.Y(n_1799)
);

INVx6_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1763),
.Y(n_1801)
);

INVx6_ASAP7_75t_L g1802 ( 
.A(n_1754),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1753),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1725),
.A2(n_669),
.B1(n_706),
.B2(n_672),
.Y(n_1804)
);

AOI22x1_ASAP7_75t_SL g1805 ( 
.A1(n_1751),
.A2(n_479),
.B1(n_481),
.B2(n_471),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1746),
.A2(n_717),
.B1(n_695),
.B2(n_597),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1727),
.Y(n_1807)
);

BUFx4f_ASAP7_75t_SL g1808 ( 
.A(n_1707),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1737),
.A2(n_1684),
.B1(n_481),
.B2(n_679),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1773),
.B(n_1683),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1750),
.A2(n_1433),
.B1(n_1688),
.B2(n_1497),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1707),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1746),
.A2(n_695),
.B1(n_1684),
.B2(n_1497),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1723),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1769),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1746),
.A2(n_695),
.B1(n_1684),
.B2(n_1497),
.Y(n_1816)
);

BUFx2_ASAP7_75t_SL g1817 ( 
.A(n_1726),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1723),
.Y(n_1818)
);

INVx4_ASAP7_75t_L g1819 ( 
.A(n_1754),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1727),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1730),
.Y(n_1821)
);

INVx6_ASAP7_75t_L g1822 ( 
.A(n_1754),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1716),
.A2(n_678),
.B1(n_683),
.B2(n_479),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1763),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1746),
.A2(n_1752),
.B1(n_1741),
.B2(n_1750),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1730),
.Y(n_1827)
);

BUFx8_ASAP7_75t_L g1828 ( 
.A(n_1723),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1777),
.Y(n_1829)
);

OAI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1765),
.A2(n_1433),
.B1(n_1688),
.B2(n_1572),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1712),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1777),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1752),
.A2(n_695),
.B1(n_1320),
.B2(n_1683),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1752),
.A2(n_695),
.B1(n_1320),
.B2(n_1683),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1712),
.Y(n_1835)
);

BUFx4f_ASAP7_75t_SL g1836 ( 
.A(n_1707),
.Y(n_1836)
);

INVx6_ASAP7_75t_L g1837 ( 
.A(n_1723),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1723),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1693),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1723),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1745),
.A2(n_679),
.B1(n_683),
.B2(n_678),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1696),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1752),
.A2(n_695),
.B1(n_1320),
.B2(n_532),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1752),
.A2(n_695),
.B1(n_1320),
.B2(n_569),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1751),
.B(n_1517),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1768),
.Y(n_1846)
);

INVx6_ASAP7_75t_L g1847 ( 
.A(n_1699),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1693),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1772),
.Y(n_1849)
);

BUFx2_ASAP7_75t_SL g1850 ( 
.A(n_1726),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1693),
.Y(n_1851)
);

BUFx12f_ASAP7_75t_L g1852 ( 
.A(n_1744),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1705),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1768),
.Y(n_1854)
);

NAND2x1p5_ASAP7_75t_L g1855 ( 
.A(n_1699),
.B(n_1585),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1696),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1773),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1752),
.A2(n_695),
.B1(n_588),
.B2(n_591),
.Y(n_1858)
);

INVx8_ASAP7_75t_L g1859 ( 
.A(n_1728),
.Y(n_1859)
);

CKINVDCx6p67_ASAP7_75t_R g1860 ( 
.A(n_1728),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1733),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1741),
.A2(n_598),
.B1(n_605),
.B2(n_548),
.Y(n_1862)
);

INVx6_ASAP7_75t_L g1863 ( 
.A(n_1699),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1734),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1699),
.Y(n_1865)
);

INVx6_ASAP7_75t_L g1866 ( 
.A(n_1739),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1734),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1756),
.A2(n_691),
.B1(n_696),
.B2(n_686),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1739),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1705),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1768),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1705),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1756),
.A2(n_691),
.B1(n_696),
.B2(n_686),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1774),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1711),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1778),
.A2(n_1572),
.B1(n_699),
.B2(n_704),
.Y(n_1876)
);

INVx6_ASAP7_75t_L g1877 ( 
.A(n_1739),
.Y(n_1877)
);

BUFx12f_ASAP7_75t_L g1878 ( 
.A(n_1744),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1740),
.B(n_1520),
.Y(n_1879)
);

INVx8_ASAP7_75t_L g1880 ( 
.A(n_1728),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1716),
.A2(n_699),
.B1(n_704),
.B2(n_698),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1741),
.A2(n_618),
.B1(n_619),
.B2(n_608),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1741),
.A2(n_650),
.B1(n_659),
.B2(n_647),
.Y(n_1883)
);

BUFx8_ASAP7_75t_L g1884 ( 
.A(n_1709),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1744),
.Y(n_1885)
);

INVx6_ASAP7_75t_L g1886 ( 
.A(n_1739),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1711),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1711),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1740),
.B(n_675),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1714),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1703),
.A2(n_681),
.B1(n_682),
.B2(n_676),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1703),
.A2(n_697),
.B1(n_716),
.B2(n_694),
.Y(n_1892)
);

INVx6_ASAP7_75t_L g1893 ( 
.A(n_1744),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1709),
.A2(n_1761),
.B1(n_1733),
.B2(n_1748),
.Y(n_1894)
);

INVx6_ASAP7_75t_L g1895 ( 
.A(n_1749),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1774),
.Y(n_1896)
);

INVx6_ASAP7_75t_L g1897 ( 
.A(n_1749),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1774),
.Y(n_1898)
);

BUFx4_ASAP7_75t_SL g1899 ( 
.A(n_1728),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1713),
.A2(n_828),
.B1(n_829),
.B2(n_825),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1733),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1716),
.A2(n_718),
.B1(n_719),
.B2(n_698),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1714),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1748),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1755),
.A2(n_719),
.B1(n_720),
.B2(n_718),
.Y(n_1905)
);

CKINVDCx8_ASAP7_75t_R g1906 ( 
.A(n_1749),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1713),
.A2(n_833),
.B1(n_834),
.B2(n_831),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1749),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1714),
.Y(n_1909)
);

CKINVDCx16_ASAP7_75t_R g1910 ( 
.A(n_1761),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1728),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_SL g1912 ( 
.A1(n_1716),
.A2(n_721),
.B1(n_725),
.B2(n_720),
.Y(n_1912)
);

BUFx2_ASAP7_75t_SL g1913 ( 
.A(n_1772),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1755),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1772),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1772),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1760),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1755),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1758),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1770),
.A2(n_1638),
.B1(n_836),
.B2(n_840),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1758),
.B(n_1529),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1708),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1757),
.B(n_835),
.Y(n_1923)
);

BUFx3_ASAP7_75t_L g1924 ( 
.A(n_1771),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1771),
.Y(n_1925)
);

CKINVDCx11_ASAP7_75t_R g1926 ( 
.A(n_1747),
.Y(n_1926)
);

INVx6_ASAP7_75t_L g1927 ( 
.A(n_1713),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1760),
.A2(n_725),
.B1(n_721),
.B2(n_537),
.Y(n_1928)
);

BUFx10_ASAP7_75t_L g1929 ( 
.A(n_1713),
.Y(n_1929)
);

CKINVDCx6p67_ASAP7_75t_R g1930 ( 
.A(n_1747),
.Y(n_1930)
);

O2A1O1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1905),
.A2(n_1731),
.B(n_1771),
.C(n_1718),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1807),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1837),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1795),
.B(n_1760),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1824),
.A2(n_1729),
.B(n_1736),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1824),
.A2(n_1729),
.B(n_1736),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1814),
.B(n_1842),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1841),
.A2(n_1718),
.B(n_1717),
.C(n_1708),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1820),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1803),
.B(n_1717),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1917),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1917),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1821),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1827),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1818),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1910),
.B(n_1747),
.Y(n_1946)
);

OA21x2_ASAP7_75t_L g1947 ( 
.A1(n_1923),
.A2(n_1757),
.B(n_1776),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1864),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1857),
.B(n_1747),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1881),
.A2(n_1747),
.B1(n_1759),
.B2(n_1736),
.Y(n_1950)
);

AO31x2_ASAP7_75t_L g1951 ( 
.A1(n_1865),
.A2(n_1715),
.A3(n_1719),
.B(n_1732),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1867),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1904),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1881),
.A2(n_1747),
.B1(n_1759),
.B2(n_1766),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1922),
.B(n_1747),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1810),
.B(n_1747),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1785),
.B(n_1747),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1902),
.A2(n_1759),
.B(n_1766),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1801),
.B(n_1698),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1789),
.B(n_1742),
.Y(n_1960)
);

OA21x2_ASAP7_75t_L g1961 ( 
.A1(n_1923),
.A2(n_1776),
.B(n_1722),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1831),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1801),
.Y(n_1963)
);

A2O1A1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1809),
.A2(n_578),
.B(n_617),
.C(n_568),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1902),
.A2(n_1732),
.B(n_1702),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1799),
.B(n_1586),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1825),
.B(n_1764),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1825),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1835),
.B(n_1698),
.Y(n_1969)
);

A2O1A1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1809),
.A2(n_602),
.B(n_627),
.C(n_580),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1839),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1912),
.A2(n_1766),
.B(n_1718),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1848),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1851),
.Y(n_1974)
);

AO21x2_ASAP7_75t_L g1975 ( 
.A1(n_1811),
.A2(n_1783),
.B(n_1830),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1818),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1853),
.Y(n_1977)
);

AO31x2_ASAP7_75t_L g1978 ( 
.A1(n_1865),
.A2(n_1715),
.A3(n_1719),
.B(n_1694),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1894),
.B(n_1698),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1855),
.A2(n_1722),
.B(n_1743),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1912),
.A2(n_1764),
.B(n_1702),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1796),
.B(n_1815),
.Y(n_1982)
);

OAI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1920),
.A2(n_1698),
.B1(n_1721),
.B2(n_1720),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1829),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1823),
.B(n_1720),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1894),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1870),
.B(n_1764),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1872),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1875),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1884),
.A2(n_1721),
.B1(n_1742),
.B2(n_1720),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1832),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1887),
.B(n_1720),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1846),
.Y(n_1993)
);

AO31x2_ASAP7_75t_L g1994 ( 
.A1(n_1869),
.A2(n_1715),
.A3(n_1719),
.B(n_1694),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1784),
.B(n_1721),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1849),
.Y(n_1996)
);

OA21x2_ASAP7_75t_L g1997 ( 
.A1(n_1888),
.A2(n_1903),
.B(n_1890),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1909),
.B(n_1854),
.Y(n_1998)
);

OAI21x1_ASAP7_75t_L g1999 ( 
.A1(n_1855),
.A2(n_1743),
.B(n_1724),
.Y(n_1999)
);

OAI21x1_ASAP7_75t_L g2000 ( 
.A1(n_1845),
.A2(n_1724),
.B(n_1697),
.Y(n_2000)
);

AO31x2_ASAP7_75t_L g2001 ( 
.A1(n_1869),
.A2(n_1694),
.A3(n_1697),
.B(n_860),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1927),
.B(n_1721),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1871),
.Y(n_2003)
);

AO31x2_ASAP7_75t_L g2004 ( 
.A1(n_1779),
.A2(n_1697),
.A3(n_861),
.B(n_862),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1891),
.A2(n_544),
.B1(n_547),
.B2(n_530),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1874),
.B(n_1742),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1841),
.A2(n_552),
.B1(n_557),
.B2(n_551),
.C(n_549),
.Y(n_2007)
);

CKINVDCx20_ASAP7_75t_R g2008 ( 
.A(n_1782),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1892),
.A2(n_1742),
.B(n_848),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1927),
.B(n_1710),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1896),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1818),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1898),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1919),
.A2(n_559),
.B1(n_562),
.B2(n_558),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1859),
.A2(n_1880),
.B(n_1779),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1814),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1901),
.B(n_1710),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1901),
.B(n_1710),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1845),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1859),
.A2(n_1880),
.B(n_1862),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1791),
.A2(n_854),
.B(n_852),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1787),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1787),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1859),
.A2(n_1880),
.B(n_1882),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1790),
.B(n_1797),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1813),
.A2(n_841),
.B1(n_854),
.B2(n_852),
.Y(n_2026)
);

AO31x2_ASAP7_75t_L g2027 ( 
.A1(n_1819),
.A2(n_1697),
.A3(n_1504),
.B(n_1513),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1816),
.A2(n_856),
.B1(n_577),
.B2(n_579),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1915),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1927),
.B(n_856),
.Y(n_2030)
);

AOI21xp33_ASAP7_75t_SL g2031 ( 
.A1(n_1876),
.A2(n_1183),
.B(n_1486),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1781),
.Y(n_2032)
);

AOI21xp33_ASAP7_75t_SL g2033 ( 
.A1(n_1928),
.A2(n_1486),
.B(n_586),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1861),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1921),
.A2(n_1396),
.B(n_1374),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1916),
.B(n_1842),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1883),
.A2(n_590),
.B1(n_593),
.B2(n_576),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1916),
.B(n_1921),
.Y(n_2038)
);

OAI21x1_ASAP7_75t_SL g2039 ( 
.A1(n_1879),
.A2(n_1826),
.B(n_1819),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1788),
.B(n_596),
.Y(n_2040)
);

OAI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_1793),
.A2(n_626),
.B1(n_628),
.B2(n_612),
.C(n_607),
.Y(n_2041)
);

AOI21x1_ASAP7_75t_L g2042 ( 
.A1(n_1868),
.A2(n_894),
.B(n_892),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1787),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1884),
.B(n_630),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1792),
.A2(n_1437),
.B(n_1585),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1798),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1885),
.B(n_0),
.Y(n_2047)
);

INVx6_ASAP7_75t_L g2048 ( 
.A(n_1828),
.Y(n_2048)
);

OA21x2_ASAP7_75t_L g2049 ( 
.A1(n_1879),
.A2(n_641),
.B(n_640),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1798),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1914),
.B(n_1563),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_SL g2052 ( 
.A1(n_1808),
.A2(n_646),
.B1(n_648),
.B2(n_642),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1889),
.A2(n_1411),
.B(n_1400),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1798),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1840),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_1868),
.A2(n_1873),
.B1(n_1928),
.B2(n_668),
.C(n_654),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1837),
.Y(n_2057)
);

CKINVDCx20_ASAP7_75t_R g2058 ( 
.A(n_1895),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1893),
.A2(n_653),
.B1(n_660),
.B2(n_649),
.Y(n_2059)
);

NAND2x1p5_ASAP7_75t_L g2060 ( 
.A(n_1918),
.B(n_1506),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1900),
.A2(n_1267),
.B(n_1261),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1856),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1800),
.Y(n_2063)
);

AO21x2_ASAP7_75t_L g2064 ( 
.A1(n_1873),
.A2(n_1426),
.B(n_1420),
.Y(n_2064)
);

A2O1A1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_1794),
.A2(n_1804),
.B(n_1858),
.C(n_1806),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1800),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1800),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1780),
.A2(n_667),
.B1(n_662),
.B2(n_1564),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1802),
.B(n_1),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1907),
.A2(n_1267),
.B(n_1478),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1908),
.B(n_2),
.Y(n_2071)
);

OA21x2_ASAP7_75t_L g2072 ( 
.A1(n_1786),
.A2(n_894),
.B(n_892),
.Y(n_2072)
);

AOI21x1_ASAP7_75t_L g2073 ( 
.A1(n_1812),
.A2(n_1436),
.B(n_1435),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1893),
.A2(n_1192),
.B1(n_1202),
.B2(n_986),
.Y(n_2074)
);

BUFx8_ASAP7_75t_L g2075 ( 
.A(n_1852),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1833),
.A2(n_1834),
.B(n_1843),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1802),
.Y(n_2077)
);

A2O1A1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_1924),
.A2(n_430),
.B(n_431),
.C(n_428),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1802),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1822),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1822),
.Y(n_2081)
);

AOI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_1805),
.A2(n_433),
.B1(n_435),
.B2(n_431),
.C(n_430),
.Y(n_2082)
);

BUFx3_ASAP7_75t_L g2083 ( 
.A(n_1837),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1822),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1893),
.A2(n_1192),
.B1(n_1202),
.B2(n_986),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1929),
.B(n_1838),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1895),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1929),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1844),
.A2(n_1218),
.B(n_1236),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2016),
.Y(n_2090)
);

AOI22xp33_ASAP7_75t_SL g2091 ( 
.A1(n_2049),
.A2(n_1836),
.B1(n_1911),
.B2(n_1878),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2019),
.B(n_1897),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2034),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1963),
.B(n_1897),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2049),
.A2(n_1975),
.B1(n_1935),
.B2(n_1936),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1958),
.A2(n_1925),
.B(n_1911),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1937),
.Y(n_2097)
);

AOI222xp33_ASAP7_75t_L g2098 ( 
.A1(n_2056),
.A2(n_446),
.B1(n_435),
.B2(n_449),
.C1(n_444),
.C2(n_433),
.Y(n_2098)
);

A2O1A1Ixp33_ASAP7_75t_L g2099 ( 
.A1(n_2056),
.A2(n_1911),
.B(n_446),
.C(n_449),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_2000),
.A2(n_1980),
.B(n_1999),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2007),
.A2(n_1860),
.B1(n_1897),
.B2(n_1926),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_SL g2102 ( 
.A1(n_1975),
.A2(n_1828),
.B1(n_1850),
.B2(n_1817),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1968),
.B(n_1838),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1997),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2007),
.A2(n_454),
.B1(n_456),
.B2(n_444),
.Y(n_2105)
);

NAND4xp25_ASAP7_75t_L g2106 ( 
.A(n_2082),
.B(n_1458),
.C(n_1475),
.D(n_1456),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2041),
.A2(n_456),
.B1(n_457),
.B2(n_454),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1965),
.A2(n_2009),
.B1(n_2041),
.B2(n_1972),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1950),
.A2(n_461),
.B1(n_462),
.B2(n_457),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2082),
.A2(n_462),
.B1(n_468),
.B2(n_461),
.Y(n_2110)
);

A2O1A1Ixp33_ASAP7_75t_L g2111 ( 
.A1(n_2033),
.A2(n_474),
.B(n_573),
.C(n_468),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_2009),
.A2(n_573),
.B1(n_671),
.B2(n_474),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2005),
.A2(n_673),
.B1(n_688),
.B2(n_671),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1997),
.Y(n_2114)
);

AOI221xp5_ASAP7_75t_L g2115 ( 
.A1(n_1964),
.A2(n_693),
.B1(n_700),
.B2(n_688),
.C(n_673),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1996),
.Y(n_2116)
);

NOR2x1_ASAP7_75t_L g2117 ( 
.A(n_2083),
.B(n_1913),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1941),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1932),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1937),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2005),
.A2(n_700),
.B1(n_701),
.B2(n_693),
.Y(n_2121)
);

AOI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_1970),
.A2(n_705),
.B1(n_707),
.B2(n_702),
.C(n_701),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1954),
.A2(n_705),
.B1(n_707),
.B2(n_702),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1939),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1942),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2076),
.A2(n_1930),
.B1(n_1847),
.B2(n_1866),
.Y(n_2126)
);

OAI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_1986),
.A2(n_1906),
.B(n_711),
.C(n_713),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2076),
.A2(n_1847),
.B1(n_1866),
.B2(n_1863),
.Y(n_2128)
);

BUFx4f_ASAP7_75t_SL g2129 ( 
.A(n_2008),
.Y(n_2129)
);

AOI222xp33_ASAP7_75t_L g2130 ( 
.A1(n_2037),
.A2(n_2014),
.B1(n_2068),
.B2(n_2052),
.C1(n_2044),
.C2(n_1965),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2088),
.B(n_1899),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2039),
.A2(n_1847),
.B1(n_1866),
.B2(n_1863),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2068),
.A2(n_713),
.B1(n_715),
.B2(n_711),
.C(n_709),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_2032),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1962),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1990),
.A2(n_1780),
.B1(n_1877),
.B2(n_1863),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2064),
.A2(n_715),
.B1(n_722),
.B2(n_709),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_1955),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2050),
.B(n_1899),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1993),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2058),
.A2(n_1877),
.B1(n_1886),
.B2(n_1563),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2014),
.A2(n_722),
.B1(n_512),
.B2(n_513),
.C(n_504),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2003),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2065),
.A2(n_1877),
.B1(n_1886),
.B2(n_1563),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1956),
.B(n_1886),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2015),
.A2(n_986),
.B1(n_1541),
.B2(n_1483),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_1955),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_2015),
.A2(n_986),
.B1(n_1541),
.B2(n_1493),
.Y(n_2148)
);

BUFx12f_ASAP7_75t_L g2149 ( 
.A(n_2075),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2013),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2064),
.A2(n_1995),
.B1(n_2030),
.B2(n_2045),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2038),
.B(n_2),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1943),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1944),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1983),
.A2(n_1482),
.B1(n_1513),
.B2(n_1504),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2048),
.A2(n_1563),
.B1(n_1564),
.B2(n_1523),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1971),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_1973),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1931),
.A2(n_515),
.B(n_501),
.Y(n_2159)
);

AOI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_1981),
.A2(n_1328),
.B(n_1321),
.Y(n_2160)
);

A2O1A1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_2031),
.A2(n_534),
.B(n_535),
.C(n_533),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1946),
.B(n_3),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1974),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2069),
.A2(n_1555),
.B1(n_1554),
.B2(n_1528),
.Y(n_2164)
);

BUFx2_ASAP7_75t_L g2165 ( 
.A(n_2081),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1957),
.B(n_3),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2063),
.B(n_1506),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2061),
.A2(n_1342),
.B(n_1336),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1977),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_1988),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2040),
.A2(n_554),
.B1(n_561),
.B2(n_553),
.C(n_539),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2038),
.B(n_4),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_2037),
.A2(n_570),
.B1(n_571),
.B2(n_563),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1989),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_2028),
.A2(n_575),
.B1(n_583),
.B2(n_574),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2048),
.A2(n_1523),
.B1(n_1506),
.B2(n_1512),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1949),
.B(n_5),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1945),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_2021),
.A2(n_595),
.B1(n_613),
.B2(n_592),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2029),
.A2(n_1523),
.B1(n_1506),
.B2(n_1547),
.Y(n_2180)
);

NOR4xp25_ASAP7_75t_L g2181 ( 
.A(n_1938),
.B(n_10),
.C(n_6),
.D(n_7),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2011),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1998),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1948),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_L g2185 ( 
.A(n_2017),
.B(n_2018),
.C(n_2069),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1952),
.Y(n_2186)
);

OAI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2059),
.A2(n_620),
.B1(n_635),
.B2(n_615),
.C(n_614),
.Y(n_2187)
);

OAI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2020),
.A2(n_1523),
.B1(n_637),
.B2(n_638),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2002),
.B(n_6),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2021),
.A2(n_644),
.B1(n_651),
.B2(n_636),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2087),
.A2(n_1546),
.B1(n_1419),
.B2(n_1428),
.Y(n_2191)
);

OAI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2024),
.A2(n_2078),
.B1(n_2055),
.B2(n_1979),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2017),
.A2(n_664),
.B1(n_670),
.B2(n_663),
.C(n_652),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_2062),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1998),
.Y(n_2195)
);

INVx4_ASAP7_75t_L g2196 ( 
.A(n_2062),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1982),
.B(n_7),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_1992),
.Y(n_2198)
);

BUFx2_ASAP7_75t_L g2199 ( 
.A(n_2086),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_2067),
.B(n_10),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2077),
.B(n_11),
.Y(n_2201)
);

AOI21xp33_ASAP7_75t_L g2202 ( 
.A1(n_2018),
.A2(n_12),
.B(n_13),
.Y(n_2202)
);

AOI222xp33_ASAP7_75t_L g2203 ( 
.A1(n_2047),
.A2(n_726),
.B1(n_15),
.B2(n_17),
.C1(n_12),
.C2(n_13),
.Y(n_2203)
);

OAI21xp33_ASAP7_75t_L g2204 ( 
.A1(n_1967),
.A2(n_1441),
.B(n_1416),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2062),
.Y(n_2205)
);

OAI33xp33_ASAP7_75t_L g2206 ( 
.A1(n_1967),
.A2(n_1940),
.A3(n_1987),
.B1(n_1953),
.B2(n_1934),
.B3(n_1992),
.Y(n_2206)
);

AOI222xp33_ASAP7_75t_L g2207 ( 
.A1(n_1966),
.A2(n_17),
.B1(n_20),
.B2(n_15),
.C1(n_16),
.C2(n_19),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2075),
.A2(n_1443),
.B1(n_1546),
.B2(n_1312),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2022),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_SL g2210 ( 
.A1(n_2025),
.A2(n_2080),
.B1(n_2084),
.B2(n_2079),
.Y(n_2210)
);

AOI221xp5_ASAP7_75t_L g2211 ( 
.A1(n_2071),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.C(n_23),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2023),
.B(n_24),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_1987),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2010),
.A2(n_1546),
.B1(n_1312),
.B2(n_1094),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2026),
.A2(n_1546),
.B1(n_1319),
.B2(n_1466),
.Y(n_2215)
);

AOI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_1934),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.C(n_29),
.Y(n_2216)
);

INVx4_ASAP7_75t_L g2217 ( 
.A(n_1945),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2074),
.A2(n_1359),
.B1(n_1399),
.B2(n_1398),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_1945),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1940),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2043),
.B(n_25),
.Y(n_2221)
);

AOI221xp5_ASAP7_75t_L g2222 ( 
.A1(n_1984),
.A2(n_35),
.B1(n_30),
.B2(n_31),
.C(n_36),
.Y(n_2222)
);

OAI21x1_ASAP7_75t_L g2223 ( 
.A1(n_2073),
.A2(n_1466),
.B(n_1401),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2085),
.A2(n_1410),
.B1(n_1413),
.B2(n_1406),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2006),
.Y(n_2225)
);

BUFx3_ASAP7_75t_L g2226 ( 
.A(n_2046),
.Y(n_2226)
);

OAI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2042),
.A2(n_40),
.B1(n_36),
.B2(n_38),
.Y(n_2227)
);

AOI21xp33_ASAP7_75t_L g2228 ( 
.A1(n_2051),
.A2(n_41),
.B(n_42),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_1947),
.B(n_1311),
.C(n_886),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1991),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2054),
.A2(n_1546),
.B1(n_1031),
.B2(n_1043),
.Y(n_2231)
);

BUFx2_ASAP7_75t_L g2232 ( 
.A(n_1976),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2006),
.Y(n_2233)
);

AND2x2_ASAP7_75t_SL g2234 ( 
.A(n_2072),
.B(n_41),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2066),
.B(n_1960),
.Y(n_2235)
);

OAI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2053),
.A2(n_1031),
.B(n_1029),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1985),
.B(n_42),
.Y(n_2237)
);

OAI21xp33_ASAP7_75t_L g2238 ( 
.A1(n_2036),
.A2(n_1969),
.B(n_1959),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2070),
.A2(n_1043),
.B1(n_1044),
.B2(n_1029),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2036),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2060),
.A2(n_1423),
.B1(n_1424),
.B2(n_1421),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2060),
.A2(n_1499),
.B1(n_1473),
.B2(n_1487),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1933),
.B(n_43),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2057),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_SL g2245 ( 
.A1(n_2072),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1976),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1976),
.Y(n_2247)
);

AOI22xp33_ASAP7_75t_L g2248 ( 
.A1(n_1947),
.A2(n_1044),
.B1(n_1090),
.B2(n_1152),
.Y(n_2248)
);

OAI222xp33_ASAP7_75t_L g2249 ( 
.A1(n_2089),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C1(n_48),
.C2(n_50),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2104),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2114),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2158),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2129),
.B(n_2012),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_2117),
.B(n_2012),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2158),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2097),
.B(n_2120),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_2100),
.B(n_2012),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2170),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2185),
.B(n_2004),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_2096),
.A2(n_2035),
.B(n_2001),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2199),
.B(n_1978),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2170),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2165),
.B(n_1978),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2233),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2145),
.B(n_1978),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2205),
.B(n_1994),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_2116),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_2116),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2234),
.A2(n_1961),
.B1(n_2089),
.B2(n_2004),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_2149),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2240),
.B(n_2004),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2225),
.B(n_1994),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2198),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2225),
.B(n_1994),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2131),
.B(n_1951),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2198),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2138),
.B(n_2001),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2138),
.B(n_2147),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2217),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_2196),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2157),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2108),
.A2(n_1961),
.B1(n_1090),
.B2(n_1152),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2220),
.B(n_2001),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2147),
.B(n_1951),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2235),
.B(n_2226),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2183),
.B(n_1951),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2169),
.Y(n_2287)
);

CKINVDCx20_ASAP7_75t_R g2288 ( 
.A(n_2129),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2195),
.Y(n_2289)
);

INVx4_ASAP7_75t_SL g2290 ( 
.A(n_2200),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2232),
.B(n_2027),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2238),
.B(n_2027),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2174),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2246),
.B(n_2027),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2213),
.B(n_47),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2119),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2124),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2213),
.B(n_2244),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2153),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2154),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2209),
.B(n_50),
.Y(n_2301)
);

INVxp67_ASAP7_75t_SL g2302 ( 
.A(n_2103),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2163),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2247),
.B(n_51),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2182),
.Y(n_2305)
);

HB1xp67_ASAP7_75t_L g2306 ( 
.A(n_2093),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2135),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_2178),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2140),
.Y(n_2309)
);

NAND2x1p5_ASAP7_75t_L g2310 ( 
.A(n_2234),
.B(n_1403),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2178),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2090),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2118),
.Y(n_2313)
);

BUFx2_ASAP7_75t_L g2314 ( 
.A(n_2196),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2194),
.B(n_51),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2143),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2125),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2150),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2230),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2184),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2102),
.B(n_884),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2092),
.B(n_53),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2186),
.B(n_55),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2178),
.Y(n_2324)
);

NOR2x1p5_ASAP7_75t_L g2325 ( 
.A(n_2106),
.B(n_56),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2095),
.B(n_56),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2178),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2201),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2194),
.B(n_57),
.Y(n_2329)
);

AND2x4_ASAP7_75t_L g2330 ( 
.A(n_2131),
.B(n_58),
.Y(n_2330)
);

BUFx3_ASAP7_75t_L g2331 ( 
.A(n_2134),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_R g2332 ( 
.A(n_2101),
.B(n_60),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2094),
.B(n_60),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2152),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2172),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2167),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2095),
.B(n_61),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2102),
.B(n_61),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2167),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2132),
.B(n_62),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2139),
.B(n_63),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2223),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2139),
.B(n_64),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2219),
.B(n_64),
.Y(n_2344)
);

AO21x2_ASAP7_75t_L g2345 ( 
.A1(n_2108),
.A2(n_1327),
.B(n_1401),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2221),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2126),
.B(n_65),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2151),
.B(n_65),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2217),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2237),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2197),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2166),
.B(n_66),
.Y(n_2352)
);

BUFx3_ASAP7_75t_L g2353 ( 
.A(n_2200),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2177),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2212),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_2212),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2243),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2204),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2189),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2162),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2210),
.Y(n_2361)
);

CKINVDCx20_ASAP7_75t_R g2362 ( 
.A(n_2192),
.Y(n_2362)
);

AND2x2_ASAP7_75t_SL g2363 ( 
.A(n_2181),
.B(n_67),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2144),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2128),
.B(n_2141),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2136),
.B(n_2091),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2229),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2130),
.A2(n_1125),
.B1(n_1127),
.B2(n_1121),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2164),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2180),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_2206),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2137),
.B(n_2091),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_2188),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2101),
.B(n_67),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2155),
.B(n_68),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2164),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2334),
.B(n_2137),
.Y(n_2377)
);

OAI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2361),
.A2(n_2216),
.B1(n_2202),
.B2(n_2159),
.Y(n_2378)
);

AO31x2_ASAP7_75t_L g2379 ( 
.A1(n_2367),
.A2(n_2176),
.A3(n_2156),
.B(n_2242),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2281),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2250),
.Y(n_2381)
);

AO31x2_ASAP7_75t_L g2382 ( 
.A1(n_2367),
.A2(n_2160),
.A3(n_2241),
.B(n_2099),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2267),
.Y(n_2383)
);

INVx1_ASAP7_75t_SL g2384 ( 
.A(n_2288),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_2256),
.B(n_2146),
.Y(n_2385)
);

AOI21xp33_ASAP7_75t_L g2386 ( 
.A1(n_2366),
.A2(n_2207),
.B(n_2203),
.Y(n_2386)
);

AOI221xp5_ASAP7_75t_L g2387 ( 
.A1(n_2371),
.A2(n_2249),
.B1(n_2206),
.B2(n_2211),
.C(n_2110),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2250),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2366),
.A2(n_2112),
.B(n_2123),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_2270),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2281),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2251),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2363),
.A2(n_2112),
.B1(n_2098),
.B2(n_2222),
.Y(n_2393)
);

AOI211xp5_ASAP7_75t_L g2394 ( 
.A1(n_2361),
.A2(n_2227),
.B(n_2228),
.C(n_2127),
.Y(n_2394)
);

INVxp67_ASAP7_75t_SL g2395 ( 
.A(n_2361),
.Y(n_2395)
);

OAI221xp5_ASAP7_75t_L g2396 ( 
.A1(n_2372),
.A2(n_2110),
.B1(n_2105),
.B2(n_2109),
.C(n_2107),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2256),
.B(n_2148),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2251),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2287),
.Y(n_2399)
);

AOI211xp5_ASAP7_75t_L g2400 ( 
.A1(n_2326),
.A2(n_2227),
.B(n_2133),
.C(n_2111),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2363),
.A2(n_2109),
.B1(n_2105),
.B2(n_2107),
.Y(n_2401)
);

AOI22xp33_ASAP7_75t_L g2402 ( 
.A1(n_2363),
.A2(n_2123),
.B1(n_2121),
.B2(n_2113),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2287),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2293),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2293),
.Y(n_2405)
);

HB1xp67_ASAP7_75t_L g2406 ( 
.A(n_2267),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2268),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2362),
.A2(n_2121),
.B1(n_2113),
.B2(n_2173),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2296),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2360),
.B(n_2214),
.Y(n_2410)
);

INVxp67_ASAP7_75t_L g2411 ( 
.A(n_2335),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2360),
.B(n_2302),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2296),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2337),
.A2(n_2193),
.B(n_2245),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2369),
.B(n_2248),
.Y(n_2415)
);

OA21x2_ASAP7_75t_L g2416 ( 
.A1(n_2286),
.A2(n_2236),
.B(n_2190),
.Y(n_2416)
);

OAI21x1_ASAP7_75t_L g2417 ( 
.A1(n_2283),
.A2(n_2168),
.B(n_2179),
.Y(n_2417)
);

OAI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2371),
.A2(n_2245),
.B(n_2173),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2268),
.Y(n_2419)
);

AO21x2_ASAP7_75t_L g2420 ( 
.A1(n_2295),
.A2(n_2161),
.B(n_2171),
.Y(n_2420)
);

NAND4xp25_ASAP7_75t_L g2421 ( 
.A(n_2269),
.B(n_2122),
.C(n_2115),
.D(n_2142),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2297),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2369),
.B(n_2191),
.Y(n_2423)
);

O2A1O1Ixp5_ASAP7_75t_L g2424 ( 
.A1(n_2371),
.A2(n_2224),
.B(n_2218),
.C(n_2179),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2278),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2360),
.B(n_2208),
.Y(n_2426)
);

AOI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_2325),
.A2(n_2175),
.B1(n_2187),
.B2(n_2190),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2325),
.A2(n_2175),
.B1(n_2208),
.B2(n_2215),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2297),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2278),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2374),
.A2(n_2215),
.B1(n_2239),
.B2(n_2231),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2307),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2311),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2376),
.B(n_68),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2307),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2334),
.B(n_69),
.Y(n_2436)
);

BUFx8_ASAP7_75t_L g2437 ( 
.A(n_2270),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2299),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2285),
.B(n_69),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_2290),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2374),
.A2(n_886),
.B1(n_884),
.B2(n_74),
.Y(n_2441)
);

INVxp67_ASAP7_75t_SL g2442 ( 
.A(n_2311),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_2373),
.B(n_884),
.Y(n_2443)
);

AO21x2_ASAP7_75t_L g2444 ( 
.A1(n_2295),
.A2(n_1442),
.B(n_1403),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2350),
.B(n_71),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2285),
.B(n_71),
.Y(n_2446)
);

AOI21xp33_ASAP7_75t_L g2447 ( 
.A1(n_2348),
.A2(n_73),
.B(n_74),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2299),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2312),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2348),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.C(n_78),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2300),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2336),
.B(n_76),
.Y(n_2452)
);

NAND2x1_ASAP7_75t_L g2453 ( 
.A(n_2254),
.B(n_1209),
.Y(n_2453)
);

INVx3_ASAP7_75t_L g2454 ( 
.A(n_2311),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2376),
.B(n_2350),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2300),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2252),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2312),
.Y(n_2458)
);

OAI21x1_ASAP7_75t_L g2459 ( 
.A1(n_2277),
.A2(n_1442),
.B(n_1098),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2252),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2374),
.A2(n_886),
.B1(n_884),
.B2(n_80),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2313),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2336),
.B(n_78),
.Y(n_2463)
);

OAI211xp5_ASAP7_75t_L g2464 ( 
.A1(n_2332),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2313),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2317),
.Y(n_2466)
);

OAI221xp5_ASAP7_75t_L g2467 ( 
.A1(n_2373),
.A2(n_84),
.B1(n_79),
.B2(n_83),
.C(n_86),
.Y(n_2467)
);

AO21x2_ASAP7_75t_L g2468 ( 
.A1(n_2345),
.A2(n_88),
.B(n_89),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_2351),
.B(n_88),
.Y(n_2469)
);

A2O1A1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2374),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_2470)
);

AOI21x1_ASAP7_75t_L g2471 ( 
.A1(n_2280),
.A2(n_1327),
.B(n_1098),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2317),
.Y(n_2472)
);

AO31x2_ASAP7_75t_L g2473 ( 
.A1(n_2280),
.A2(n_94),
.A3(n_92),
.B(n_93),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2277),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_SL g2475 ( 
.A1(n_2330),
.A2(n_97),
.B1(n_94),
.B2(n_95),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2255),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2255),
.Y(n_2477)
);

INVxp67_ASAP7_75t_SL g2478 ( 
.A(n_2311),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2258),
.Y(n_2479)
);

OAI21x1_ASAP7_75t_L g2480 ( 
.A1(n_2271),
.A2(n_1098),
.B(n_1058),
.Y(n_2480)
);

OAI21x1_ASAP7_75t_L g2481 ( 
.A1(n_2284),
.A2(n_1098),
.B(n_1058),
.Y(n_2481)
);

AOI21xp33_ASAP7_75t_L g2482 ( 
.A1(n_2345),
.A2(n_95),
.B(n_98),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2353),
.B(n_98),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2365),
.B(n_99),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2258),
.Y(n_2485)
);

OAI21xp33_ASAP7_75t_L g2486 ( 
.A1(n_2282),
.A2(n_100),
.B(n_101),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2262),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2365),
.B(n_100),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2321),
.A2(n_1180),
.B(n_102),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2390),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2440),
.B(n_2314),
.Y(n_2491)
);

AND2x4_ASAP7_75t_L g2492 ( 
.A(n_2383),
.B(n_2290),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2377),
.B(n_2357),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2383),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_2390),
.Y(n_2495)
);

AOI211x1_ASAP7_75t_L g2496 ( 
.A1(n_2418),
.A2(n_2386),
.B(n_2389),
.C(n_2464),
.Y(n_2496)
);

INVxp67_ASAP7_75t_L g2497 ( 
.A(n_2395),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2406),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2406),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2412),
.B(n_2425),
.Y(n_2500)
);

INVx1_ASAP7_75t_SL g2501 ( 
.A(n_2384),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2380),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2437),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2391),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2407),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2425),
.B(n_2314),
.Y(n_2506)
);

AND2x4_ASAP7_75t_SL g2507 ( 
.A(n_2439),
.B(n_2330),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2484),
.B(n_2357),
.Y(n_2508)
);

NAND3xp33_ASAP7_75t_SL g2509 ( 
.A(n_2387),
.B(n_2338),
.C(n_2347),
.Y(n_2509)
);

OAI33xp33_ASAP7_75t_L g2510 ( 
.A1(n_2411),
.A2(n_2259),
.A3(n_2262),
.B1(n_2276),
.B2(n_2273),
.B3(n_2358),
.Y(n_2510)
);

INVx2_ASAP7_75t_SL g2511 ( 
.A(n_2437),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2433),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2430),
.B(n_2275),
.Y(n_2513)
);

HB1xp67_ASAP7_75t_L g2514 ( 
.A(n_2407),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2437),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2433),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2455),
.B(n_2430),
.Y(n_2517)
);

OAI221xp5_ASAP7_75t_L g2518 ( 
.A1(n_2394),
.A2(n_2338),
.B1(n_2364),
.B2(n_2358),
.C(n_2259),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2419),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2433),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2454),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2426),
.B(n_2275),
.Y(n_2522)
);

OAI211xp5_ASAP7_75t_L g2523 ( 
.A1(n_2393),
.A2(n_2347),
.B(n_2340),
.C(n_2375),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2442),
.B(n_2275),
.Y(n_2524)
);

OAI211xp5_ASAP7_75t_L g2525 ( 
.A1(n_2393),
.A2(n_2340),
.B(n_2375),
.C(n_2364),
.Y(n_2525)
);

INVx2_ASAP7_75t_SL g2526 ( 
.A(n_2419),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_L g2527 ( 
.A1(n_2401),
.A2(n_2345),
.B1(n_2330),
.B2(n_2351),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2399),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2403),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2454),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2488),
.B(n_2328),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2378),
.A2(n_2401),
.B1(n_2402),
.B2(n_2421),
.Y(n_2532)
);

NAND3xp33_ASAP7_75t_L g2533 ( 
.A(n_2424),
.B(n_2368),
.C(n_2342),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2381),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2478),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2410),
.B(n_2279),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2446),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2385),
.B(n_2279),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_2381),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2404),
.Y(n_2540)
);

INVx3_ASAP7_75t_L g2541 ( 
.A(n_2388),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2388),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2392),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2405),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2397),
.B(n_2279),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2449),
.B(n_2339),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2474),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2434),
.B(n_2423),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2449),
.B(n_2339),
.Y(n_2549)
);

OAI221xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2402),
.A2(n_2343),
.B1(n_2341),
.B2(n_2292),
.C(n_2356),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2392),
.Y(n_2551)
);

AOI221xp5_ASAP7_75t_L g2552 ( 
.A1(n_2378),
.A2(n_2354),
.B1(n_2322),
.B2(n_2333),
.C(n_2330),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2398),
.Y(n_2553)
);

AOI221xp5_ASAP7_75t_L g2554 ( 
.A1(n_2414),
.A2(n_2354),
.B1(n_2333),
.B2(n_2346),
.C(n_2328),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2474),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_2473),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2398),
.Y(n_2557)
);

AOI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2447),
.A2(n_2346),
.B1(n_2356),
.B2(n_2276),
.C(n_2273),
.Y(n_2558)
);

AOI222xp33_ASAP7_75t_L g2559 ( 
.A1(n_2396),
.A2(n_2352),
.B1(n_2343),
.B2(n_2341),
.C1(n_2355),
.C2(n_2290),
.Y(n_2559)
);

INVxp67_ASAP7_75t_L g2560 ( 
.A(n_2443),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2452),
.B(n_2359),
.Y(n_2561)
);

BUFx2_ASAP7_75t_L g2562 ( 
.A(n_2473),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2458),
.B(n_2265),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2458),
.B(n_2265),
.Y(n_2564)
);

CKINVDCx20_ASAP7_75t_R g2565 ( 
.A(n_2475),
.Y(n_2565)
);

AND2x4_ASAP7_75t_SL g2566 ( 
.A(n_2463),
.B(n_2254),
.Y(n_2566)
);

BUFx2_ASAP7_75t_L g2567 ( 
.A(n_2473),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2409),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2432),
.B(n_2264),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2432),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2413),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_SL g2572 ( 
.A1(n_2408),
.A2(n_2331),
.B1(n_2253),
.B2(n_2353),
.Y(n_2572)
);

AO21x2_ASAP7_75t_L g2573 ( 
.A1(n_2482),
.A2(n_2468),
.B(n_2417),
.Y(n_2573)
);

OR2x2_ASAP7_75t_L g2574 ( 
.A(n_2435),
.B(n_2264),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2462),
.B(n_2298),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2422),
.B(n_2290),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2483),
.Y(n_2577)
);

INVx2_ASAP7_75t_SL g2578 ( 
.A(n_2492),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2491),
.B(n_2417),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2491),
.B(n_2379),
.Y(n_2580)
);

AND2x4_ASAP7_75t_L g2581 ( 
.A(n_2492),
.B(n_2457),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2497),
.B(n_2443),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2496),
.B(n_2532),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2547),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2501),
.B(n_2483),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2515),
.B(n_2331),
.Y(n_2586)
);

NAND2x1p5_ASAP7_75t_L g2587 ( 
.A(n_2535),
.B(n_2323),
.Y(n_2587)
);

OR2x2_ASAP7_75t_L g2588 ( 
.A(n_2548),
.B(n_2415),
.Y(n_2588)
);

AND2x4_ASAP7_75t_SL g2589 ( 
.A(n_2492),
.B(n_2495),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2495),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2538),
.B(n_2379),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2495),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2555),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2537),
.B(n_2436),
.Y(n_2594)
);

AND2x4_ASAP7_75t_SL g2595 ( 
.A(n_2495),
.B(n_2254),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2535),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2538),
.B(n_2349),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2493),
.B(n_2469),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2495),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2545),
.B(n_2379),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2490),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2545),
.B(n_2379),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2494),
.Y(n_2603)
);

BUFx2_ASAP7_75t_L g2604 ( 
.A(n_2490),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2536),
.B(n_2324),
.Y(n_2605)
);

INVx1_ASAP7_75t_SL g2606 ( 
.A(n_2503),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2505),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2536),
.B(n_2522),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2490),
.B(n_2460),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2522),
.B(n_2324),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2503),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2537),
.B(n_2445),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2566),
.B(n_2349),
.Y(n_2613)
);

NAND4xp25_ASAP7_75t_L g2614 ( 
.A(n_2559),
.B(n_2408),
.C(n_2427),
.D(n_2400),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2526),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2498),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2554),
.B(n_2420),
.Y(n_2617)
);

INVxp67_ASAP7_75t_L g2618 ( 
.A(n_2572),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2552),
.B(n_2420),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2531),
.B(n_2508),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2499),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2517),
.B(n_2476),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2566),
.B(n_2355),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2517),
.B(n_2477),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2514),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2524),
.B(n_2327),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2576),
.B(n_2479),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2525),
.B(n_2359),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2526),
.Y(n_2629)
);

NOR2xp67_ASAP7_75t_L g2630 ( 
.A(n_2515),
.B(n_2485),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2519),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_2515),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2528),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2528),
.Y(n_2634)
);

INVx1_ASAP7_75t_SL g2635 ( 
.A(n_2577),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2502),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2550),
.B(n_2487),
.Y(n_2637)
);

BUFx2_ASAP7_75t_SL g2638 ( 
.A(n_2511),
.Y(n_2638)
);

OR2x2_ASAP7_75t_L g2639 ( 
.A(n_2561),
.B(n_2429),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2504),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2539),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2524),
.B(n_2327),
.Y(n_2642)
);

INVxp67_ASAP7_75t_L g2643 ( 
.A(n_2577),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2506),
.B(n_2435),
.Y(n_2644)
);

OR2x2_ASAP7_75t_L g2645 ( 
.A(n_2533),
.B(n_2438),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2506),
.B(n_2462),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2539),
.Y(n_2647)
);

NAND2x1_ASAP7_75t_L g2648 ( 
.A(n_2576),
.B(n_2254),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2500),
.B(n_2465),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2576),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2539),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2541),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2541),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2529),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2556),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2560),
.B(n_2315),
.Y(n_2656)
);

OR2x2_ASAP7_75t_L g2657 ( 
.A(n_2509),
.B(n_2448),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2523),
.B(n_2315),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2500),
.B(n_2451),
.Y(n_2659)
);

BUFx3_ASAP7_75t_L g2660 ( 
.A(n_2611),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2638),
.B(n_2511),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2589),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2635),
.B(n_2565),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2589),
.B(n_2507),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2619),
.A2(n_2565),
.B1(n_2518),
.B2(n_2510),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2607),
.Y(n_2666)
);

NOR4xp25_ASAP7_75t_L g2667 ( 
.A(n_2583),
.B(n_2467),
.C(n_2450),
.D(n_2470),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2607),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2655),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2608),
.B(n_2507),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_2655),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2608),
.B(n_2575),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2606),
.B(n_2575),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2587),
.Y(n_2674)
);

NOR2x1_ASAP7_75t_L g2675 ( 
.A(n_2604),
.B(n_2556),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2596),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2650),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2584),
.B(n_2593),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2615),
.Y(n_2679)
);

NAND4xp75_ASAP7_75t_SL g2680 ( 
.A(n_2586),
.B(n_2416),
.C(n_2549),
.D(n_2546),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2587),
.Y(n_2681)
);

INVx1_ASAP7_75t_SL g2682 ( 
.A(n_2611),
.Y(n_2682)
);

NAND4xp75_ASAP7_75t_SL g2683 ( 
.A(n_2586),
.B(n_2416),
.C(n_2549),
.D(n_2546),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2615),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2629),
.Y(n_2685)
);

XNOR2xp5_ASAP7_75t_L g2686 ( 
.A(n_2614),
.B(n_2427),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2629),
.Y(n_2687)
);

OA22x2_ASAP7_75t_L g2688 ( 
.A1(n_2617),
.A2(n_2567),
.B1(n_2562),
.B2(n_2530),
.Y(n_2688)
);

OR2x2_ASAP7_75t_L g2689 ( 
.A(n_2658),
.B(n_2527),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2633),
.Y(n_2690)
);

INVxp67_ASAP7_75t_L g2691 ( 
.A(n_2585),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2623),
.B(n_2521),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2618),
.A2(n_2632),
.B1(n_2643),
.B2(n_2573),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2634),
.Y(n_2694)
);

XOR2x2_ASAP7_75t_L g2695 ( 
.A(n_2657),
.B(n_2558),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2613),
.B(n_2521),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2650),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2610),
.B(n_2530),
.Y(n_2698)
);

NAND4xp75_ASAP7_75t_L g2699 ( 
.A(n_2630),
.B(n_2489),
.C(n_2516),
.D(n_2512),
.Y(n_2699)
);

INVxp67_ASAP7_75t_SL g2700 ( 
.A(n_2590),
.Y(n_2700)
);

NOR3xp33_ASAP7_75t_L g2701 ( 
.A(n_2601),
.B(n_2470),
.C(n_2562),
.Y(n_2701)
);

NAND4xp75_ASAP7_75t_SL g2702 ( 
.A(n_2579),
.B(n_2416),
.C(n_2329),
.D(n_2513),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2637),
.A2(n_2567),
.B1(n_2645),
.B2(n_2428),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2625),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2610),
.B(n_2597),
.Y(n_2705)
);

NAND4xp75_ASAP7_75t_L g2706 ( 
.A(n_2578),
.B(n_2516),
.C(n_2520),
.D(n_2512),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2631),
.B(n_2540),
.Y(n_2707)
);

INVx2_ASAP7_75t_SL g2708 ( 
.A(n_2595),
.Y(n_2708)
);

NAND3xp33_ASAP7_75t_L g2709 ( 
.A(n_2628),
.B(n_2461),
.C(n_2441),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2605),
.B(n_2513),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2588),
.B(n_2573),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2659),
.Y(n_2712)
);

NOR3xp33_ASAP7_75t_L g2713 ( 
.A(n_2601),
.B(n_2486),
.C(n_2520),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2648),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2622),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2590),
.B(n_2544),
.Y(n_2716)
);

NAND4xp75_ASAP7_75t_L g2717 ( 
.A(n_2578),
.B(n_2329),
.C(n_2344),
.D(n_2534),
.Y(n_2717)
);

AO22x2_ASAP7_75t_L g2718 ( 
.A1(n_2603),
.A2(n_2571),
.B1(n_2568),
.B2(n_2534),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2605),
.B(n_2563),
.Y(n_2719)
);

NOR2x1_ASAP7_75t_L g2720 ( 
.A(n_2592),
.B(n_2573),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2624),
.Y(n_2721)
);

OAI21xp33_ASAP7_75t_SL g2722 ( 
.A1(n_2680),
.A2(n_2579),
.B(n_2591),
.Y(n_2722)
);

NOR4xp25_ASAP7_75t_L g2723 ( 
.A(n_2703),
.B(n_2592),
.C(n_2599),
.D(n_2616),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2661),
.B(n_2595),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2671),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2667),
.B(n_2599),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2682),
.B(n_2598),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2671),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2668),
.Y(n_2729)
);

OR2x2_ASAP7_75t_L g2730 ( 
.A(n_2678),
.B(n_2594),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2686),
.B(n_2621),
.Y(n_2731)
);

A2O1A1Ixp33_ASAP7_75t_L g2732 ( 
.A1(n_2665),
.A2(n_2582),
.B(n_2580),
.C(n_2591),
.Y(n_2732)
);

AOI32xp33_ASAP7_75t_L g2733 ( 
.A1(n_2703),
.A2(n_2580),
.A3(n_2600),
.B1(n_2602),
.B2(n_2650),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2697),
.Y(n_2734)
);

INVxp33_ASAP7_75t_L g2735 ( 
.A(n_2663),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2700),
.B(n_2636),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_2674),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2660),
.B(n_2612),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2673),
.B(n_2609),
.Y(n_2739)
);

A2O1A1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2709),
.A2(n_2602),
.B(n_2600),
.C(n_2656),
.Y(n_2740)
);

AOI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2695),
.A2(n_2609),
.B(n_2581),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_2664),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2678),
.B(n_2620),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2714),
.Y(n_2744)
);

INVxp67_ASAP7_75t_SL g2745 ( 
.A(n_2714),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2679),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2670),
.B(n_2626),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2700),
.B(n_2679),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2718),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2718),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2664),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2677),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2718),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2669),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2666),
.Y(n_2755)
);

OR2x6_ASAP7_75t_L g2756 ( 
.A(n_2662),
.B(n_2708),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2675),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2684),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2685),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2691),
.B(n_2639),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2687),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2691),
.B(n_2649),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2710),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2701),
.B(n_2640),
.Y(n_2764)
);

NAND2x1_ASAP7_75t_L g2765 ( 
.A(n_2681),
.B(n_2609),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2701),
.B(n_2654),
.Y(n_2766)
);

INVx3_ASAP7_75t_SL g2767 ( 
.A(n_2692),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2705),
.B(n_2626),
.Y(n_2768)
);

OAI21xp33_ASAP7_75t_L g2769 ( 
.A1(n_2732),
.A2(n_2689),
.B(n_2693),
.Y(n_2769)
);

AOI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2742),
.A2(n_2717),
.B1(n_2672),
.B2(n_2688),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2746),
.Y(n_2771)
);

OAI21xp33_ASAP7_75t_L g2772 ( 
.A1(n_2735),
.A2(n_2723),
.B(n_2726),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2748),
.Y(n_2773)
);

OAI22xp33_ASAP7_75t_SL g2774 ( 
.A1(n_2749),
.A2(n_2711),
.B1(n_2720),
.B2(n_2715),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2726),
.A2(n_2688),
.B1(n_2699),
.B2(n_2696),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2722),
.A2(n_2713),
.B1(n_2698),
.B2(n_2706),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2723),
.A2(n_2707),
.B(n_2721),
.Y(n_2777)
);

OAI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2731),
.A2(n_2712),
.B1(n_2676),
.B2(n_2704),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2748),
.Y(n_2779)
);

OAI21xp33_ASAP7_75t_L g2780 ( 
.A1(n_2751),
.A2(n_2719),
.B(n_2713),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2725),
.Y(n_2781)
);

OAI21xp33_ASAP7_75t_SL g2782 ( 
.A1(n_2733),
.A2(n_2683),
.B(n_2680),
.Y(n_2782)
);

OAI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2741),
.A2(n_2707),
.B(n_2716),
.Y(n_2783)
);

AOI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2724),
.A2(n_2642),
.B1(n_2581),
.B2(n_2627),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_2767),
.B(n_2716),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2756),
.A2(n_2642),
.B1(n_2581),
.B2(n_2627),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2756),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2731),
.A2(n_2428),
.B1(n_2627),
.B2(n_2461),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2756),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2765),
.Y(n_2790)
);

OAI21xp33_ASAP7_75t_L g2791 ( 
.A1(n_2738),
.A2(n_2649),
.B(n_2646),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2728),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2727),
.B(n_2644),
.Y(n_2793)
);

AOI22xp33_ASAP7_75t_SL g2794 ( 
.A1(n_2757),
.A2(n_2683),
.B1(n_2702),
.B2(n_2646),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2747),
.A2(n_2644),
.B1(n_2468),
.B2(n_2690),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2768),
.B(n_2694),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2740),
.A2(n_2441),
.B1(n_2647),
.B2(n_2641),
.Y(n_2797)
);

INVx1_ASAP7_75t_SL g2798 ( 
.A(n_2762),
.Y(n_2798)
);

OAI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2764),
.A2(n_2702),
.B(n_2647),
.Y(n_2799)
);

AOI211xp5_ASAP7_75t_L g2800 ( 
.A1(n_2764),
.A2(n_2352),
.B(n_2323),
.C(n_2641),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2744),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2737),
.A2(n_2763),
.B1(n_2745),
.B2(n_2734),
.Y(n_2802)
);

AOI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2739),
.A2(n_2651),
.B1(n_2653),
.B2(n_2652),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2766),
.A2(n_2651),
.B1(n_2653),
.B2(n_2652),
.Y(n_2804)
);

OAI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2766),
.A2(n_2551),
.B(n_2543),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2729),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2771),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2772),
.B(n_2730),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2787),
.B(n_2752),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2789),
.B(n_2743),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2790),
.Y(n_2811)
);

OAI21xp5_ASAP7_75t_SL g2812 ( 
.A1(n_2776),
.A2(n_2753),
.B(n_2750),
.Y(n_2812)
);

INVx1_ASAP7_75t_SL g2813 ( 
.A(n_2798),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2796),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2802),
.Y(n_2815)
);

OAI21xp33_ASAP7_75t_L g2816 ( 
.A1(n_2769),
.A2(n_2755),
.B(n_2754),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2777),
.A2(n_2774),
.B(n_2783),
.Y(n_2817)
);

AOI211x1_ASAP7_75t_SL g2818 ( 
.A1(n_2797),
.A2(n_2736),
.B(n_2551),
.C(n_2557),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2793),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2780),
.B(n_2758),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2798),
.B(n_2761),
.Y(n_2821)
);

XNOR2xp5_ASAP7_75t_L g2822 ( 
.A(n_2784),
.B(n_2760),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2773),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2775),
.A2(n_2788),
.B1(n_2782),
.B2(n_2791),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2801),
.B(n_2806),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2770),
.B(n_2736),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2779),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2781),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2794),
.A2(n_2759),
.B1(n_2344),
.B2(n_2304),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2792),
.Y(n_2830)
);

AOI31xp33_ASAP7_75t_L g2831 ( 
.A1(n_2785),
.A2(n_2304),
.A3(n_2557),
.B(n_2543),
.Y(n_2831)
);

OAI21x1_ASAP7_75t_SL g2832 ( 
.A1(n_2786),
.A2(n_2570),
.B(n_2308),
.Y(n_2832)
);

OAI32xp33_ASAP7_75t_L g2833 ( 
.A1(n_2799),
.A2(n_2541),
.A3(n_2553),
.B1(n_2542),
.B2(n_2570),
.Y(n_2833)
);

OA22x2_ASAP7_75t_L g2834 ( 
.A1(n_2803),
.A2(n_2553),
.B1(n_2542),
.B2(n_2563),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2805),
.Y(n_2835)
);

OAI22x1_ASAP7_75t_L g2836 ( 
.A1(n_2795),
.A2(n_2308),
.B1(n_2553),
.B2(n_2542),
.Y(n_2836)
);

OA222x2_ASAP7_75t_L g2837 ( 
.A1(n_2778),
.A2(n_2473),
.B1(n_2574),
.B2(n_2569),
.C1(n_2456),
.C2(n_2472),
.Y(n_2837)
);

AOI22xp33_ASAP7_75t_L g2838 ( 
.A1(n_2804),
.A2(n_2444),
.B1(n_2564),
.B2(n_2431),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2817),
.A2(n_2800),
.B(n_2574),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2826),
.A2(n_2800),
.B1(n_2569),
.B2(n_2564),
.Y(n_2840)
);

AOI31xp33_ASAP7_75t_L g2841 ( 
.A1(n_2813),
.A2(n_2808),
.A3(n_2811),
.B(n_2821),
.Y(n_2841)
);

NAND3xp33_ASAP7_75t_SL g2842 ( 
.A(n_2818),
.B(n_2301),
.C(n_2453),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2810),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2812),
.A2(n_2370),
.B1(n_2311),
.B2(n_2444),
.Y(n_2844)
);

INVxp33_ASAP7_75t_L g2845 ( 
.A(n_2822),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2814),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2829),
.B(n_2465),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2829),
.B(n_2466),
.Y(n_2848)
);

INVx2_ASAP7_75t_SL g2849 ( 
.A(n_2825),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2819),
.B(n_2466),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2809),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2834),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2815),
.A2(n_2370),
.B1(n_2301),
.B2(n_2257),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2824),
.B(n_2472),
.Y(n_2854)
);

NAND2xp67_ASAP7_75t_L g2855 ( 
.A(n_2820),
.B(n_2266),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2832),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2816),
.A2(n_2257),
.B(n_2431),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2807),
.Y(n_2858)
);

OAI21xp33_ASAP7_75t_L g2859 ( 
.A1(n_2831),
.A2(n_2257),
.B(n_2342),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2835),
.B(n_2828),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2830),
.Y(n_2861)
);

OAI322xp33_ASAP7_75t_L g2862 ( 
.A1(n_2823),
.A2(n_2284),
.A3(n_2274),
.B1(n_2272),
.B2(n_2310),
.C1(n_2263),
.C2(n_2266),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2827),
.B(n_2261),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2843),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2841),
.A2(n_2833),
.B(n_2836),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_2845),
.B(n_2838),
.Y(n_2866)
);

BUFx2_ASAP7_75t_L g2867 ( 
.A(n_2849),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2841),
.A2(n_2837),
.B(n_2257),
.Y(n_2868)
);

NOR2x1_ASAP7_75t_L g2869 ( 
.A(n_2856),
.B(n_2837),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2846),
.Y(n_2870)
);

AOI21xp33_ASAP7_75t_L g2871 ( 
.A1(n_2851),
.A2(n_102),
.B(n_103),
.Y(n_2871)
);

AOI211xp5_ASAP7_75t_L g2872 ( 
.A1(n_2839),
.A2(n_2261),
.B(n_2263),
.C(n_2291),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2847),
.Y(n_2873)
);

NOR2x1_ASAP7_75t_SL g2874 ( 
.A(n_2840),
.B(n_2298),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2854),
.B(n_2306),
.Y(n_2875)
);

OR2x2_ASAP7_75t_L g2876 ( 
.A(n_2852),
.B(n_2319),
.Y(n_2876)
);

INVxp67_ASAP7_75t_SL g2877 ( 
.A(n_2848),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2857),
.B(n_2272),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2860),
.Y(n_2879)
);

AOI211xp5_ASAP7_75t_L g2880 ( 
.A1(n_2842),
.A2(n_2291),
.B(n_2274),
.C(n_2459),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2858),
.B(n_2289),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2855),
.B(n_2289),
.Y(n_2882)
);

AOI221xp5_ASAP7_75t_L g2883 ( 
.A1(n_2865),
.A2(n_2861),
.B1(n_2863),
.B2(n_2850),
.C(n_2859),
.Y(n_2883)
);

AOI221xp5_ASAP7_75t_L g2884 ( 
.A1(n_2868),
.A2(n_2862),
.B1(n_2844),
.B2(n_2853),
.C(n_2294),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2867),
.B(n_2382),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2864),
.B(n_2382),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_SL g2887 ( 
.A(n_2879),
.B(n_2862),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2866),
.B(n_2382),
.Y(n_2888)
);

NOR3xp33_ASAP7_75t_L g2889 ( 
.A(n_2877),
.B(n_2459),
.C(n_2480),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2874),
.B(n_2382),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2870),
.B(n_2305),
.Y(n_2891)
);

NAND4xp25_ASAP7_75t_L g2892 ( 
.A(n_2876),
.B(n_2294),
.C(n_2316),
.D(n_2309),
.Y(n_2892)
);

OAI211xp5_ASAP7_75t_L g2893 ( 
.A1(n_2869),
.A2(n_107),
.B(n_104),
.C(n_106),
.Y(n_2893)
);

NOR2x1_ASAP7_75t_L g2894 ( 
.A(n_2873),
.B(n_104),
.Y(n_2894)
);

OAI21xp33_ASAP7_75t_L g2895 ( 
.A1(n_2875),
.A2(n_2310),
.B(n_2471),
.Y(n_2895)
);

INVx2_ASAP7_75t_SL g2896 ( 
.A(n_2894),
.Y(n_2896)
);

OAI22xp33_ASAP7_75t_SL g2897 ( 
.A1(n_2887),
.A2(n_2878),
.B1(n_2882),
.B2(n_2881),
.Y(n_2897)
);

A2O1A1Ixp33_ASAP7_75t_SL g2898 ( 
.A1(n_2893),
.A2(n_2872),
.B(n_2885),
.C(n_2871),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2886),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2891),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2890),
.Y(n_2901)
);

BUFx2_ASAP7_75t_L g2902 ( 
.A(n_2883),
.Y(n_2902)
);

AOI221xp5_ASAP7_75t_L g2903 ( 
.A1(n_2884),
.A2(n_2871),
.B1(n_2880),
.B2(n_2316),
.C(n_2318),
.Y(n_2903)
);

OAI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2888),
.A2(n_2320),
.B1(n_2309),
.B2(n_2318),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2892),
.Y(n_2905)
);

O2A1O1Ixp33_ASAP7_75t_L g2906 ( 
.A1(n_2895),
.A2(n_2310),
.B(n_109),
.C(n_107),
.Y(n_2906)
);

AOI221xp5_ASAP7_75t_L g2907 ( 
.A1(n_2889),
.A2(n_2303),
.B1(n_2305),
.B2(n_2320),
.C(n_111),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2887),
.A2(n_2260),
.B1(n_2303),
.B2(n_2480),
.Y(n_2908)
);

AOI221x1_ASAP7_75t_L g2909 ( 
.A1(n_2897),
.A2(n_2901),
.B1(n_2899),
.B2(n_2900),
.C(n_2905),
.Y(n_2909)
);

AOI221xp5_ASAP7_75t_L g2910 ( 
.A1(n_2902),
.A2(n_2903),
.B1(n_2906),
.B2(n_2896),
.C(n_2907),
.Y(n_2910)
);

AOI221x1_ASAP7_75t_L g2911 ( 
.A1(n_2904),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2898),
.A2(n_2481),
.B(n_2260),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2908),
.A2(n_2481),
.B(n_2260),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2896),
.B(n_2260),
.Y(n_2914)
);

OAI221xp5_ASAP7_75t_L g2915 ( 
.A1(n_2898),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.C(n_115),
.Y(n_2915)
);

NAND4xp25_ASAP7_75t_SL g2916 ( 
.A(n_2903),
.B(n_117),
.C(n_114),
.D(n_116),
.Y(n_2916)
);

OAI21xp33_ASAP7_75t_SL g2917 ( 
.A1(n_2896),
.A2(n_118),
.B(n_119),
.Y(n_2917)
);

AOI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2902),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2902),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2896),
.Y(n_2920)
);

NAND2xp33_ASAP7_75t_SL g2921 ( 
.A(n_2896),
.B(n_122),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_R g2922 ( 
.A(n_2896),
.B(n_125),
.Y(n_2922)
);

OAI211xp5_ASAP7_75t_SL g2923 ( 
.A1(n_2905),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_2923)
);

AOI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2897),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_2924)
);

AOI211xp5_ASAP7_75t_L g2925 ( 
.A1(n_2897),
.A2(n_132),
.B(n_129),
.C(n_131),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2920),
.Y(n_2926)
);

AOI211xp5_ASAP7_75t_L g2927 ( 
.A1(n_2915),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_2927)
);

AOI222xp33_ASAP7_75t_L g2928 ( 
.A1(n_2924),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.C1(n_138),
.C2(n_141),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2925),
.B(n_2918),
.Y(n_2929)
);

OAI211xp5_ASAP7_75t_L g2930 ( 
.A1(n_2917),
.A2(n_2910),
.B(n_2909),
.C(n_2911),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2919),
.Y(n_2931)
);

OAI221xp5_ASAP7_75t_L g2932 ( 
.A1(n_2921),
.A2(n_138),
.B1(n_143),
.B2(n_145),
.C(n_146),
.Y(n_2932)
);

OAI211xp5_ASAP7_75t_L g2933 ( 
.A1(n_2922),
.A2(n_148),
.B(n_145),
.C(n_147),
.Y(n_2933)
);

AOI311xp33_ASAP7_75t_L g2934 ( 
.A1(n_2912),
.A2(n_148),
.A3(n_151),
.B(n_153),
.C(n_154),
.Y(n_2934)
);

A2O1A1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_2923),
.A2(n_157),
.B(n_151),
.C(n_156),
.Y(n_2935)
);

AOI221xp5_ASAP7_75t_L g2936 ( 
.A1(n_2916),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.C(n_160),
.Y(n_2936)
);

AND3x2_ASAP7_75t_L g2937 ( 
.A(n_2914),
.B(n_159),
.C(n_161),
.Y(n_2937)
);

OAI211xp5_ASAP7_75t_L g2938 ( 
.A1(n_2913),
.A2(n_165),
.B(n_162),
.C(n_163),
.Y(n_2938)
);

A2O1A1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2917),
.A2(n_165),
.B(n_162),
.C(n_163),
.Y(n_2939)
);

AOI221x1_ASAP7_75t_L g2940 ( 
.A1(n_2921),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_2940)
);

NOR2x1p5_ASAP7_75t_L g2941 ( 
.A(n_2926),
.B(n_2929),
.Y(n_2941)
);

NAND3x1_ASAP7_75t_SL g2942 ( 
.A(n_2936),
.B(n_169),
.C(n_171),
.Y(n_2942)
);

OAI22xp5_ASAP7_75t_SL g2943 ( 
.A1(n_2932),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_2943)
);

OAI321xp33_ASAP7_75t_L g2944 ( 
.A1(n_2930),
.A2(n_173),
.A3(n_175),
.B1(n_176),
.B2(n_177),
.C(n_179),
.Y(n_2944)
);

AOI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2939),
.A2(n_1180),
.B(n_179),
.Y(n_2945)
);

NAND3xp33_ASAP7_75t_SL g2946 ( 
.A(n_2927),
.B(n_2928),
.C(n_2933),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2937),
.B(n_180),
.Y(n_2947)
);

AOI31xp33_ASAP7_75t_L g2948 ( 
.A1(n_2931),
.A2(n_180),
.A3(n_181),
.B(n_182),
.Y(n_2948)
);

NAND2xp33_ASAP7_75t_SL g2949 ( 
.A(n_2940),
.B(n_184),
.Y(n_2949)
);

NOR3xp33_ASAP7_75t_L g2950 ( 
.A(n_2935),
.B(n_185),
.C(n_186),
.Y(n_2950)
);

AOI21xp33_ASAP7_75t_SL g2951 ( 
.A1(n_2938),
.A2(n_187),
.B(n_188),
.Y(n_2951)
);

AOI221xp5_ASAP7_75t_L g2952 ( 
.A1(n_2934),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.C(n_193),
.Y(n_2952)
);

AND2x2_ASAP7_75t_SL g2953 ( 
.A(n_2950),
.B(n_193),
.Y(n_2953)
);

OA22x2_ASAP7_75t_L g2954 ( 
.A1(n_2943),
.A2(n_195),
.B1(n_196),
.B2(n_1468),
.Y(n_2954)
);

AOI221xp5_ASAP7_75t_L g2955 ( 
.A1(n_2944),
.A2(n_196),
.B1(n_884),
.B2(n_886),
.C(n_1125),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2947),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2942),
.Y(n_2957)
);

OAI221xp5_ASAP7_75t_SL g2958 ( 
.A1(n_2952),
.A2(n_1244),
.B1(n_1270),
.B2(n_202),
.C(n_203),
.Y(n_2958)
);

NOR2xp67_ASAP7_75t_L g2959 ( 
.A(n_2951),
.B(n_199),
.Y(n_2959)
);

NOR2xp67_ASAP7_75t_SL g2960 ( 
.A(n_2945),
.B(n_886),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2941),
.Y(n_2961)
);

NAND4xp25_ASAP7_75t_L g2962 ( 
.A(n_2946),
.B(n_1218),
.C(n_1197),
.D(n_1304),
.Y(n_2962)
);

NOR4xp75_ASAP7_75t_L g2963 ( 
.A(n_2949),
.B(n_2948),
.C(n_1304),
.D(n_210),
.Y(n_2963)
);

OAI22xp5_ASAP7_75t_SL g2964 ( 
.A1(n_2957),
.A2(n_1216),
.B1(n_1232),
.B2(n_1263),
.Y(n_2964)
);

NAND5xp2_ASAP7_75t_L g2965 ( 
.A(n_2956),
.B(n_201),
.C(n_204),
.D(n_213),
.E(n_215),
.Y(n_2965)
);

OAI22xp5_ASAP7_75t_L g2966 ( 
.A1(n_2961),
.A2(n_1468),
.B1(n_1270),
.B2(n_1244),
.Y(n_2966)
);

INVxp67_ASAP7_75t_SL g2967 ( 
.A(n_2959),
.Y(n_2967)
);

OAI211xp5_ASAP7_75t_L g2968 ( 
.A1(n_2955),
.A2(n_218),
.B(n_219),
.C(n_220),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_SL g2969 ( 
.A(n_2953),
.B(n_1326),
.Y(n_2969)
);

NAND3xp33_ASAP7_75t_SL g2970 ( 
.A(n_2963),
.B(n_223),
.C(n_226),
.Y(n_2970)
);

NOR3xp33_ASAP7_75t_L g2971 ( 
.A(n_2958),
.B(n_1127),
.C(n_1121),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2954),
.Y(n_2972)
);

NOR4xp25_ASAP7_75t_L g2973 ( 
.A(n_2960),
.B(n_2962),
.C(n_230),
.D(n_234),
.Y(n_2973)
);

OAI321xp33_ASAP7_75t_L g2974 ( 
.A1(n_2961),
.A2(n_227),
.A3(n_236),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2954),
.Y(n_2975)
);

NAND3x1_ASAP7_75t_L g2976 ( 
.A(n_2963),
.B(n_244),
.C(n_247),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2954),
.Y(n_2977)
);

NOR3xp33_ASAP7_75t_L g2978 ( 
.A(n_2961),
.B(n_875),
.C(n_1247),
.Y(n_2978)
);

AND4x1_ASAP7_75t_L g2979 ( 
.A(n_2973),
.B(n_248),
.C(n_249),
.D(n_253),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2967),
.B(n_255),
.Y(n_2980)
);

NAND2x1p5_ASAP7_75t_L g2981 ( 
.A(n_2972),
.B(n_1247),
.Y(n_2981)
);

NOR3xp33_ASAP7_75t_L g2982 ( 
.A(n_2975),
.B(n_875),
.C(n_259),
.Y(n_2982)
);

NOR4xp25_ASAP7_75t_L g2983 ( 
.A(n_2977),
.B(n_265),
.C(n_267),
.D(n_268),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_SL g2984 ( 
.A1(n_2970),
.A2(n_1235),
.B(n_275),
.Y(n_2984)
);

OR3x1_ASAP7_75t_L g2985 ( 
.A(n_2965),
.B(n_276),
.C(n_279),
.Y(n_2985)
);

INVx3_ASAP7_75t_L g2986 ( 
.A(n_2976),
.Y(n_2986)
);

INVxp67_ASAP7_75t_L g2987 ( 
.A(n_2969),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2985),
.Y(n_2988)
);

AOI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_2986),
.A2(n_2968),
.B1(n_2971),
.B2(n_2964),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2980),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2982),
.A2(n_2978),
.B1(n_2974),
.B2(n_2966),
.Y(n_2991)
);

NAND4xp75_ASAP7_75t_L g2992 ( 
.A(n_2979),
.B(n_280),
.C(n_281),
.D(n_286),
.Y(n_2992)
);

OAI22x1_ASAP7_75t_L g2993 ( 
.A1(n_2987),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_2993)
);

AOI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2984),
.A2(n_1332),
.B1(n_1326),
.B2(n_1209),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2981),
.A2(n_1197),
.B1(n_1290),
.B2(n_1279),
.Y(n_2995)
);

O2A1O1Ixp33_ASAP7_75t_SL g2996 ( 
.A1(n_2983),
.A2(n_1326),
.B(n_1332),
.C(n_302),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2985),
.Y(n_2997)
);

AOI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2985),
.A2(n_1332),
.B1(n_1287),
.B2(n_916),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2985),
.A2(n_1287),
.B1(n_916),
.B2(n_972),
.Y(n_2999)
);

AO22x1_ASAP7_75t_L g3000 ( 
.A1(n_2986),
.A2(n_916),
.B1(n_300),
.B2(n_305),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2985),
.A2(n_1232),
.B1(n_1216),
.B2(n_1279),
.Y(n_3001)
);

AOI22x1_ASAP7_75t_L g3002 ( 
.A1(n_2986),
.A2(n_297),
.B1(n_307),
.B2(n_311),
.Y(n_3002)
);

AOI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2985),
.A2(n_1287),
.B1(n_916),
.B2(n_972),
.Y(n_3003)
);

AO22x2_ASAP7_75t_L g3004 ( 
.A1(n_2986),
.A2(n_312),
.B1(n_316),
.B2(n_323),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2985),
.Y(n_3005)
);

INVxp67_ASAP7_75t_SL g3006 ( 
.A(n_2980),
.Y(n_3006)
);

AO22x2_ASAP7_75t_L g3007 ( 
.A1(n_2986),
.A2(n_324),
.B1(n_331),
.B2(n_334),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_SL g3008 ( 
.A1(n_2986),
.A2(n_916),
.B1(n_972),
.B2(n_338),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2985),
.Y(n_3009)
);

INVx3_ASAP7_75t_SL g3010 ( 
.A(n_3005),
.Y(n_3010)
);

BUFx6f_ASAP7_75t_L g3011 ( 
.A(n_2990),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2988),
.B(n_336),
.Y(n_3012)
);

OAI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2994),
.A2(n_1263),
.B1(n_1290),
.B2(n_1232),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2992),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2999),
.Y(n_3015)
);

NAND3xp33_ASAP7_75t_L g3016 ( 
.A(n_2997),
.B(n_3009),
.C(n_2989),
.Y(n_3016)
);

OAI31xp33_ASAP7_75t_SL g3017 ( 
.A1(n_3006),
.A2(n_337),
.A3(n_339),
.B(n_340),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_3003),
.B(n_341),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_3002),
.Y(n_3019)
);

NAND3xp33_ASAP7_75t_L g3020 ( 
.A(n_2998),
.B(n_2991),
.C(n_3008),
.Y(n_3020)
);

HB1xp67_ASAP7_75t_L g3021 ( 
.A(n_2993),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2995),
.A2(n_916),
.B1(n_972),
.B2(n_1339),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_3001),
.A2(n_916),
.B1(n_972),
.B2(n_1272),
.Y(n_3023)
);

AO22x2_ASAP7_75t_L g3024 ( 
.A1(n_2996),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_3004),
.Y(n_3025)
);

OAI31xp33_ASAP7_75t_L g3026 ( 
.A1(n_3004),
.A2(n_354),
.A3(n_356),
.B(n_357),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_3000),
.B(n_360),
.Y(n_3027)
);

INVx4_ASAP7_75t_L g3028 ( 
.A(n_3007),
.Y(n_3028)
);

AO22x2_ASAP7_75t_L g3029 ( 
.A1(n_2988),
.A2(n_362),
.B1(n_364),
.B2(n_369),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_3005),
.A2(n_972),
.B1(n_1216),
.B2(n_1339),
.Y(n_3030)
);

AOI22xp33_ASAP7_75t_L g3031 ( 
.A1(n_3005),
.A2(n_1263),
.B1(n_1290),
.B2(n_1339),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_3005),
.A2(n_1263),
.B1(n_1290),
.B2(n_1279),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2999),
.B(n_370),
.Y(n_3033)
);

AOI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2988),
.A2(n_1347),
.B1(n_1279),
.B2(n_1058),
.Y(n_3034)
);

AOI31xp33_ASAP7_75t_L g3035 ( 
.A1(n_2988),
.A2(n_375),
.A3(n_377),
.B(n_379),
.Y(n_3035)
);

OAI22xp33_ASAP7_75t_L g3036 ( 
.A1(n_2994),
.A2(n_1254),
.B1(n_1324),
.B2(n_1222),
.Y(n_3036)
);

AOI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_2988),
.A2(n_1058),
.B1(n_1254),
.B2(n_1324),
.Y(n_3037)
);

AOI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2988),
.A2(n_1278),
.B1(n_1259),
.B2(n_1237),
.Y(n_3038)
);

OAI31xp33_ASAP7_75t_L g3039 ( 
.A1(n_2996),
.A2(n_382),
.A3(n_386),
.B(n_393),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_3012),
.A2(n_1278),
.B1(n_1259),
.B2(n_1237),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_3016),
.A2(n_998),
.B1(n_1016),
.B2(n_1008),
.Y(n_3041)
);

INVx2_ASAP7_75t_SL g3042 ( 
.A(n_3024),
.Y(n_3042)
);

AOI22x1_ASAP7_75t_L g3043 ( 
.A1(n_3028),
.A2(n_399),
.B1(n_407),
.B2(n_409),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_3010),
.A2(n_1008),
.B1(n_1016),
.B2(n_1278),
.Y(n_3044)
);

OAI211xp5_ASAP7_75t_SL g3045 ( 
.A1(n_3025),
.A2(n_412),
.B(n_413),
.C(n_415),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_SL g3046 ( 
.A1(n_3019),
.A2(n_418),
.B1(n_1237),
.B2(n_1259),
.Y(n_3046)
);

OAI22x1_ASAP7_75t_L g3047 ( 
.A1(n_3021),
.A2(n_3014),
.B1(n_3020),
.B2(n_3018),
.Y(n_3047)
);

NAND4xp75_ASAP7_75t_L g3048 ( 
.A(n_3026),
.B(n_1113),
.C(n_1106),
.D(n_1114),
.Y(n_3048)
);

NAND4xp25_ASAP7_75t_L g3049 ( 
.A(n_3039),
.B(n_875),
.C(n_1106),
.D(n_1113),
.Y(n_3049)
);

NOR4xp75_ASAP7_75t_L g3050 ( 
.A(n_3027),
.B(n_1083),
.C(n_1149),
.D(n_1131),
.Y(n_3050)
);

OAI22xp5_ASAP7_75t_SL g3051 ( 
.A1(n_3011),
.A2(n_919),
.B1(n_937),
.B2(n_928),
.Y(n_3051)
);

XNOR2xp5_ASAP7_75t_L g3052 ( 
.A(n_3029),
.B(n_1114),
.Y(n_3052)
);

OAI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_3011),
.A2(n_1344),
.B1(n_1181),
.B2(n_1217),
.Y(n_3053)
);

AND3x4_ASAP7_75t_L g3054 ( 
.A(n_3017),
.B(n_1048),
.C(n_1097),
.Y(n_3054)
);

NAND4xp25_ASAP7_75t_L g3055 ( 
.A(n_3033),
.B(n_875),
.C(n_1149),
.D(n_1148),
.Y(n_3055)
);

OAI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_3015),
.A2(n_937),
.B1(n_928),
.B2(n_906),
.Y(n_3056)
);

AOI222xp33_ASAP7_75t_L g3057 ( 
.A1(n_3013),
.A2(n_919),
.B1(n_937),
.B2(n_906),
.C1(n_928),
.C2(n_882),
.Y(n_3057)
);

AOI221xp5_ASAP7_75t_L g3058 ( 
.A1(n_3036),
.A2(n_919),
.B1(n_937),
.B2(n_906),
.C(n_928),
.Y(n_3058)
);

OAI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_3031),
.A2(n_919),
.B1(n_906),
.B2(n_882),
.Y(n_3059)
);

OAI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_3032),
.A2(n_878),
.B1(n_882),
.B2(n_1075),
.Y(n_3060)
);

NOR2x1p5_ASAP7_75t_L g3061 ( 
.A(n_3035),
.B(n_1130),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_3038),
.B(n_878),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_3030),
.A2(n_3022),
.B1(n_3023),
.B2(n_3037),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_3034),
.A2(n_882),
.B1(n_1130),
.B2(n_1149),
.Y(n_3064)
);

OAI22x1_ASAP7_75t_L g3065 ( 
.A1(n_3028),
.A2(n_1344),
.B1(n_1181),
.B2(n_1097),
.Y(n_3065)
);

AOI211xp5_ASAP7_75t_L g3066 ( 
.A1(n_3012),
.A2(n_882),
.B(n_1129),
.C(n_1100),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_SL g3067 ( 
.A1(n_3028),
.A2(n_1048),
.B1(n_1054),
.B2(n_1071),
.Y(n_3067)
);

OAI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_3016),
.A2(n_1079),
.B1(n_1075),
.B2(n_1074),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_3061),
.A2(n_3054),
.B1(n_3042),
.B2(n_3049),
.Y(n_3069)
);

AOI22xp33_ASAP7_75t_L g3070 ( 
.A1(n_3046),
.A2(n_1085),
.B1(n_1100),
.B2(n_1056),
.Y(n_3070)
);

AOI22xp33_ASAP7_75t_L g3071 ( 
.A1(n_3047),
.A2(n_1085),
.B1(n_1100),
.B2(n_1056),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_3055),
.A2(n_1085),
.B1(n_1100),
.B2(n_1056),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_3045),
.A2(n_1085),
.B1(n_1100),
.B2(n_1056),
.Y(n_3073)
);

AOI31xp33_ASAP7_75t_L g3074 ( 
.A1(n_3052),
.A2(n_1071),
.A3(n_1054),
.B(n_1082),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_3053),
.A2(n_1085),
.B1(n_1129),
.B2(n_1017),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_3051),
.A2(n_1129),
.B1(n_1140),
.B2(n_1056),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_3067),
.A2(n_1129),
.B1(n_1021),
.B2(n_1140),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_3043),
.A2(n_1129),
.B1(n_1021),
.B2(n_1140),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_3041),
.A2(n_1129),
.B1(n_1021),
.B2(n_1140),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_3068),
.A2(n_3063),
.B1(n_3065),
.B2(n_3059),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_L g3081 ( 
.A1(n_3058),
.A2(n_1021),
.B1(n_1017),
.B2(n_1140),
.Y(n_3081)
);

AOI31xp33_ASAP7_75t_L g3082 ( 
.A1(n_3066),
.A2(n_1082),
.A3(n_1081),
.B(n_1074),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_L g3083 ( 
.A1(n_3060),
.A2(n_1017),
.B1(n_1021),
.B2(n_1140),
.Y(n_3083)
);

OAI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_3069),
.A2(n_3048),
.B1(n_3064),
.B2(n_3062),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_3074),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_SL g3086 ( 
.A1(n_3080),
.A2(n_3044),
.B1(n_3056),
.B2(n_3050),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_3071),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_3070),
.A2(n_3040),
.B1(n_3057),
.B2(n_1148),
.Y(n_3088)
);

AOI22xp5_ASAP7_75t_L g3089 ( 
.A1(n_3073),
.A2(n_1131),
.B1(n_1149),
.B2(n_1148),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_3078),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3082),
.Y(n_3091)
);

OAI22x1_ASAP7_75t_L g3092 ( 
.A1(n_3072),
.A2(n_3081),
.B1(n_3079),
.B2(n_3076),
.Y(n_3092)
);

OR3x1_ASAP7_75t_L g3093 ( 
.A(n_3083),
.B(n_3075),
.C(n_3077),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3074),
.Y(n_3094)
);

NAND4xp75_ASAP7_75t_L g3095 ( 
.A(n_3094),
.B(n_1081),
.C(n_1131),
.D(n_1021),
.Y(n_3095)
);

AOI221x1_ASAP7_75t_SL g3096 ( 
.A1(n_3084),
.A2(n_1017),
.B1(n_1055),
.B2(n_1053),
.C(n_1057),
.Y(n_3096)
);

OA21x2_ASAP7_75t_L g3097 ( 
.A1(n_3091),
.A2(n_3085),
.B(n_3087),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_3090),
.B(n_1057),
.Y(n_3098)
);

INVx1_ASAP7_75t_SL g3099 ( 
.A(n_3093),
.Y(n_3099)
);

AOI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_3086),
.A2(n_1053),
.B1(n_1057),
.B2(n_1055),
.Y(n_3100)
);

OA21x2_ASAP7_75t_L g3101 ( 
.A1(n_3089),
.A2(n_1057),
.B(n_1055),
.Y(n_3101)
);

AOI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_3092),
.A2(n_1055),
.B(n_1053),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3088),
.Y(n_3103)
);

AOI222xp33_ASAP7_75t_L g3104 ( 
.A1(n_3099),
.A2(n_1009),
.B1(n_1053),
.B2(n_989),
.C1(n_1285),
.C2(n_1282),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_3098),
.A2(n_989),
.B(n_1009),
.Y(n_3105)
);

AOI21xp33_ASAP7_75t_L g3106 ( 
.A1(n_3103),
.A2(n_876),
.B(n_951),
.Y(n_3106)
);

BUFx2_ASAP7_75t_L g3107 ( 
.A(n_3104),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3105),
.Y(n_3108)
);

NOR2x1_ASAP7_75t_L g3109 ( 
.A(n_3108),
.B(n_3097),
.Y(n_3109)
);

AOI221xp5_ASAP7_75t_L g3110 ( 
.A1(n_3109),
.A2(n_3102),
.B1(n_3106),
.B2(n_3107),
.C(n_3096),
.Y(n_3110)
);

AOI211xp5_ASAP7_75t_L g3111 ( 
.A1(n_3110),
.A2(n_3100),
.B(n_3095),
.C(n_3101),
.Y(n_3111)
);


endmodule