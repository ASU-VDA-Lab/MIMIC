module fake_jpeg_1756_n_378 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_0),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_53),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_16),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_13),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_70),
.Y(n_147)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_26),
.B(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_91),
.Y(n_116)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_88),
.Y(n_106)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_97),
.B(n_33),
.Y(n_114)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_40),
.B(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_14),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_14),
.C(n_13),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_22),
.C(n_38),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_98),
.Y(n_125)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_12),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_100),
.A2(n_102),
.B1(n_112),
.B2(n_114),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_48),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_53),
.A2(n_97),
.B1(n_89),
.B2(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_131),
.B1(n_138),
.B2(n_144),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_128),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_45),
.B1(n_20),
.B2(n_22),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_96),
.B1(n_3),
.B2(n_5),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_20),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_44),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_44),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_38),
.B(n_2),
.C(n_3),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_65),
.B(n_54),
.C(n_78),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_49),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_67),
.A2(n_43),
.B1(n_42),
.B2(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_95),
.Y(n_160)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_135),
.B(n_101),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_160),
.Y(n_208)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_162),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_58),
.B1(n_51),
.B2(n_52),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_135),
.B(n_143),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_38),
.B1(n_94),
.B2(n_92),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_112),
.A2(n_100),
.B1(n_77),
.B2(n_102),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_169),
.B1(n_176),
.B2(n_197),
.Y(n_201)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_144),
.B1(n_151),
.B2(n_152),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_12),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_171),
.B(n_182),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_183),
.Y(n_199)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_175),
.Y(n_206)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_177),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_184),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_121),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_133),
.B1(n_150),
.B2(n_135),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_3),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_7),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_187),
.Y(n_202)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_191),
.Y(n_216)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_7),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_132),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_115),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_150),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_219),
.B1(n_169),
.B2(n_166),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_119),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_218),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_99),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_228),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_211),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_172),
.B(n_149),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_163),
.A2(n_148),
.B1(n_111),
.B2(n_142),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_134),
.B1(n_110),
.B2(n_140),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_176),
.B1(n_168),
.B2(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_141),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_185),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_154),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_184),
.C(n_190),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_190),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_236),
.B1(n_202),
.B2(n_216),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_248),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_190),
.B1(n_208),
.B2(n_220),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_239),
.B(n_254),
.Y(n_274)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_227),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_186),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_158),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_250),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_219),
.B1(n_211),
.B2(n_209),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_252),
.B1(n_206),
.B2(n_215),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_101),
.B(n_162),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_200),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_201),
.A2(n_197),
.B1(n_142),
.B2(n_108),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_170),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_225),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_198),
.B(n_187),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_202),
.B(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_199),
.B1(n_218),
.B2(n_226),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_258),
.B1(n_264),
.B2(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_226),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_276),
.C(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_273),
.Y(n_290)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_203),
.B1(n_217),
.B2(n_224),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_266),
.B1(n_237),
.B2(n_250),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_277),
.B(n_254),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_202),
.B1(n_216),
.B2(n_173),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_212),
.B1(n_224),
.B2(n_207),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_270),
.B1(n_237),
.B2(n_234),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_236),
.A2(n_212),
.B1(n_224),
.B2(n_207),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_210),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_210),
.C(n_195),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_217),
.B(n_200),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_177),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_244),
.C(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_205),
.Y(n_279)
);

AO221x1_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_253),
.B1(n_252),
.B2(n_256),
.C(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_280),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_233),
.B1(n_272),
.B2(n_238),
.Y(n_318)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_294),
.B1(n_270),
.B2(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_232),
.C(n_234),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_274),
.C(n_269),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_267),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_258),
.B1(n_266),
.B2(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_300),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_232),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_245),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_261),
.B(n_240),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_205),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_262),
.B(n_252),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

OAI322xp33_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_273),
.A3(n_254),
.B1(n_257),
.B2(n_263),
.C1(n_260),
.C2(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_301),
.B(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_312),
.B1(n_318),
.B2(n_286),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_276),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_311),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_310),
.Y(n_323)
);

NOR4xp25_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_251),
.C(n_277),
.D(n_260),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_262),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_285),
.A2(n_293),
.B1(n_300),
.B2(n_292),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_283),
.B(n_299),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_288),
.C(n_291),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_327),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_331),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_290),
.B(n_284),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_324),
.C(n_314),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_305),
.B(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_318),
.B1(n_316),
.B2(n_304),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_290),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_292),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_311),
.CI(n_305),
.CON(n_331),
.SN(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_287),
.C(n_281),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_313),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_321),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_339),
.Y(n_350)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_344),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_324),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_306),
.B1(n_297),
.B2(n_313),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_345),
.B(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_347),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_320),
.B(n_326),
.Y(n_348)
);

AOI21xp33_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_338),
.B(n_334),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_341),
.B(n_306),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_352),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_337),
.A2(n_333),
.B1(n_280),
.B2(n_331),
.Y(n_351)
);

AOI21x1_ASAP7_75t_L g360 ( 
.A1(n_351),
.A2(n_331),
.B(n_323),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_342),
.B(n_319),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_350),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_358),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_344),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_346),
.A2(n_323),
.B(n_329),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_360),
.B(n_361),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_348),
.A2(n_335),
.B1(n_343),
.B2(n_328),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_351),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_364),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_357),
.A2(n_354),
.B1(n_335),
.B2(n_328),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_272),
.C(n_243),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_366),
.C(n_217),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_357),
.A2(n_137),
.B(n_174),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_108),
.C(n_164),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_372),
.C(n_109),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_130),
.C(n_109),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_373),
.A2(n_374),
.B(n_375),
.C(n_8),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_189),
.C(n_167),
.Y(n_375)
);

AOI321xp33_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_155),
.A3(n_161),
.B1(n_111),
.B2(n_148),
.C(n_11),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_377),
.Y(n_378)
);


endmodule