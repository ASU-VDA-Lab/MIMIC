module fake_jpeg_21475_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_31),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_26),
.B(n_16),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_23),
.B1(n_30),
.B2(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_84),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_48),
.A3(n_19),
.B1(n_17),
.B2(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_71),
.Y(n_94)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_75),
.B1(n_61),
.B2(n_44),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_38),
.B1(n_34),
.B2(n_28),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_17),
.B1(n_27),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_24),
.B1(n_51),
.B2(n_55),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_38),
.B1(n_34),
.B2(n_27),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_85),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_21),
.B1(n_32),
.B2(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_31),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_93),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_110),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_115),
.B1(n_85),
.B2(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_16),
.B(n_18),
.C(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_31),
.Y(n_133)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_69),
.B1(n_87),
.B2(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_13),
.C(n_8),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_29),
.B1(n_20),
.B2(n_31),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_79),
.B(n_64),
.C(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_116),
.A2(n_119),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_121),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_68),
.B(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_68),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_83),
.B(n_72),
.C(n_66),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_83),
.C(n_72),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_142),
.C(n_59),
.Y(n_162)
);

OAI22x1_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_72),
.B1(n_85),
.B2(n_18),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_18),
.B1(n_59),
.B2(n_20),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_16),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_82),
.B1(n_81),
.B2(n_57),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_141),
.B1(n_113),
.B2(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_26),
.B(n_28),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_16),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_37),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_102),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_57),
.B1(n_47),
.B2(n_36),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_37),
.C(n_36),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_93),
.B1(n_95),
.B2(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_144),
.B1(n_149),
.B2(n_165),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_109),
.B1(n_103),
.B2(n_97),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_152),
.B1(n_161),
.B2(n_166),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_114),
.A3(n_26),
.B1(n_29),
.B2(n_20),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_150),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_101),
.B1(n_98),
.B2(n_36),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_35),
.B1(n_62),
.B2(n_14),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_154),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_26),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_156),
.B(n_162),
.CI(n_0),
.CON(n_199),
.SN(n_199)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_160),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_59),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_139),
.B(n_129),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_62),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_116),
.B1(n_127),
.B2(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_29),
.B1(n_20),
.B2(n_28),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_118),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_141),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_134),
.C(n_125),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_181),
.B(n_185),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_184),
.C(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_134),
.B(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_190),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_130),
.C(n_139),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_130),
.B1(n_20),
.B2(n_9),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_189),
.B1(n_193),
.B2(n_161),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_167),
.A2(n_148),
.B1(n_157),
.B2(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_188),
.B1(n_152),
.B2(n_156),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_29),
.B1(n_28),
.B2(n_2),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_13),
.B1(n_11),
.B2(n_9),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_11),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_154),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_200),
.B(n_172),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_206),
.C(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_171),
.C(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_208),
.B1(n_179),
.B2(n_174),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_211),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

FAx1_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_146),
.CI(n_158),
.CON(n_215),
.SN(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_155),
.C(n_11),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_174),
.B(n_189),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_197),
.B1(n_173),
.B2(n_175),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_0),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_1),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_199),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_212),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_199),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_178),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_178),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_219),
.B(n_210),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_241),
.B1(n_204),
.B2(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_195),
.C(n_175),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_218),
.C(n_205),
.Y(n_246)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_179),
.B1(n_173),
.B2(n_194),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_252),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_259),
.B1(n_248),
.B2(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_220),
.C(n_214),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_238),
.C(n_231),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_242),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_215),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_229),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_201),
.B1(n_215),
.B2(n_194),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_226),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_193),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_268),
.C(n_271),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_239),
.B(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_230),
.C(n_237),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_237),
.C(n_3),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_273),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_250),
.B1(n_245),
.B2(n_259),
.Y(n_274)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_247),
.B(n_258),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_263),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_268),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_247),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_251),
.B1(n_5),
.B2(n_7),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_275),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_279),
.A2(n_4),
.B(n_7),
.Y(n_292)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_4),
.B(n_7),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_281),
.B(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_297),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_286),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_282),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_284),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_289),
.C(n_288),
.Y(n_303)
);

O2A1O1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.C(n_301),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_302),
.B(n_299),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_298),
.B(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_300),
.C(n_304),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_277),
.B(n_294),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_294),
.Y(n_311)
);


endmodule