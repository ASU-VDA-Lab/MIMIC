module fake_jpeg_28967_n_488 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_488);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_488;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_51),
.Y(n_149)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_29),
.B(n_13),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_13),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_32),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_87),
.B(n_47),
.Y(n_140)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_46),
.B(n_13),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_93),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_12),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_98),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_102),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_153),
.B1(n_38),
.B2(n_31),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_41),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_26),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_51),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_51),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_38),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_150),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_79),
.B(n_0),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_70),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_58),
.B(n_35),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_84),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_54),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_158),
.A2(n_114),
.B1(n_72),
.B2(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_161),
.Y(n_219)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_75),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_188),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_170),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_184),
.Y(n_215)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_83),
.B1(n_90),
.B2(n_60),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_176),
.B1(n_204),
.B2(n_149),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_88),
.B1(n_93),
.B2(n_71),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx11_ASAP7_75t_SL g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_59),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_181),
.B(n_189),
.Y(n_238)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_53),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_193),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_34),
.B(n_45),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_105),
.B(n_145),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_236)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_42),
.Y(n_247)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_196),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_107),
.B(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_41),
.Y(n_213)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_201),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_133),
.A2(n_93),
.B1(n_71),
.B2(n_61),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_246)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_147),
.C(n_143),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_197),
.C(n_185),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_143),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_130),
.B1(n_140),
.B2(n_73),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_231),
.B1(n_127),
.B2(n_165),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_122),
.B1(n_62),
.B2(n_146),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_223),
.A2(n_228),
.B1(n_245),
.B2(n_134),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_155),
.B1(n_154),
.B2(n_144),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_154),
.B1(n_133),
.B2(n_34),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_163),
.B(n_47),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_249),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_181),
.A2(n_106),
.B1(n_111),
.B2(n_123),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_186),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_115),
.B1(n_123),
.B2(n_134),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_172),
.B(n_45),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_171),
.B(n_67),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_22),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_257),
.C(n_239),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_168),
.C(n_78),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_178),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_263),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_175),
.B(n_176),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_274),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_157),
.B(n_169),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_281),
.B(n_219),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_207),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_265),
.B(n_269),
.Y(n_300)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_204),
.B(n_187),
.C(n_200),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_268),
.A2(n_290),
.B(n_218),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_187),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_271),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_217),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_278),
.B1(n_282),
.B2(n_237),
.Y(n_311)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_276),
.B(n_279),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_223),
.B1(n_246),
.B2(n_226),
.Y(n_299)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_285),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_27),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_222),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_288),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_286),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_213),
.B(n_209),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_229),
.B(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_227),
.B(n_190),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_127),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_296),
.C(n_321),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_289),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_310),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_238),
.C(n_225),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_299),
.B1(n_268),
.B2(n_255),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_229),
.B(n_235),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_305),
.A2(n_0),
.B(n_1),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_214),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_270),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_211),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_230),
.B1(n_240),
.B2(n_239),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_299),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_254),
.A2(n_230),
.B1(n_240),
.B2(n_182),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_254),
.A2(n_192),
.B1(n_203),
.B2(n_206),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_235),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_324),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_283),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_254),
.A2(n_237),
.B1(n_243),
.B2(n_225),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_274),
.B1(n_266),
.B2(n_275),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_257),
.B(n_243),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_261),
.A2(n_233),
.B1(n_252),
.B2(n_237),
.Y(n_322)
);

OAI22x1_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_268),
.B1(n_255),
.B2(n_262),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_253),
.A2(n_252),
.A3(n_241),
.B1(n_233),
.B2(n_22),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_258),
.B(n_219),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_340),
.B1(n_315),
.B2(n_313),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_330),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_292),
.C(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_332),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_303),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_333),
.Y(n_377)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_334),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_335),
.A2(n_349),
.B1(n_353),
.B2(n_319),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_300),
.B(n_280),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_345),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_339),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_316),
.B(n_281),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_295),
.A2(n_269),
.B1(n_290),
.B2(n_268),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_344),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_283),
.B1(n_282),
.B2(n_278),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_317),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_166),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_347),
.B(n_348),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_307),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_91),
.B1(n_96),
.B2(n_74),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_303),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_354),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_293),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_329),
.C(n_301),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_48),
.B1(n_37),
.B2(n_3),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_306),
.B(n_296),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_362),
.C(n_382),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_294),
.B(n_324),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_358),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_361),
.A2(n_326),
.B1(n_338),
.B2(n_328),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_352),
.C(n_301),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_336),
.B(n_317),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_366),
.B(n_371),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_367),
.A2(n_374),
.B(n_364),
.Y(n_403)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_332),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_341),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_351),
.B(n_337),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_328),
.A2(n_318),
.B(n_305),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_376),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_294),
.Y(n_378)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_318),
.Y(n_379)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_333),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_323),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_343),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_310),
.C(n_308),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_334),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_377),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_395),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_372),
.A2(n_361),
.B1(n_363),
.B2(n_379),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_391),
.A2(n_398),
.B1(n_405),
.B2(n_408),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_344),
.C(n_339),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_396),
.C(n_406),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_376),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_394),
.B(n_400),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_350),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_349),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_372),
.A2(n_339),
.B1(n_346),
.B2(n_353),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_340),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_364),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_402),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_403),
.A2(n_407),
.B(n_370),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_363),
.A2(n_346),
.B1(n_309),
.B2(n_308),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_309),
.C(n_22),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_374),
.A2(n_48),
.B(n_27),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_381),
.C(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_411),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_360),
.C(n_378),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_418),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_370),
.C(n_377),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_420),
.Y(n_430)
);

INVx13_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_424),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_416),
.B(n_417),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_368),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_374),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_403),
.B(n_402),
.CI(n_391),
.CON(n_420),
.SN(n_420)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_359),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_427),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_426),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_384),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_406),
.C(n_404),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_431),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_396),
.C(n_387),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_434),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_388),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_389),
.B1(n_398),
.B2(n_405),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_420),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_423),
.A2(n_407),
.B(n_386),
.Y(n_438)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_438),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_425),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_419),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_442),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_409),
.C(n_413),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_444),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_415),
.C(n_416),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_456),
.B1(n_446),
.B2(n_439),
.Y(n_466)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_448),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_440),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_450),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_415),
.C(n_418),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_422),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_452),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_420),
.C(n_426),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_439),
.A2(n_412),
.B(n_384),
.Y(n_453)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_453),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_437),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_447),
.B(n_443),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_460),
.B(n_464),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_437),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_465),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_432),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_466),
.B(n_467),
.C(n_448),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_454),
.A2(n_365),
.B1(n_408),
.B2(n_414),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_473),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_444),
.C(n_450),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_471),
.B(n_4),
.Y(n_478)
);

O2A1O1Ixp33_ASAP7_75t_SL g472 ( 
.A1(n_458),
.A2(n_459),
.B(n_462),
.C(n_461),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_472),
.A2(n_474),
.B1(n_467),
.B2(n_463),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_462),
.A2(n_365),
.B(n_27),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_466),
.A2(n_1),
.B(n_2),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_476),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_1),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_478),
.A2(n_11),
.B(n_6),
.Y(n_481)
);

A2O1A1O1Ixp25_ASAP7_75t_L g479 ( 
.A1(n_477),
.A2(n_468),
.B(n_474),
.C(n_8),
.D(n_9),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_5),
.B(n_6),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_5),
.C(n_6),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_483),
.C(n_480),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_484),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_11),
.C(n_9),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_486),
.B(n_9),
.Y(n_487)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_487),
.B(n_10),
.CI(n_11),
.CON(n_488),
.SN(n_488)
);


endmodule