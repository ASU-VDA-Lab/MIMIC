module fake_jpeg_18313_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_53),
.Y(n_82)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_60),
.B1(n_54),
.B2(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_91),
.B1(n_80),
.B2(n_62),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_60),
.B1(n_65),
.B2(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_81),
.B1(n_53),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_103),
.B1(n_64),
.B2(n_66),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_101),
.B1(n_105),
.B2(n_64),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_65),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_86),
.B1(n_90),
.B2(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_78),
.B1(n_77),
.B2(n_70),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_67),
.B1(n_55),
.B2(n_68),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_115),
.B(n_4),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_73),
.Y(n_110)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_117),
.CI(n_72),
.CON(n_126),
.SN(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_120),
.B1(n_121),
.B2(n_1),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_47),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_0),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_107),
.C(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_130),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_133),
.B(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_23),
.B(n_43),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_116),
.B(n_7),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_123),
.B1(n_129),
.B2(n_125),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_6),
.B(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_140),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_137),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_139),
.B1(n_9),
.B2(n_12),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_44),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_8),
.C(n_13),
.Y(n_150)
);

OAI21x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_14),
.B(n_15),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_17),
.Y(n_152)
);

OAI321xp33_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_19),
.A3(n_27),
.B1(n_28),
.B2(n_29),
.C(n_34),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_36),
.Y(n_154)
);


endmodule