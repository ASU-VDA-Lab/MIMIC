module fake_jpeg_28386_n_82 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_17),
.C(n_21),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_12),
.B1(n_16),
.B2(n_14),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_40),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_15),
.B(n_20),
.C(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_51),
.B1(n_33),
.B2(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_11),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_53),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_42),
.C(n_51),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.C(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_50),
.C(n_30),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_65),
.B(n_2),
.Y(n_73)
);

OAI322xp33_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_53),
.A3(n_14),
.B1(n_9),
.B2(n_16),
.C1(n_6),
.C2(n_48),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_6),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_65),
.B1(n_67),
.B2(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_76),
.A2(n_1),
.B1(n_3),
.B2(n_18),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_77),
.C(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_1),
.Y(n_82)
);


endmodule