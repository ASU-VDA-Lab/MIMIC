module fake_jpeg_17069_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

HB1xp67_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_25),
.B1(n_12),
.B2(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_13),
.C(n_18),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_17),
.B(n_11),
.C(n_12),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_39),
.B1(n_41),
.B2(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_26),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_48),
.C(n_50),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_45),
.C(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

AOI21x1_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_62),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_2),
.B(n_3),
.Y(n_61)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_50),
.B(n_52),
.C(n_2),
.D(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_45),
.C(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_55),
.B1(n_59),
.B2(n_56),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_71),
.Y(n_77)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_75),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_79),
.B(n_61),
.Y(n_81)
);

AOI21x1_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_72),
.B(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_81),
.C(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_4),
.C(n_6),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_7),
.C(n_8),
.Y(n_84)
);


endmodule