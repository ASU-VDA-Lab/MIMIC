module fake_jpeg_17090_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_8),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_9),
.B(n_6),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_11),
.B1(n_9),
.B2(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_32),
.B(n_26),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_25),
.B(n_24),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_29),
.C(n_26),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.C(n_17),
.Y(n_36)
);

OAI322xp33_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_26),
.A3(n_28),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_13),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.C(n_16),
.Y(n_37)
);

OAI31xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_18),
.A3(n_8),
.B(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);


endmodule