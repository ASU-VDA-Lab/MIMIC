module fake_jpeg_14127_n_569 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_569);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_569;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_9),
.B(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_23),
.B(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_81),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_30),
.B(n_9),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_12),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_83),
.B(n_97),
.Y(n_148)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_12),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_34),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_117),
.Y(n_160)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_18),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_119),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_12),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_22),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_16),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_85),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_142),
.B(n_161),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_23),
.C(n_52),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_147),
.B(n_50),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_57),
.B1(n_56),
.B2(n_52),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_150),
.A2(n_200),
.B1(n_80),
.B2(n_111),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_32),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_32),
.B1(n_36),
.B2(n_49),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_152),
.A2(n_185),
.B1(n_196),
.B2(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_117),
.B(n_39),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_84),
.A2(n_39),
.B1(n_36),
.B2(n_49),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_167),
.A2(n_175),
.B1(n_38),
.B2(n_35),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_68),
.B(n_20),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_60),
.A2(n_33),
.B1(n_24),
.B2(n_47),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_90),
.B(n_66),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_50),
.B(n_43),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_78),
.A2(n_33),
.B1(n_24),
.B2(n_47),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_87),
.A2(n_57),
.B1(n_56),
.B2(n_25),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_44),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_201),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_82),
.A2(n_28),
.B1(n_35),
.B2(n_46),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_96),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_61),
.A2(n_66),
.B1(n_80),
.B2(n_69),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_61),
.B(n_44),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_205),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_148),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_206),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_208),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_236),
.Y(n_278)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_211),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_135),
.B(n_86),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_212),
.A2(n_43),
.B(n_124),
.Y(n_296)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_214),
.Y(n_307)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_215),
.Y(n_315)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_219),
.B(n_226),
.Y(n_308)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_220),
.Y(n_327)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_143),
.A2(n_88),
.B1(n_109),
.B2(n_105),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_148),
.B(n_25),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_222),
.B(n_227),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_184),
.Y(n_223)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_225),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_132),
.B(n_40),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_228),
.Y(n_323)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_137),
.Y(n_232)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_145),
.A2(n_131),
.B1(n_56),
.B2(n_57),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_234),
.A2(n_238),
.B1(n_244),
.B2(n_250),
.Y(n_320)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx4_ASAP7_75t_SL g302 ( 
.A(n_237),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_145),
.A2(n_56),
.B1(n_57),
.B2(n_92),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_192),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_241),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_243),
.Y(n_288)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_134),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_195),
.A2(n_57),
.B1(n_99),
.B2(n_91),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_248),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_246),
.A2(n_196),
.B1(n_21),
.B2(n_40),
.Y(n_289)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_247),
.Y(n_275)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_249),
.B(n_253),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_190),
.A2(n_89),
.B1(n_75),
.B2(n_70),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_200),
.A2(n_62),
.B1(n_74),
.B2(n_71),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_297)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_252),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_184),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_184),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_255),
.Y(n_281)
);

BUFx4f_ASAP7_75t_SL g256 ( 
.A(n_128),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_256),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_192),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_257),
.B(n_259),
.Y(n_287)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_127),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_130),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_128),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_138),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_158),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_133),
.Y(n_264)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_129),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_46),
.B(n_28),
.C(n_38),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_267),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_175),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_170),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_160),
.B(n_21),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_165),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_159),
.B1(n_178),
.B2(n_171),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_213),
.A2(n_217),
.A3(n_160),
.B1(n_206),
.B2(n_221),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_204),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_279),
.B(n_296),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_289),
.A2(n_309),
.B1(n_325),
.B2(n_328),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_216),
.A2(n_150),
.B1(n_189),
.B2(n_126),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_297),
.B1(n_317),
.B2(n_324),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_209),
.C(n_230),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_304),
.C(n_261),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_231),
.B(n_244),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_126),
.B1(n_189),
.B2(n_139),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_208),
.A2(n_65),
.B1(n_179),
.B2(n_202),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_250),
.A2(n_178),
.B1(n_171),
.B2(n_176),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_218),
.A2(n_141),
.B1(n_140),
.B2(n_169),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_229),
.A2(n_169),
.B1(n_166),
.B2(n_88),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_332),
.Y(n_379)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_330),
.Y(n_375)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_336),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_247),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_341),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_238),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_335),
.B(n_337),
.C(n_368),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_234),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_289),
.Y(n_372)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_265),
.B(n_256),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g373 ( 
.A1(n_340),
.A2(n_316),
.B(n_327),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g341 ( 
.A1(n_277),
.A2(n_252),
.B1(n_225),
.B2(n_243),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_269),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_343),
.B(n_346),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_282),
.B(n_214),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_353),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_263),
.B1(n_248),
.B2(n_273),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_345),
.A2(n_351),
.B1(n_358),
.B2(n_327),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_321),
.A2(n_207),
.B1(n_166),
.B2(n_228),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_317),
.A2(n_291),
.B1(n_320),
.B2(n_300),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_354),
.B(n_359),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_237),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_361),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_220),
.B(n_205),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_316),
.B(n_328),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_223),
.B1(n_240),
.B2(n_265),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_278),
.B(n_261),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_296),
.A2(n_256),
.B1(n_13),
.B2(n_16),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_367),
.B1(n_311),
.B2(n_318),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_363),
.A2(n_322),
.B(n_319),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_314),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_366),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_294),
.A2(n_14),
.B1(n_15),
.B2(n_2),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_SL g394 ( 
.A(n_365),
.B(n_302),
.C(n_303),
.Y(n_394)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_14),
.B1(n_15),
.B2(n_2),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_295),
.B(n_0),
.C(n_1),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_281),
.B(n_0),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_0),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_371),
.A2(n_373),
.B(n_378),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_397),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_392),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_334),
.A2(n_325),
.B1(n_288),
.B2(n_281),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_383),
.B1(n_384),
.B2(n_396),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_356),
.A2(n_298),
.B1(n_301),
.B2(n_292),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_280),
.B(n_275),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_398),
.B(n_371),
.Y(n_416)
);

OAI32xp33_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_280),
.A3(n_303),
.B1(n_319),
.B2(n_290),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_401),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_369),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_394),
.A2(n_342),
.B1(n_351),
.B2(n_360),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_356),
.A2(n_292),
.B1(n_283),
.B2(n_322),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_338),
.A2(n_307),
.B(n_323),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_330),
.A2(n_283),
.B1(n_299),
.B2(n_307),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_341),
.Y(n_419)
);

AOI32xp33_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_302),
.A3(n_305),
.B1(n_279),
.B2(n_323),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_405),
.A2(n_340),
.B(n_368),
.Y(n_425)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_406),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_331),
.B1(n_348),
.B2(n_339),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_410),
.B1(n_413),
.B2(n_414),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_409),
.B(n_425),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_380),
.A2(n_329),
.B1(n_332),
.B2(n_370),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_398),
.A2(n_357),
.B1(n_370),
.B2(n_341),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_341),
.B1(n_362),
.B2(n_340),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_400),
.A2(n_360),
.B(n_344),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_415),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_416),
.Y(n_452)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_381),
.B1(n_390),
.B2(n_394),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_337),
.B(n_335),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_401),
.Y(n_464)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_373),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_431),
.Y(n_437)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_424),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_341),
.B1(n_347),
.B2(n_364),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_426),
.A2(n_427),
.B1(n_434),
.B2(n_383),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_347),
.B1(n_366),
.B2(n_354),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_428),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_397),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_436),
.C(n_393),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_392),
.B(n_349),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_382),
.A2(n_367),
.B(n_358),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_413),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_390),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_435),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_375),
.A2(n_345),
.B1(n_350),
.B2(n_353),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_315),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_411),
.C(n_421),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_447),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_412),
.A2(n_378),
.B1(n_385),
.B2(n_399),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_450),
.B1(n_453),
.B2(n_462),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_372),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_412),
.A2(n_399),
.B1(n_375),
.B2(n_376),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_451),
.A2(n_454),
.B1(n_449),
.B2(n_428),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_424),
.A2(n_378),
.B1(n_376),
.B2(n_372),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_377),
.B1(n_396),
.B2(n_384),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_382),
.Y(n_455)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_455),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_423),
.B1(n_414),
.B2(n_431),
.Y(n_476)
);

AO22x1_ASAP7_75t_SL g458 ( 
.A1(n_422),
.A2(n_387),
.B1(n_389),
.B2(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_458),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_404),
.Y(n_460)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_417),
.A2(n_387),
.B(n_391),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_464),
.B(n_432),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_417),
.A2(n_403),
.B1(n_404),
.B2(n_388),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_408),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_433),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_429),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_472),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_473),
.B1(n_486),
.B2(n_461),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_463),
.B(n_403),
.Y(n_470)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_449),
.A2(n_416),
.B1(n_420),
.B2(n_423),
.Y(n_473)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_411),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_464),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_476),
.A2(n_438),
.B1(n_443),
.B2(n_439),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_425),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_477),
.B(n_442),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_448),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_478),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_407),
.Y(n_480)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_481),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_455),
.B(n_435),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_487),
.B1(n_456),
.B2(n_439),
.Y(n_500)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_450),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_483),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_458),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_452),
.A2(n_418),
.B(n_415),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_485),
.A2(n_444),
.B(n_452),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_454),
.A2(n_419),
.B1(n_410),
.B2(n_418),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_453),
.A2(n_440),
.B1(n_461),
.B2(n_438),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_488),
.A2(n_437),
.B(n_440),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_492),
.B(n_476),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_485),
.A2(n_437),
.B(n_460),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_495),
.A2(n_467),
.B(n_479),
.Y(n_518)
);

MAJx2_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_498),
.C(n_504),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_500),
.A2(n_508),
.B1(n_471),
.B2(n_443),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_468),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_488),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_503),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_468),
.B(n_451),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_472),
.B(n_458),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_506),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_481),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_490),
.B(n_477),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_511),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_496),
.B(n_467),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_475),
.C(n_483),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_520),
.C(n_523),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_514),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_502),
.A2(n_471),
.B(n_473),
.Y(n_515)
);

XNOR2x1_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_305),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_487),
.Y(n_517)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_518),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_469),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_521),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_486),
.C(n_479),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_466),
.C(n_406),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_466),
.C(n_459),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_497),
.C(n_459),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_515),
.A2(n_494),
.B1(n_499),
.B2(n_491),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_526),
.A2(n_528),
.B1(n_530),
.B2(n_523),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_520),
.A2(n_506),
.B(n_507),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_527),
.B(n_532),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_515),
.A2(n_491),
.B1(n_492),
.B2(n_505),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_495),
.B1(n_489),
.B2(n_434),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_535),
.C(n_524),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_315),
.C(n_290),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_536),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_539),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_512),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_516),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_543),
.Y(n_549)
);

AOI31xp33_ASAP7_75t_L g542 ( 
.A1(n_537),
.A2(n_514),
.A3(n_513),
.B(n_509),
.Y(n_542)
);

OAI21xp33_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_529),
.B(n_533),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_522),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_546),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_528),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_517),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_547),
.Y(n_553)
);

A2O1A1O1Ixp25_ASAP7_75t_L g550 ( 
.A1(n_546),
.A2(n_525),
.B(n_509),
.C(n_535),
.D(n_529),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_550),
.B(n_555),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_544),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_554),
.B(n_530),
.Y(n_557)
);

OAI21xp33_ASAP7_75t_L g556 ( 
.A1(n_548),
.A2(n_541),
.B(n_540),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_557),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_553),
.B(n_311),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_318),
.Y(n_562)
);

AOI21x1_ASAP7_75t_SL g560 ( 
.A1(n_552),
.A2(n_549),
.B(n_551),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_558),
.C(n_14),
.Y(n_563)
);

OAI321xp33_ASAP7_75t_L g564 ( 
.A1(n_562),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_5),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_563),
.A2(n_0),
.B(n_1),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_564),
.A2(n_565),
.B(n_561),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_2),
.B(n_3),
.Y(n_568)
);

BUFx24_ASAP7_75t_SL g569 ( 
.A(n_568),
.Y(n_569)
);


endmodule