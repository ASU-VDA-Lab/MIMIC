module fake_jpeg_11035_n_201 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_3),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_1),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_101),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_65),
.B1(n_75),
.B2(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_82),
.B1(n_78),
.B2(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_82),
.B1(n_65),
.B2(n_63),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_78),
.B1(n_61),
.B2(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_74),
.B1(n_61),
.B2(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_74),
.B1(n_81),
.B2(n_69),
.Y(n_127)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_67),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_129),
.C(n_60),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_80),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_133),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_131),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_71),
.B(n_4),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_77),
.B1(n_84),
.B2(n_70),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_66),
.B(n_79),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_1),
.Y(n_142)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_85),
.A3(n_76),
.B1(n_73),
.B2(n_59),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_144),
.B(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_30),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_145),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_34),
.B1(n_40),
.B2(n_42),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_55),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_8),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_37),
.C(n_53),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_139),
.C(n_45),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_161),
.B1(n_165),
.B2(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_13),
.B1(n_17),
.B2(n_19),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_134),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_54),
.B1(n_35),
.B2(n_38),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_135),
.B1(n_147),
.B2(n_47),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_177),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_183),
.C(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_143),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_165),
.B1(n_163),
.B2(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_164),
.B1(n_180),
.B2(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_157),
.Y(n_189)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_176),
.A3(n_177),
.B1(n_173),
.B2(n_181),
.C(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_189),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_192),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_186),
.B(n_46),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_43),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_50),
.Y(n_201)
);


endmodule