module fake_netlist_5_1680_n_1696 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1696);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1696;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_49),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_110),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_92),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_43),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_27),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_35),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_91),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_61),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_49),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_51),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_34),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_52),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_30),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_43),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_54),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_23),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_17),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_130),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_33),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_75),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_6),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_9),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_35),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_5),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_4),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_27),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_122),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_119),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_44),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_104),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_58),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_46),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_30),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_39),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_11),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_107),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_143),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_88),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_41),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_28),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_115),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_94),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_70),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_33),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_56),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_100),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_106),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_21),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_125),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_18),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_111),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_7),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_138),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_1),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_74),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_89),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_42),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_39),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_55),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_13),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_71),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_96),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_38),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_109),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_76),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_80),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_24),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_137),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_84),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_105),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_101),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_69),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_48),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_145),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_21),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_158),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_187),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_161),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_161),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_289),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_206),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_151),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_153),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_161),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_161),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_157),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_205),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_205),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_205),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_205),
.Y(n_321)
);

BUFx6f_ASAP7_75t_SL g322 ( 
.A(n_181),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_173),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_246),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_187),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_162),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_292),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_160),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_162),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_186),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_153),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_201),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_186),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_191),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_192),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_163),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_164),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_176),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_192),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_201),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_203),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_166),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_168),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_203),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_227),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_152),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_171),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_215),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_261),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_220),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_227),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_220),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_175),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_221),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_177),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_221),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_223),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_223),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_229),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_154),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_178),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_180),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_229),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_156),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_184),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_303),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_344),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_271),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_164),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_315),
.A2(n_209),
.B1(n_324),
.B2(n_308),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_367),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_170),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_271),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_311),
.A2(n_341),
.B(n_334),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_369),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_319),
.B(n_275),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_324),
.A2(n_259),
.B1(n_284),
.B2(n_251),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_309),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_275),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_165),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_159),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_310),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_366),
.B(n_307),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_304),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_304),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_336),
.B(n_176),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_338),
.B(n_188),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_313),
.B(n_181),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_339),
.B(n_189),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_170),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_388),
.B(n_331),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_398),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_388),
.B(n_179),
.C(n_174),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_398),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_399),
.Y(n_449)
);

BUFx8_ASAP7_75t_SL g450 ( 
.A(n_374),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_317),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_431),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_398),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_330),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_385),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_340),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_399),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_346),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_404),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_385),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_347),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_SL g471 ( 
.A(n_436),
.B(n_355),
.C(n_371),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_348),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_386),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_416),
.B(n_313),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_416),
.B(n_353),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_371),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_359),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_401),
.B(n_339),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_409),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_376),
.B(n_361),
.Y(n_483)
);

CKINVDCx6p67_ASAP7_75t_R g484 ( 
.A(n_374),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_431),
.B(n_368),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_411),
.B(n_373),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_376),
.B(n_167),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_398),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_376),
.B(n_200),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_381),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_193),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_420),
.B(n_181),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_391),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_398),
.B(n_247),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_377),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_401),
.B(n_343),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_396),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_420),
.B(n_397),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_402),
.B(n_288),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_384),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_382),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_402),
.B(n_322),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_322),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_406),
.A2(n_322),
.B1(n_181),
.B2(n_248),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_194),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_382),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_397),
.A2(n_214),
.B1(n_262),
.B2(n_172),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_383),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_406),
.B(n_322),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_377),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_412),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_410),
.B(n_337),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_384),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_412),
.B(n_197),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_412),
.B(n_198),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_422),
.B(n_343),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_410),
.B(n_210),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_386),
.B(n_179),
.C(n_174),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_392),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_412),
.B(n_217),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_392),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_390),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_386),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_414),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_384),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_394),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_422),
.B(n_362),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_419),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_384),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

CKINVDCx6p67_ASAP7_75t_R g557 ( 
.A(n_391),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_386),
.A2(n_232),
.B1(n_264),
.B2(n_256),
.Y(n_558)
);

OAI21xp33_ASAP7_75t_SL g559 ( 
.A1(n_430),
.A2(n_248),
.B(n_242),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_390),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_386),
.B(n_202),
.C(n_185),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_386),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_434),
.Y(n_563)
);

CKINVDCx6p67_ASAP7_75t_R g564 ( 
.A(n_434),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_405),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_419),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_434),
.B(n_218),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_434),
.B(n_219),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_408),
.B(n_362),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_421),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_390),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_395),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_395),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_400),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_408),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_400),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_403),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_439),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_442),
.A2(n_272),
.B1(n_302),
.B2(n_290),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_580),
.B(n_390),
.Y(n_585)
);

AOI221xp5_ASAP7_75t_L g586 ( 
.A1(n_510),
.A2(n_272),
.B1(n_290),
.B2(n_280),
.C(n_265),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_390),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_533),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_457),
.B(n_190),
.C(n_182),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_459),
.B(n_384),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_491),
.B(n_403),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_450),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_533),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_459),
.B(n_384),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_491),
.B(n_417),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_459),
.B(n_384),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_483),
.B(n_478),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_417),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_492),
.B(n_375),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_442),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_527),
.B(n_418),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_439),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_441),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_474),
.B(n_204),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_563),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_507),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_375),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_497),
.A2(n_268),
.B1(n_222),
.B2(n_228),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_441),
.Y(n_610)
);

AOI221xp5_ASAP7_75t_L g611 ( 
.A1(n_535),
.A2(n_523),
.B1(n_528),
.B2(n_302),
.C(n_280),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_468),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_446),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_456),
.B(n_430),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_507),
.B(n_375),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_446),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_504),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_375),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_527),
.B(n_418),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_508),
.B(n_418),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_508),
.B(n_418),
.Y(n_622)
);

BUFx6f_ASAP7_75t_SL g623 ( 
.A(n_519),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_456),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_479),
.A2(n_238),
.B1(n_301),
.B2(n_299),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_451),
.B(n_230),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_508),
.B(n_379),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_463),
.B(n_379),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_548),
.B(n_418),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_471),
.B(n_211),
.C(n_240),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_463),
.B(n_379),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_548),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_443),
.B(n_433),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_449),
.Y(n_634)
);

NAND2x1_ASAP7_75t_L g635 ( 
.A(n_473),
.B(n_379),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_512),
.B(n_387),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_562),
.B(n_442),
.Y(n_638)
);

INVx8_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_453),
.B(n_207),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_481),
.B(n_387),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_442),
.B(n_418),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_448),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_481),
.B(n_387),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_452),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_452),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_506),
.B(n_387),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_460),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_506),
.B(n_389),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_468),
.B(n_425),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_516),
.B(n_389),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_468),
.B(n_425),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_521),
.B(n_389),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_472),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_489),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_487),
.B(n_216),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_515),
.B(n_389),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_465),
.B(n_433),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_464),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_461),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_479),
.A2(n_273),
.B1(n_297),
.B2(n_295),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_443),
.B(n_437),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_493),
.B(n_438),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_489),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_490),
.B(n_438),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_461),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_490),
.Y(n_672)
);

NAND2x1_ASAP7_75t_L g673 ( 
.A(n_473),
.B(n_423),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_572),
.A2(n_437),
.B(n_438),
.C(n_265),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_423),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_546),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_455),
.B(n_237),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_494),
.B(n_495),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_477),
.B(n_224),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_495),
.B(n_423),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_496),
.B(n_423),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_582),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_496),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_440),
.B(n_425),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_577),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_466),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_514),
.B(n_423),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_449),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_546),
.A2(n_564),
.B1(n_445),
.B2(n_532),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_440),
.B(n_425),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_440),
.B(n_425),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_445),
.B(n_345),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_485),
.A2(n_243),
.B1(n_244),
.B2(n_250),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_226),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_480),
.A2(n_258),
.B1(n_252),
.B2(n_253),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_462),
.B(n_266),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_522),
.B(n_185),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_559),
.A2(n_552),
.B(n_558),
.C(n_523),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_484),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_440),
.B(n_425),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_528),
.B(n_231),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_465),
.B(n_526),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_522),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_526),
.B(n_345),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_520),
.A2(n_195),
.B1(n_196),
.B2(n_199),
.C(n_276),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_525),
.B(n_274),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_466),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_524),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_524),
.B(n_202),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_539),
.B(n_208),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_539),
.B(n_208),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_500),
.B(n_534),
.C(n_486),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_542),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_531),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_537),
.A2(n_213),
.B1(n_212),
.B2(n_225),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_542),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_544),
.B(n_212),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_467),
.B(n_503),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_551),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_545),
.B(n_560),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_469),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_551),
.B(n_213),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_498),
.B(n_279),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_285),
.C(n_233),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_469),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_579),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_579),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_558),
.B(n_235),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_556),
.B(n_225),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_543),
.B(n_239),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_556),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_560),
.B(n_576),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_564),
.A2(n_291),
.B1(n_287),
.B2(n_282),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_578),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_578),
.B(n_234),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_547),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_560),
.B(n_576),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_349),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_581),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_502),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_559),
.A2(n_296),
.B(n_234),
.C(n_236),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_547),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_582),
.B(n_236),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_598),
.B(n_498),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_601),
.B(n_498),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_SL g752 ( 
.A1(n_740),
.A2(n_549),
.B1(n_458),
.B2(n_277),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_742),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_592),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_633),
.B(n_444),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_601),
.B(n_498),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_633),
.B(n_444),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_682),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_605),
.B(n_464),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_605),
.B(n_464),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_685),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_658),
.B(n_464),
.Y(n_763)
);

NOR2x1_ASAP7_75t_L g764 ( 
.A(n_614),
.B(n_537),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_685),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_601),
.B(n_529),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_730),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_640),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_660),
.B(n_624),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_730),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_666),
.B(n_588),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_700),
.A2(n_561),
.B(n_241),
.C(n_245),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_640),
.Y(n_774)
);

BUFx4f_ASAP7_75t_L g775 ( 
.A(n_639),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_658),
.B(n_513),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_696),
.B(n_519),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_745),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_612),
.B(n_619),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_585),
.B(n_513),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_706),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_607),
.A2(n_476),
.B1(n_473),
.B2(n_447),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_584),
.A2(n_561),
.B1(n_294),
.B2(n_298),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_696),
.B(n_519),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_584),
.A2(n_294),
.B1(n_298),
.B2(n_296),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_744),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_587),
.B(n_513),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_719),
.B(n_519),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_639),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_667),
.B(n_513),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_732),
.A2(n_603),
.B1(n_604),
.B2(n_583),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_606),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_716),
.A2(n_568),
.B1(n_567),
.B2(n_473),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_639),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_648),
.B(n_555),
.Y(n_797)
);

OR2x2_ASAP7_75t_SL g798 ( 
.A(n_589),
.B(n_549),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_583),
.A2(n_454),
.B1(n_488),
.B2(n_189),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_SL g800 ( 
.A1(n_747),
.A2(n_300),
.B1(n_269),
.B2(n_286),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_689),
.A2(n_454),
.B1(n_488),
.B2(n_555),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_732),
.A2(n_263),
.B(n_241),
.C(n_293),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_666),
.B(n_349),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_597),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_703),
.B(n_484),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_601),
.B(n_529),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_700),
.A2(n_263),
.B(n_293),
.C(n_283),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_612),
.B(n_529),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_634),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_694),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_657),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_734),
.A2(n_555),
.B1(n_281),
.B2(n_260),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_593),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_688),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_669),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_644),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_672),
.B(n_555),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_603),
.A2(n_257),
.B1(n_283),
.B2(n_270),
.Y(n_819)
);

AND2x6_ASAP7_75t_SL g820 ( 
.A(n_703),
.B(n_557),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_699),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_619),
.B(n_529),
.Y(n_822)
);

NOR2x1_ASAP7_75t_L g823 ( 
.A(n_636),
.B(n_550),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_646),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_636),
.B(n_550),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_647),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_650),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_604),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_734),
.A2(n_260),
.B1(n_249),
.B2(n_257),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_683),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_668),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_692),
.Y(n_832)
);

NOR2x2_ASAP7_75t_L g833 ( 
.A(n_611),
.B(n_557),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_679),
.A2(n_249),
.B1(n_270),
.B2(n_245),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_674),
.B(n_678),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_663),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_641),
.B(n_351),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_691),
.B(n_550),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_610),
.A2(n_254),
.B1(n_575),
.B2(n_573),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_610),
.B(n_613),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_613),
.B(n_529),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_705),
.B(n_710),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_671),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_722),
.A2(n_575),
.B(n_574),
.C(n_573),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_668),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_715),
.B(n_550),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_686),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_679),
.A2(n_254),
.B1(n_571),
.B2(n_475),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_L g850 ( 
.A1(n_718),
.A2(n_720),
.B1(n_735),
.B2(n_738),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_723),
.B(n_351),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_632),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_701),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_641),
.B(n_470),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_623),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_354),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_642),
.B(n_354),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_616),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_616),
.B(n_470),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_R g860 ( 
.A(n_623),
.B(n_59),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_717),
.A2(n_574),
.B1(n_571),
.B2(n_475),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_676),
.B(n_482),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_676),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_727),
.B(n_482),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_714),
.B(n_356),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_722),
.A2(n_501),
.B1(n_569),
.B2(n_566),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_653),
.A2(n_501),
.B(n_499),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_645),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_649),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_725),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_651),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_711),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_729),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_717),
.A2(n_505),
.B1(n_569),
.B2(n_566),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_670),
.B(n_499),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_728),
.B(n_356),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_637),
.B(n_505),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_724),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_358),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_630),
.B(n_625),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_724),
.B(n_358),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_628),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_675),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_746),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_591),
.A2(n_509),
.B1(n_554),
.B2(n_553),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_707),
.B(n_365),
.C(n_360),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_662),
.B(n_509),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_638),
.A2(n_530),
.B1(n_554),
.B2(n_553),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_673),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_638),
.A2(n_518),
.B1(n_511),
.B2(n_540),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_708),
.B(n_518),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_631),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_643),
.A2(n_536),
.B(n_511),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_713),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_665),
.B(n_363),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_695),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_680),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_655),
.B(n_536),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_736),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_721),
.B(n_530),
.Y(n_902)
);

CKINVDCx11_ASAP7_75t_R g903 ( 
.A(n_586),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_726),
.B(n_363),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_643),
.B(n_540),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_681),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_538),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_626),
.A2(n_538),
.B1(n_517),
.B2(n_427),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_739),
.B(n_517),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_687),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_748),
.Y(n_911)
);

BUFx4f_ASAP7_75t_SL g912 ( 
.A(n_602),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_595),
.B(n_432),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_600),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_697),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_659),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_608),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_599),
.B(n_432),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_746),
.A2(n_360),
.B(n_364),
.C(n_372),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_749),
.B(n_615),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_791),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_792),
.A2(n_590),
.B(n_594),
.Y(n_922)
);

AOI21xp33_ASAP7_75t_L g923 ( 
.A1(n_808),
.A2(n_749),
.B(n_882),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_814),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_884),
.A2(n_590),
.B(n_594),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_837),
.B(n_618),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_769),
.B(n_737),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_754),
.B(n_677),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_777),
.B(n_609),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_884),
.A2(n_596),
.B(n_627),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_858),
.A2(n_596),
.B(n_652),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_855),
.B(n_698),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_771),
.B(n_602),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_787),
.A2(n_702),
.B1(n_693),
.B2(n_690),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_898),
.B(n_364),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_791),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_845),
.A2(n_622),
.B(n_621),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_786),
.B(n_654),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_773),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_831),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_773),
.B(n_652),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_814),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_802),
.A2(n_620),
.B(n_693),
.C(n_690),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_888),
.A2(n_874),
.B(n_772),
.C(n_808),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_807),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_760),
.A2(n_620),
.B(n_629),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_868),
.A2(n_654),
.B(n_684),
.C(n_702),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_791),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_812),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_781),
.Y(n_950)
);

AO22x1_ASAP7_75t_L g951 ( 
.A1(n_805),
.A2(n_372),
.B1(n_370),
.B2(n_365),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_791),
.B(n_796),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_856),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_805),
.B(n_622),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_858),
.A2(n_621),
.B(n_684),
.Y(n_955)
);

AO32x1_ASAP7_75t_L g956 ( 
.A1(n_887),
.A2(n_370),
.A3(n_428),
.B1(n_427),
.B2(n_432),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_903),
.B(n_635),
.Y(n_957)
);

AO32x1_ASAP7_75t_L g958 ( 
.A1(n_799),
.A2(n_432),
.A3(n_428),
.B1(n_427),
.B2(n_426),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_915),
.A2(n_428),
.B1(n_427),
.B2(n_426),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_778),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_888),
.A2(n_428),
.B(n_426),
.C(n_7),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_787),
.A2(n_426),
.B1(n_425),
.B2(n_570),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_886),
.A2(n_425),
.B(n_570),
.C(n_541),
.Y(n_963)
);

OAI22x1_ASAP7_75t_L g964 ( 
.A1(n_866),
.A2(n_0),
.B1(n_2),
.B2(n_8),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_810),
.Y(n_965)
);

AO31x2_ASAP7_75t_L g966 ( 
.A1(n_772),
.A2(n_0),
.A3(n_2),
.B(n_8),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_874),
.B(n_10),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_752),
.B(n_12),
.C(n_13),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_831),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_SL g970 ( 
.A1(n_864),
.A2(n_570),
.B(n_541),
.C(n_149),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_896),
.B(n_14),
.Y(n_971)
);

OAI221xp5_ASAP7_75t_L g972 ( 
.A1(n_834),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_796),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_790),
.B(n_811),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_886),
.A2(n_541),
.B(n_570),
.C(n_19),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_850),
.A2(n_15),
.B(n_18),
.C(n_19),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_821),
.B(n_20),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_846),
.Y(n_978)
);

OA22x2_ASAP7_75t_L g979 ( 
.A1(n_800),
.A2(n_866),
.B1(n_771),
.B2(n_803),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_816),
.Y(n_980)
);

CKINVDCx16_ASAP7_75t_R g981 ( 
.A(n_815),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_916),
.B(n_20),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_775),
.B(n_768),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_803),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_759),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_916),
.B(n_869),
.Y(n_986)
);

NAND2x1_ASAP7_75t_L g987 ( 
.A(n_846),
.B(n_570),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_775),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_830),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_798),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_853),
.B(n_146),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_850),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_870),
.B(n_25),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_878),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_761),
.A2(n_541),
.B(n_131),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_794),
.B(n_26),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_763),
.A2(n_541),
.B(n_128),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_851),
.B(n_31),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_829),
.A2(n_764),
.B(n_854),
.C(n_873),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_878),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_776),
.A2(n_541),
.B(n_112),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_833),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_894),
.B(n_854),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_911),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_912),
.B(n_755),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_912),
.B(n_72),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_755),
.B(n_81),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_883),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_813),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_842),
.A2(n_47),
.B(n_48),
.C(n_86),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_793),
.B(n_97),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_793),
.B(n_904),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_828),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_757),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_845),
.A2(n_895),
.B(n_859),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_751),
.B(n_753),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_765),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_864),
.A2(n_893),
.B(n_809),
.C(n_822),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_762),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_780),
.A2(n_789),
.B(n_840),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_785),
.A2(n_819),
.B1(n_828),
.B2(n_839),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_904),
.B(n_883),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_914),
.B(n_917),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_770),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_852),
.B(n_885),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_767),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_809),
.A2(n_822),
.B(n_900),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_863),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_881),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_919),
.B(n_750),
.C(n_756),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_881),
.B(n_857),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_840),
.A2(n_918),
.B(n_913),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_879),
.A2(n_838),
.B(n_847),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_899),
.B(n_906),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_785),
.A2(n_819),
.B1(n_828),
.B2(n_839),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_880),
.B(n_901),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_783),
.Y(n_1037)
);

AO21x1_ASAP7_75t_L g1038 ( 
.A1(n_905),
.A2(n_900),
.B(n_877),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_897),
.A2(n_758),
.B1(n_795),
.B2(n_857),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_828),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_766),
.A2(n_806),
.B(n_889),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_880),
.B(n_901),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_857),
.A2(n_861),
.B1(n_876),
.B2(n_901),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_766),
.A2(n_806),
.B(n_907),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_881),
.B(n_875),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_910),
.B(n_872),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_774),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_871),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_861),
.A2(n_876),
.B1(n_835),
.B2(n_832),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_782),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_938),
.A2(n_877),
.B(n_756),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_960),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_1015),
.A2(n_1027),
.B(n_1020),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_945),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_949),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_922),
.A2(n_859),
.B(n_818),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_SL g1058 ( 
.A1(n_1021),
.A2(n_779),
.B(n_750),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_925),
.A2(n_835),
.B(n_902),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1003),
.B(n_872),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_930),
.A2(n_797),
.B(n_867),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_935),
.B(n_779),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1034),
.B(n_926),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_931),
.A2(n_801),
.B(n_841),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_939),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_953),
.B(n_844),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_986),
.B(n_872),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_929),
.A2(n_849),
.B(n_824),
.C(n_865),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_980),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_946),
.A2(n_919),
.A3(n_784),
.B(n_909),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1023),
.B(n_954),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_989),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1032),
.A2(n_841),
.B(n_892),
.Y(n_1073)
);

BUFx8_ASAP7_75t_L g1074 ( 
.A(n_988),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1033),
.A2(n_825),
.B(n_871),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_935),
.B(n_820),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_1013),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_981),
.B(n_860),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_920),
.A2(n_862),
.B(n_871),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_923),
.A2(n_890),
.B(n_908),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_923),
.A2(n_836),
.B(n_804),
.C(n_817),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1014),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_1013),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_950),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_927),
.A2(n_863),
.B1(n_848),
.B2(n_843),
.Y(n_1085)
);

INVx3_ASAP7_75t_SL g1086 ( 
.A(n_988),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_999),
.A2(n_825),
.B(n_871),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1021),
.A2(n_788),
.B1(n_826),
.B2(n_827),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1022),
.B(n_862),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1044),
.A2(n_823),
.B(n_891),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_937),
.A2(n_891),
.B(n_860),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_937),
.A2(n_1041),
.B(n_947),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1035),
.A2(n_891),
.B(n_955),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1018),
.A2(n_944),
.B(n_1049),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_997),
.A2(n_1001),
.B(n_995),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1043),
.A2(n_1035),
.B(n_1049),
.Y(n_1096)
);

NAND2x1_ASAP7_75t_L g1097 ( 
.A(n_1048),
.B(n_940),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1043),
.A2(n_934),
.B(n_1046),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_934),
.A2(n_943),
.B(n_963),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_988),
.Y(n_1100)
);

INVx8_ASAP7_75t_L g1101 ( 
.A(n_948),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1012),
.B(n_1025),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1038),
.A2(n_987),
.B(n_1011),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_921),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_969),
.A2(n_1028),
.B(n_978),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1030),
.A2(n_959),
.B(n_961),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_990),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1036),
.B(n_1042),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1050),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_921),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_994),
.B(n_1005),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_974),
.B(n_1039),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1048),
.A2(n_969),
.B(n_978),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_941),
.B(n_933),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_970),
.A2(n_975),
.B(n_993),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_SL g1117 ( 
.A1(n_972),
.A2(n_976),
.B(n_992),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_948),
.B(n_973),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_967),
.A2(n_977),
.B(n_982),
.C(n_1009),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_979),
.A2(n_1008),
.B1(n_1019),
.B2(n_1024),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_924),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_1004),
.A2(n_985),
.B(n_1017),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_983),
.A2(n_962),
.B(n_1037),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1040),
.B(n_1026),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_942),
.B(n_1045),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_956),
.A2(n_958),
.A3(n_996),
.B(n_964),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1016),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1029),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_956),
.A2(n_958),
.B(n_1007),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_SL g1131 ( 
.A1(n_1006),
.A2(n_1047),
.B(n_956),
.C(n_966),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_958),
.A2(n_979),
.B(n_1016),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_998),
.B(n_1031),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_951),
.A2(n_1010),
.B(n_984),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_921),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1002),
.A2(n_971),
.A3(n_966),
.B(n_957),
.Y(n_1136)
);

INVx6_ASAP7_75t_L g1137 ( 
.A(n_936),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_928),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_936),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_936),
.B(n_966),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_952),
.A2(n_973),
.B(n_991),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_952),
.B(n_968),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_991),
.A2(n_787),
.B1(n_584),
.B2(n_749),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_932),
.A2(n_1035),
.B(n_1021),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1015),
.A2(n_946),
.B(n_1018),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_923),
.A2(n_922),
.B(n_925),
.Y(n_1147)
);

NOR4xp25_ASAP7_75t_L g1148 ( 
.A(n_976),
.B(n_992),
.C(n_972),
.D(n_923),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_960),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1000),
.B(n_994),
.Y(n_1150)
);

AOI221x1_ASAP7_75t_L g1151 ( 
.A1(n_923),
.A2(n_605),
.B1(n_975),
.B2(n_1009),
.C(n_749),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1033),
.A2(n_619),
.B(n_612),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_945),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1003),
.B(n_598),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_953),
.B(n_456),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1033),
.A2(n_619),
.B(n_612),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_923),
.A2(n_808),
.B(n_944),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_960),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_923),
.A2(n_922),
.B(n_925),
.Y(n_1160)
);

BUFx2_ASAP7_75t_R g1161 ( 
.A(n_965),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_946),
.A2(n_868),
.A3(n_1038),
.B(n_963),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1013),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1003),
.B(n_598),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_939),
.Y(n_1167)
);

NOR2xp67_ASAP7_75t_SL g1168 ( 
.A(n_948),
.B(n_810),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_921),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_945),
.Y(n_1171)
);

NAND2x1_ASAP7_75t_L g1172 ( 
.A(n_1048),
.B(n_940),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1003),
.A2(n_787),
.B1(n_584),
.B2(n_749),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_925),
.A2(n_1033),
.B(n_922),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1015),
.A2(n_845),
.B(n_1027),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_945),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_925),
.A2(n_1033),
.B(n_922),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_925),
.A2(n_1033),
.B(n_922),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_965),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1128),
.B(n_1112),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1143),
.A2(n_1158),
.B1(n_1096),
.B2(n_1173),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1054),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_1077),
.B(n_1168),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1163),
.A2(n_1170),
.B(n_1164),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1175),
.A2(n_1093),
.B(n_1174),
.Y(n_1188)
);

CKINVDCx9p33_ASAP7_75t_R g1189 ( 
.A(n_1076),
.Y(n_1189)
);

BUFx4f_ASAP7_75t_SL g1190 ( 
.A(n_1057),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1143),
.A2(n_1173),
.B1(n_1094),
.B2(n_1107),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1115),
.B(n_1113),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1147),
.A2(n_1160),
.B(n_1099),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1147),
.A2(n_1160),
.B(n_1178),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1055),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1093),
.A2(n_1177),
.B(n_1061),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1119),
.A2(n_1117),
.B(n_1142),
.C(n_1148),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1069),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1094),
.A2(n_1098),
.B1(n_1071),
.B2(n_1063),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1115),
.B(n_1071),
.Y(n_1200)
);

CKINVDCx8_ASAP7_75t_R g1201 ( 
.A(n_1129),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1101),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1133),
.B(n_1066),
.Y(n_1203)
);

CKINVDCx6p67_ASAP7_75t_R g1204 ( 
.A(n_1086),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1063),
.B(n_1102),
.Y(n_1205)
);

BUFx4f_ASAP7_75t_L g1206 ( 
.A(n_1179),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1126),
.B(n_1156),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1109),
.A2(n_1102),
.B1(n_1108),
.B2(n_1142),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_1148),
.A2(n_1117),
.B1(n_1144),
.B2(n_1080),
.C(n_1120),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1101),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1112),
.B(n_1150),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1062),
.A2(n_1080),
.B1(n_1134),
.B2(n_1067),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1161),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1141),
.B(n_1110),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1153),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1171),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1161),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1067),
.B(n_1060),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1068),
.A2(n_1140),
.B(n_1081),
.C(n_1060),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1059),
.A2(n_1087),
.B(n_1075),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1121),
.B(n_1167),
.Y(n_1222)
);

OAI222xp33_ASAP7_75t_L g1223 ( 
.A1(n_1089),
.A2(n_1085),
.B1(n_1078),
.B2(n_1132),
.C1(n_1176),
.C2(n_1082),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1074),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1074),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1056),
.A2(n_1090),
.B(n_1073),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_1151),
.B(n_1130),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1138),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1065),
.B(n_1125),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1079),
.B(n_1058),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1125),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_L g1232 ( 
.A(n_1062),
.B(n_1084),
.C(n_1150),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1064),
.A2(n_1157),
.B(n_1152),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1095),
.A2(n_1051),
.B(n_1124),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1122),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1131),
.A2(n_1140),
.B(n_1091),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1052),
.B(n_1105),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1159),
.B(n_1136),
.Y(n_1238)
);

AO32x2_ASAP7_75t_L g1239 ( 
.A1(n_1088),
.A2(n_1162),
.A3(n_1127),
.B1(n_1146),
.B2(n_1136),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1077),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1100),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1083),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1146),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1083),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1123),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1114),
.A2(n_1118),
.B(n_1116),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1123),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1106),
.A2(n_1172),
.B(n_1097),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1165),
.A2(n_1135),
.B1(n_1136),
.B2(n_1104),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1162),
.A2(n_1070),
.B(n_1127),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1137),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1077),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1111),
.B(n_1139),
.Y(n_1253)
);

AO32x2_ASAP7_75t_L g1254 ( 
.A1(n_1162),
.A2(n_1127),
.A3(n_1070),
.B1(n_1137),
.B2(n_1104),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1169),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1169),
.A2(n_1053),
.B(n_1145),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_L g1257 ( 
.A1(n_1113),
.A2(n_749),
.B1(n_805),
.B2(n_1039),
.Y(n_1257)
);

AOI32xp33_ASAP7_75t_L g1258 ( 
.A1(n_1143),
.A2(n_935),
.A3(n_436),
.B1(n_732),
.B2(n_605),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1147),
.A2(n_1160),
.B(n_1099),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1133),
.B(n_769),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1074),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1161),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1054),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1126),
.B(n_1156),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1143),
.A2(n_972),
.B1(n_749),
.B2(n_605),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1140),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1054),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1054),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1154),
.B(n_1166),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1077),
.B(n_1168),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1133),
.B(n_769),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1054),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1119),
.A2(n_605),
.B(n_935),
.C(n_474),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1126),
.B(n_1156),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1053),
.A2(n_1155),
.B(n_1145),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1054),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1119),
.A2(n_605),
.B(n_749),
.Y(n_1286)
);

INVx4_ASAP7_75t_SL g1287 ( 
.A(n_1086),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1054),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1147),
.A2(n_1160),
.B(n_1099),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1054),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1119),
.A2(n_605),
.B(n_935),
.C(n_474),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1128),
.B(n_1112),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1054),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1149),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1054),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1161),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1119),
.A2(n_605),
.B(n_749),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1286),
.A2(n_1297),
.B(n_1223),
.C(n_1230),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1207),
.B(n_1268),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1287),
.B(n_1180),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1281),
.A2(n_1291),
.B(n_1197),
.C(n_1269),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1283),
.B(n_1229),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1181),
.B(n_1205),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1181),
.B(n_1219),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1287),
.B(n_1180),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1269),
.A2(n_1208),
.B(n_1260),
.C(n_1183),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1203),
.B(n_1261),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1279),
.B(n_1212),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1236),
.A2(n_1188),
.B(n_1196),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1224),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1192),
.B(n_1231),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1214),
.A2(n_1296),
.B1(n_1218),
.B2(n_1265),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1236),
.A2(n_1188),
.B(n_1196),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1217),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1258),
.A2(n_1191),
.B1(n_1182),
.B2(n_1277),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1187),
.A2(n_1226),
.B(n_1246),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1222),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1187),
.A2(n_1250),
.B(n_1234),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1185),
.A2(n_1278),
.B(n_1257),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1192),
.B(n_1263),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1292),
.B(n_1232),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1266),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1273),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1238),
.B(n_1273),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1288),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1228),
.B(n_1294),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1191),
.A2(n_1182),
.B1(n_1272),
.B2(n_1275),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1228),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1210),
.B(n_1213),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1213),
.A2(n_1184),
.B1(n_1290),
.B2(n_1285),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1195),
.B(n_1198),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1209),
.Y(n_1336)
);

AND2x6_ASAP7_75t_L g1337 ( 
.A(n_1215),
.B(n_1202),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1271),
.A2(n_1280),
.B1(n_1201),
.B2(n_1296),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1186),
.A2(n_1267),
.B(n_1284),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1242),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1237),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1270),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1193),
.B(n_1289),
.Y(n_1343)
);

AOI221x1_ASAP7_75t_SL g1344 ( 
.A1(n_1189),
.A2(n_1244),
.B1(n_1247),
.B2(n_1245),
.C(n_1255),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1214),
.A2(n_1218),
.B1(n_1265),
.B2(n_1224),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1254),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1204),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1185),
.A2(n_1278),
.B(n_1240),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_SL g1349 ( 
.A1(n_1189),
.A2(n_1252),
.B1(n_1243),
.B2(n_1193),
.C(n_1259),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1220),
.A2(n_1264),
.B(n_1225),
.C(n_1251),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1259),
.B(n_1289),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1253),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1259),
.B(n_1194),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1194),
.B(n_1249),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1240),
.A2(n_1211),
.B(n_1221),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1241),
.A2(n_1206),
.B1(n_1190),
.B2(n_1211),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1206),
.Y(n_1357)
);

AND2x2_ASAP7_75t_SL g1358 ( 
.A(n_1227),
.B(n_1235),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1227),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1248),
.B(n_1256),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1248),
.A2(n_1233),
.B(n_1239),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1239),
.B(n_1186),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1262),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1262),
.B(n_1274),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1274),
.A2(n_1276),
.B1(n_1282),
.B2(n_1284),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1276),
.A2(n_1160),
.B(n_1147),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1281),
.A2(n_1291),
.B(n_1286),
.C(n_1297),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1258),
.A2(n_1191),
.B1(n_1269),
.B2(n_1143),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1238),
.A2(n_1142),
.B(n_1140),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1203),
.B(n_1261),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1258),
.A2(n_1191),
.B1(n_1269),
.B2(n_1143),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1287),
.B(n_1180),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1222),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1287),
.B(n_1180),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1203),
.B(n_1261),
.Y(n_1377)
);

BUFx4f_ASAP7_75t_L g1378 ( 
.A(n_1204),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1203),
.B(n_1261),
.Y(n_1379)
);

OAI31xp33_ASAP7_75t_L g1380 ( 
.A1(n_1281),
.A2(n_605),
.A3(n_1291),
.B(n_805),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1381)
);

INVx5_ASAP7_75t_SL g1382 ( 
.A(n_1358),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1363),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1343),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1351),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1309),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_1367),
.B(n_1361),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1362),
.B(n_1354),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1302),
.B(n_1303),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1354),
.B(n_1346),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1353),
.B(n_1359),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1342),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1368),
.A2(n_1373),
.B1(n_1318),
.B2(n_1333),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1360),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1353),
.B(n_1366),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1327),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1380),
.A2(n_1373),
.B(n_1368),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_1322),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1320),
.B(n_1375),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1363),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1321),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1363),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1312),
.B(n_1316),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1349),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1325),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1301),
.B(n_1348),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1349),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1337),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1339),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1364),
.B(n_1326),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1319),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1328),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1336),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1302),
.B(n_1381),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1334),
.B(n_1318),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1303),
.A2(n_1381),
.B(n_1370),
.Y(n_1418)
);

BUFx4f_ASAP7_75t_SL g1419 ( 
.A(n_1331),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1332),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1314),
.B(n_1323),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1304),
.B(n_1314),
.Y(n_1422)
);

AOI222xp33_ASAP7_75t_L g1423 ( 
.A1(n_1330),
.A2(n_1323),
.B1(n_1305),
.B2(n_1341),
.C1(n_1306),
.C2(n_1377),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1335),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1340),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1306),
.B(n_1305),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1298),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1308),
.A2(n_1350),
.B(n_1369),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1347),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1299),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1408),
.A2(n_1356),
.B(n_1307),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1411),
.Y(n_1433)
);

OAI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1398),
.A2(n_1338),
.B1(n_1344),
.B2(n_1356),
.C(n_1357),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1388),
.B(n_1379),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1384),
.B(n_1352),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1388),
.B(n_1310),
.Y(n_1437)
);

OAI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1398),
.A2(n_1393),
.B(n_1423),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1394),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1385),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1399),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1395),
.B(n_1372),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1414),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.B(n_1311),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1414),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1391),
.B(n_1338),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1400),
.B(n_1300),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1391),
.B(n_1313),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1410),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1391),
.B(n_1313),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1390),
.B(n_1313),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1400),
.B(n_1374),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1433),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1438),
.A2(n_1393),
.B(n_1389),
.C(n_1406),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1438),
.A2(n_1408),
.B1(n_1423),
.B2(n_1389),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1442),
.B(n_1382),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1448),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1434),
.B(n_1427),
.C(n_1409),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1434),
.A2(n_1408),
.B1(n_1416),
.B2(n_1387),
.C(n_1427),
.Y(n_1459)
);

NOR4xp25_ASAP7_75t_SL g1460 ( 
.A(n_1441),
.B(n_1429),
.C(n_1403),
.D(n_1400),
.Y(n_1460)
);

AOI322xp5_ASAP7_75t_L g1461 ( 
.A1(n_1435),
.A2(n_1406),
.A3(n_1409),
.B1(n_1416),
.B2(n_1427),
.C1(n_1426),
.C2(n_1421),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1432),
.A2(n_1408),
.B(n_1400),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1442),
.B(n_1382),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1447),
.B(n_1412),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1448),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1443),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1442),
.B(n_1382),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1446),
.A2(n_1408),
.B1(n_1387),
.B2(n_1418),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.Y(n_1469)
);

OAI31xp33_ASAP7_75t_L g1470 ( 
.A1(n_1446),
.A2(n_1401),
.A3(n_1421),
.B(n_1426),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1447),
.A2(n_1408),
.B1(n_1387),
.B2(n_1401),
.C(n_1344),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1451),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1431),
.B(n_1418),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1446),
.A2(n_1408),
.B1(n_1387),
.B2(n_1417),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1431),
.B(n_1418),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1443),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1433),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1441),
.B(n_1382),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1443),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1440),
.Y(n_1480)
);

OAI211xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1450),
.A2(n_1422),
.B(n_1420),
.C(n_1415),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1450),
.B(n_1387),
.C(n_1447),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1435),
.A2(n_1418),
.B1(n_1424),
.B2(n_1396),
.C(n_1392),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1387),
.C(n_1392),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1452),
.A2(n_1417),
.B(n_1387),
.Y(n_1485)
);

OAI332xp33_ASAP7_75t_L g1486 ( 
.A1(n_1451),
.A2(n_1315),
.A3(n_1345),
.B1(n_1422),
.B2(n_1425),
.B3(n_1397),
.C1(n_1386),
.C2(n_1407),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1445),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1445),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1452),
.A2(n_1417),
.B(n_1400),
.Y(n_1489)
);

AO221x1_ASAP7_75t_L g1490 ( 
.A1(n_1439),
.A2(n_1430),
.B1(n_1383),
.B2(n_1402),
.C(n_1404),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1466),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_SL g1492 ( 
.A(n_1454),
.B(n_1329),
.C(n_1451),
.Y(n_1492)
);

INVx4_ASAP7_75t_SL g1493 ( 
.A(n_1464),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1489),
.A2(n_1405),
.B(n_1413),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1490),
.A2(n_1405),
.B(n_1403),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1466),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1465),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1465),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1464),
.Y(n_1499)
);

BUFx8_ASAP7_75t_L g1500 ( 
.A(n_1478),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1490),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1476),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1465),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1480),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1485),
.A2(n_1405),
.B(n_1403),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1458),
.A2(n_1452),
.B(n_1400),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1444),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1476),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1479),
.Y(n_1510)
);

INVx4_ASAP7_75t_SL g1511 ( 
.A(n_1478),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1453),
.Y(n_1512)
);

INVx4_ASAP7_75t_SL g1513 ( 
.A(n_1456),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1472),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1453),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1469),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1479),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.B(n_1456),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1477),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1487),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1463),
.B(n_1441),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1491),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1513),
.B(n_1457),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1512),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1498),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1461),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1491),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1508),
.B(n_1461),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1455),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1435),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1506),
.A2(n_1458),
.B(n_1459),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1496),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1496),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1513),
.B(n_1463),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1502),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1514),
.Y(n_1540)
);

NOR2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1371),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1514),
.A2(n_1468),
.B1(n_1471),
.B2(n_1462),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1509),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1506),
.B(n_1460),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1467),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1500),
.B(n_1419),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1512),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1419),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1509),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1503),
.B(n_1437),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1504),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1503),
.B(n_1437),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1513),
.B(n_1467),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1517),
.B(n_1475),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1497),
.B(n_1484),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1517),
.Y(n_1558)
);

OAI33xp33_ASAP7_75t_L g1559 ( 
.A1(n_1510),
.A2(n_1474),
.A3(n_1481),
.B1(n_1488),
.B2(n_1436),
.B3(n_1486),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1510),
.Y(n_1560)
);

NAND2x1_ASAP7_75t_L g1561 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1498),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1498),
.B(n_1449),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1518),
.B(n_1431),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1444),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1519),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1523),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1532),
.B(n_1497),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1558),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1535),
.Y(n_1570)
);

OAI211xp5_ASAP7_75t_L g1571 ( 
.A1(n_1534),
.A2(n_1483),
.B(n_1505),
.C(n_1501),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1528),
.B(n_1523),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1535),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1437),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1527),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1505),
.C(n_1498),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1561),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1527),
.B(n_1498),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1552),
.B(n_1497),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1449),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1561),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1526),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1537),
.B(n_1545),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1536),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1525),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1444),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1526),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1559),
.A2(n_1501),
.B(n_1505),
.C(n_1428),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1537),
.B(n_1545),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1536),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

AND2x2_ASAP7_75t_SL g1593 ( 
.A(n_1546),
.B(n_1378),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1538),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1538),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_SL g1596 ( 
.A(n_1533),
.B(n_1495),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1551),
.B(n_1500),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1500),
.Y(n_1599)
);

OAI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1542),
.A2(n_1494),
.B(n_1499),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1570),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1579),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1590),
.B(n_1533),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1592),
.B(n_1555),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1583),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1592),
.B(n_1555),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1589),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.B(n_1554),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1554),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1567),
.B(n_1556),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1574),
.B(n_1564),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1575),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1589),
.Y(n_1616)
);

NAND3xp33_ASAP7_75t_L g1617 ( 
.A(n_1576),
.B(n_1544),
.C(n_1505),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1585),
.B(n_1533),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1593),
.B(n_1511),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1566),
.B(n_1565),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1578),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1596),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1525),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1610),
.B(n_1598),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1588),
.B(n_1600),
.C(n_1571),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1619),
.B(n_1599),
.C(n_1597),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1598),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1617),
.B(n_1568),
.C(n_1575),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1602),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.B(n_1578),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1602),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1614),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1608),
.A2(n_1577),
.B(n_1581),
.C(n_1594),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1608),
.A2(n_1577),
.B(n_1581),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1614),
.Y(n_1638)
);

NAND2x1_ASAP7_75t_SL g1639 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1621),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1621),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1623),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1615),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1611),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1630),
.B(n_1603),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1639),
.Y(n_1647)
);

NAND2x1_ASAP7_75t_L g1648 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1628),
.A2(n_1616),
.B1(n_1607),
.B2(n_1605),
.C1(n_1622),
.C2(n_1625),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1627),
.B(n_1622),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1626),
.B(n_1618),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1609),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1628),
.A2(n_1623),
.B1(n_1604),
.B2(n_1618),
.C(n_1609),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1649),
.B(n_1637),
.C(n_1629),
.Y(n_1657)
);

NAND5xp2_ASAP7_75t_L g1658 ( 
.A(n_1656),
.B(n_1629),
.C(n_1636),
.D(n_1642),
.E(n_1638),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1651),
.A2(n_1604),
.B1(n_1624),
.B2(n_1623),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1650),
.A2(n_1641),
.B(n_1640),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1655),
.B(n_1635),
.C(n_1632),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1646),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1648),
.A2(n_1593),
.B(n_1634),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1651),
.A2(n_1624),
.B1(n_1612),
.B2(n_1563),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1647),
.B(n_1612),
.C(n_1591),
.Y(n_1665)
);

OAI222xp33_ASAP7_75t_L g1666 ( 
.A1(n_1653),
.A2(n_1580),
.B1(n_1563),
.B2(n_1613),
.C1(n_1595),
.C2(n_1586),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1654),
.C(n_1645),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1662),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1652),
.B1(n_1580),
.B2(n_1563),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1660),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1661),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1670),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1668),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1671),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1669),
.B(n_1663),
.C(n_1665),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1667),
.B(n_1666),
.C(n_1664),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1511),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1613),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1673),
.A2(n_1580),
.B1(n_1563),
.B2(n_1587),
.C(n_1582),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1676),
.A2(n_1587),
.B1(n_1582),
.B2(n_1378),
.C(n_1507),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1672),
.A2(n_1539),
.B(n_1543),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1679),
.Y(n_1683)
);

AND4x1_ASAP7_75t_L g1684 ( 
.A(n_1682),
.B(n_1674),
.C(n_1524),
.D(n_1529),
.Y(n_1684)
);

NOR3x1_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1507),
.C(n_1494),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_L g1686 ( 
.A(n_1683),
.B(n_1680),
.C(n_1678),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1686),
.B(n_1684),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1687),
.A2(n_1685),
.B(n_1550),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1548),
.B1(n_1547),
.B2(n_1560),
.Y(n_1689)
);

OAI31xp33_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1548),
.A3(n_1547),
.B(n_1499),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1499),
.B1(n_1493),
.B2(n_1564),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1515),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1692),
.B(n_1515),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1493),
.B1(n_1512),
.B2(n_1521),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1516),
.B1(n_1522),
.B2(n_1520),
.Y(n_1695)
);

AOI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1376),
.B(n_1518),
.C(n_1520),
.Y(n_1696)
);


endmodule