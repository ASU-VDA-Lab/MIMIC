module real_aes_7072_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_1106;
wire n_618;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_905;
wire n_635;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_792;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1070;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1135;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_598;
wire n_404;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1014;
wire n_1028;
wire n_1083;
wire n_727;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_922;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_1102;
wire n_1076;
wire n_463;
wire n_601;
wire n_804;
wire n_396;
wire n_661;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_1119;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_0), .A2(n_59), .B1(n_523), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_1), .A2(n_286), .B1(n_544), .B2(n_666), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g1102 ( .A(n_2), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_3), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_4), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_5), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_6), .A2(n_137), .B1(n_534), .B2(n_929), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_7), .Y(n_1014) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_8), .A2(n_225), .B1(n_408), .B2(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g1084 ( .A(n_8), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_9), .A2(n_158), .B1(n_630), .B2(n_802), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_10), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_11), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_12), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_13), .A2(n_290), .B1(n_499), .B2(n_500), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_14), .A2(n_105), .B1(n_630), .B2(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_15), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_16), .A2(n_52), .B1(n_149), .B2(n_427), .C1(n_761), .C2(n_762), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_17), .A2(n_54), .B1(n_621), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_18), .A2(n_254), .B1(n_902), .B2(n_903), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_19), .A2(n_155), .B1(n_510), .B2(n_594), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_20), .B(n_567), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_21), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_22), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_23), .A2(n_308), .B1(n_480), .B2(n_540), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_24), .A2(n_357), .B1(n_466), .B2(n_471), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g1133 ( .A1(n_25), .A2(n_304), .B1(n_545), .B2(n_902), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_26), .Y(n_953) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_27), .A2(n_58), .B1(n_341), .B2(n_425), .C1(n_521), .C2(n_523), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_28), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_29), .A2(n_123), .B1(n_515), .B2(n_789), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_30), .A2(n_55), .B1(n_479), .B2(n_804), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_31), .Y(n_780) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_32), .A2(n_112), .B1(n_408), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_33), .A2(n_373), .B1(n_598), .B2(n_905), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_34), .A2(n_255), .B1(n_513), .B2(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g625 ( .A(n_35), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_36), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_37), .A2(n_117), .B1(n_482), .B2(n_535), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_38), .A2(n_277), .B1(n_929), .B2(n_942), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_39), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_40), .B(n_763), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_41), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_42), .B(n_1046), .Y(n_1045) );
AOI22xp5_ASAP7_75t_SL g669 ( .A1(n_43), .A2(n_670), .B1(n_671), .B2(n_697), .Y(n_669) );
INVx1_ASAP7_75t_L g697 ( .A(n_43), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_44), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_45), .A2(n_293), .B1(n_522), .B2(n_585), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_46), .A2(n_334), .B1(n_458), .B2(n_545), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_47), .A2(n_219), .B1(n_433), .B2(n_522), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_48), .A2(n_252), .B1(n_486), .B2(n_605), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_49), .B(n_970), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_50), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_51), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_53), .A2(n_124), .B1(n_807), .B2(n_810), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g1123 ( .A1(n_56), .A2(n_77), .B1(n_763), .B2(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_57), .A2(n_378), .B1(n_813), .B2(n_999), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_60), .A2(n_145), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_61), .A2(n_250), .B1(n_902), .B2(n_903), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_62), .A2(n_287), .B1(n_476), .B2(n_480), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_63), .A2(n_108), .B1(n_539), .B2(n_541), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_64), .A2(n_914), .B1(n_934), .B2(n_935), .Y(n_913) );
INVx1_ASAP7_75t_L g934 ( .A(n_64), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_65), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_66), .A2(n_343), .B1(n_902), .B2(n_903), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_67), .A2(n_298), .B1(n_476), .B2(n_635), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_68), .Y(n_615) );
INVx1_ASAP7_75t_L g841 ( .A(n_69), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_70), .A2(n_188), .B1(n_534), .B2(n_1002), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_71), .A2(n_355), .B1(n_495), .B2(n_548), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_72), .A2(n_103), .B1(n_515), .B2(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_73), .A2(n_340), .B1(n_548), .B2(n_813), .Y(n_849) );
INVx1_ASAP7_75t_L g755 ( .A(n_74), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_75), .A2(n_98), .B1(n_466), .B2(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_76), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_78), .B(n_762), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_79), .A2(n_261), .B1(n_522), .B2(n_585), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_80), .A2(n_291), .B1(n_517), .B2(n_519), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_81), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_82), .A2(n_313), .B1(n_445), .B2(n_761), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_83), .A2(n_216), .B1(n_445), .B2(n_523), .Y(n_1042) );
INVx1_ASAP7_75t_L g938 ( .A(n_84), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_85), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_86), .A2(n_212), .B1(n_534), .B2(n_536), .Y(n_533) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_87), .A2(n_256), .B1(n_408), .B2(n_409), .Y(n_415) );
INVx1_ASAP7_75t_L g1081 ( .A(n_87), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_88), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_89), .A2(n_90), .B1(n_499), .B2(n_519), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_91), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_92), .A2(n_107), .B1(n_602), .B2(n_791), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_93), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_94), .A2(n_233), .B1(n_446), .B2(n_585), .Y(n_655) );
OA22x2_ASAP7_75t_L g704 ( .A1(n_95), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_95), .Y(n_705) );
AOI22x1_ASAP7_75t_L g881 ( .A1(n_96), .A2(n_882), .B1(n_906), .B2(n_907), .Y(n_881) );
INVx1_ASAP7_75t_L g906 ( .A(n_96), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_97), .Y(n_1020) );
INVx1_ASAP7_75t_L g1107 ( .A(n_99), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_100), .A2(n_144), .B1(n_676), .B2(n_678), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_101), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_102), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_104), .A2(n_184), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_106), .A2(n_359), .B1(n_689), .B2(n_690), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_109), .A2(n_364), .B1(n_486), .B2(n_732), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_110), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_111), .A2(n_150), .B1(n_479), .B2(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g1085 ( .A(n_112), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_113), .A2(n_165), .B1(n_509), .B2(n_595), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_114), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_115), .A2(n_133), .B1(n_549), .B2(n_1135), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_116), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_118), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_119), .A2(n_1088), .B1(n_1108), .B2(n_1109), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g1108 ( .A(n_119), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_120), .A2(n_289), .B1(n_517), .B2(n_541), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_121), .B(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_122), .A2(n_294), .B1(n_630), .B2(n_789), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_125), .A2(n_243), .B1(n_970), .B2(n_992), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_126), .A2(n_305), .B1(n_488), .B2(n_515), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_127), .A2(n_214), .B1(n_752), .B2(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_128), .A2(n_177), .B1(n_594), .B2(n_595), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_129), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_130), .A2(n_300), .B1(n_471), .B2(n_499), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_131), .A2(n_172), .B1(n_691), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_132), .A2(n_333), .B1(n_446), .B2(n_595), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_134), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_135), .A2(n_309), .B1(n_433), .B2(n_439), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_136), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_138), .A2(n_329), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g1069 ( .A1(n_139), .A2(n_227), .B1(n_314), .B2(n_427), .C1(n_680), .C2(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_140), .A2(n_310), .B1(n_902), .B2(n_903), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_141), .A2(n_200), .B1(n_458), .B2(n_461), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_142), .A2(n_207), .B1(n_802), .B2(n_944), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_143), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_146), .A2(n_245), .B1(n_482), .B2(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_147), .A2(n_205), .B1(n_732), .B2(n_942), .Y(n_1028) );
AND2x6_ASAP7_75t_L g385 ( .A(n_148), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_148), .Y(n_1078) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_151), .A2(n_169), .B1(n_519), .B2(n_996), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_152), .A2(n_175), .B1(n_517), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_153), .A2(n_265), .B1(n_564), .B2(n_791), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_154), .A2(n_279), .B1(n_549), .B2(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_156), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_157), .A2(n_263), .B1(n_460), .B2(n_695), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_159), .A2(n_186), .B1(n_461), .B2(n_1051), .Y(n_1050) );
AOI22xp5_ASAP7_75t_SL g833 ( .A1(n_160), .A2(n_834), .B1(n_853), .B2(n_854), .Y(n_833) );
INVx1_ASAP7_75t_L g854 ( .A(n_160), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_161), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_162), .A2(n_303), .B1(n_878), .B2(n_944), .Y(n_943) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_163), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g837 ( .A(n_164), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_166), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g1136 ( .A1(n_167), .A2(n_262), .B1(n_630), .B2(n_1051), .Y(n_1136) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_168), .A2(n_247), .B1(n_408), .B2(n_412), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_168), .B(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_170), .A2(n_181), .B1(n_496), .B2(n_549), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_171), .A2(n_260), .B1(n_604), .B2(n_605), .Y(n_603) );
XNOR2x2_ASAP7_75t_L g1057 ( .A(n_173), .B(n_1058), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_174), .A2(n_358), .B1(n_476), .B2(n_480), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_176), .A2(n_270), .B1(n_445), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_178), .A2(n_187), .B1(n_458), .B2(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_179), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_180), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_182), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_183), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_185), .A2(n_321), .B1(n_802), .B2(n_980), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_189), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_190), .A2(n_230), .B1(n_602), .B2(n_800), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_191), .A2(n_203), .B1(n_536), .B2(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_192), .A2(n_237), .B1(n_499), .B2(n_663), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_193), .A2(n_231), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_194), .A2(n_610), .B1(n_636), .B2(n_637), .Y(n_609) );
INVx1_ASAP7_75t_L g636 ( .A(n_194), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_195), .A2(n_361), .B1(n_495), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g674 ( .A(n_196), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_197), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_198), .A2(n_318), .B1(n_549), .B2(n_905), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_199), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_201), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_202), .A2(n_367), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_204), .A2(n_292), .B1(n_500), .B2(n_540), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g978 ( .A1(n_206), .A2(n_299), .B1(n_460), .B2(n_468), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_208), .A2(n_353), .B1(n_496), .B2(n_598), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_209), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_210), .B(n_567), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_211), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_213), .Y(n_1099) );
AOI22xp33_ASAP7_75t_SL g1131 ( .A1(n_215), .A2(n_248), .B1(n_439), .B2(n_678), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_217), .A2(n_224), .B1(n_445), .B2(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_218), .A2(n_330), .B1(n_486), .B2(n_488), .Y(n_485) );
XNOR2x2_ASAP7_75t_L g741 ( .A(n_220), .B(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_221), .A2(n_259), .B1(n_519), .B2(n_536), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_222), .A2(n_228), .B1(n_544), .B2(n_545), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_223), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_226), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_229), .A2(n_346), .B1(n_540), .B2(n_745), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_232), .A2(n_325), .B1(n_499), .B2(n_500), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_234), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_235), .A2(n_273), .B1(n_807), .B2(n_810), .Y(n_852) );
INVxp67_ASAP7_75t_L g1117 ( .A(n_236), .Y(n_1117) );
XNOR2xp5_ASAP7_75t_L g1118 ( .A(n_236), .B(n_1119), .Y(n_1118) );
OA22x2_ASAP7_75t_L g858 ( .A1(n_238), .A2(n_859), .B1(n_860), .B2(n_880), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_238), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_239), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_240), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_241), .A2(n_372), .B1(n_752), .B2(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_242), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g389 ( .A(n_244), .B(n_390), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_246), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_249), .A2(n_258), .B1(n_476), .B2(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_251), .B(n_685), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_253), .A2(n_274), .B1(n_439), .B2(n_524), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_257), .A2(n_347), .B1(n_440), .B2(n_761), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_264), .A2(n_530), .B1(n_575), .B2(n_576), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_264), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_266), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_267), .A2(n_365), .B1(n_496), .B2(n_813), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_268), .A2(n_371), .B1(n_604), .B2(n_732), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_269), .B(n_505), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_271), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_272), .Y(n_863) );
OA22x2_ASAP7_75t_L g982 ( .A1(n_275), .A2(n_983), .B1(n_984), .B2(n_1005), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_275), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_276), .B(n_592), .Y(n_756) );
INVx1_ASAP7_75t_L g840 ( .A(n_278), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_280), .A2(n_301), .B1(n_471), .B2(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g844 ( .A(n_281), .Y(n_844) );
INVx1_ASAP7_75t_L g408 ( .A(n_282), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_282), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_283), .A2(n_369), .B1(n_515), .B2(n_791), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_284), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_285), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_288), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_295), .Y(n_1033) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_296), .A2(n_383), .B(n_391), .C(n_1086), .Y(n_382) );
INVx1_ASAP7_75t_L g1098 ( .A(n_297), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_302), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_306), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_307), .A2(n_363), .B1(n_544), .B2(n_666), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_311), .A2(n_328), .B1(n_488), .B2(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g1130 ( .A(n_312), .B(n_592), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_315), .A2(n_352), .B1(n_517), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_316), .A2(n_339), .B1(n_440), .B2(n_680), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_317), .Y(n_622) );
INVx1_ASAP7_75t_L g390 ( .A(n_319), .Y(n_390) );
INVx1_ASAP7_75t_L g626 ( .A(n_320), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_322), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_323), .Y(n_606) );
INVx1_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_326), .A2(n_360), .B1(n_519), .B2(n_534), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_327), .B(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_331), .A2(n_335), .B1(n_684), .B2(n_685), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_332), .A2(n_342), .B1(n_461), .B2(n_536), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_336), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_337), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_338), .B(n_762), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_344), .Y(n_1041) );
INVx1_ASAP7_75t_L g792 ( .A(n_345), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_348), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_349), .B(n_678), .Y(n_1017) );
INVx1_ASAP7_75t_L g838 ( .A(n_350), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_351), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_354), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_356), .Y(n_562) );
INVx1_ASAP7_75t_L g668 ( .A(n_362), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_366), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_368), .B(n_445), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_370), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_374), .A2(n_794), .B1(n_826), .B2(n_827), .Y(n_793) );
INVx1_ASAP7_75t_L g826 ( .A(n_374), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_375), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_376), .Y(n_924) );
INVx1_ASAP7_75t_L g845 ( .A(n_377), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_379), .A2(n_381), .B1(n_802), .B2(n_804), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_380), .Y(n_619) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1077 ( .A(n_386), .Y(n_1077) );
OAI21xp5_ASAP7_75t_L g1115 ( .A1(n_387), .A2(n_1076), .B(n_1116), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_641), .B2(n_1072), .C(n_1073), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_526), .B1(n_639), .B2(n_640), .Y(n_393) );
INVx1_ASAP7_75t_L g639 ( .A(n_394), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_490), .Y(n_394) );
XNOR2x1_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_456), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_423), .C(n_443), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_418), .B2(n_419), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_401), .A2(n_616), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_403), .A2(n_503), .B1(n_816), .B2(n_817), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_403), .A2(n_574), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g571 ( .A(n_404), .Y(n_571) );
BUFx3_ASAP7_75t_L g614 ( .A(n_404), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_404), .A2(n_574), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_948) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_413), .Y(n_404) );
INVx2_ASAP7_75t_L g489 ( .A(n_405), .Y(n_489) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_411), .Y(n_405) );
AND2x2_ASAP7_75t_L g422 ( .A(n_406), .B(n_411), .Y(n_422) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_437), .Y(n_464) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_407), .B(n_411), .Y(n_428) );
AND2x2_ASAP7_75t_L g438 ( .A(n_407), .B(n_417), .Y(n_438) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_410), .Y(n_412) );
INVx2_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_411), .Y(n_442) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_414), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g479 ( .A(n_414), .B(n_464), .Y(n_479) );
AND2x4_ASAP7_75t_L g507 ( .A(n_414), .B(n_489), .Y(n_507) );
AND2x6_ASAP7_75t_L g589 ( .A(n_414), .B(n_422), .Y(n_589) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
INVx1_ASAP7_75t_L g436 ( .A(n_415), .Y(n_436) );
INVx1_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_415), .B(n_417), .Y(n_474) );
AND2x2_ASAP7_75t_L g429 ( .A(n_416), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g463 ( .A(n_417), .B(n_454), .Y(n_463) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g503 ( .A(n_420), .Y(n_503) );
INVx1_ASAP7_75t_L g652 ( .A(n_420), .Y(n_652) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g574 ( .A(n_421), .Y(n_574) );
AND2x4_ASAP7_75t_L g460 ( .A(n_422), .B(n_429), .Y(n_460) );
AND2x2_ASAP7_75t_L g470 ( .A(n_422), .B(n_463), .Y(n_470) );
OAI21xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_431), .B(n_432), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_424), .A2(n_674), .B(n_675), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_424), .A2(n_819), .B1(n_820), .B2(n_821), .C(n_822), .Y(n_818) );
OAI221xp5_ASAP7_75t_SL g839 ( .A1(n_424), .A2(n_563), .B1(n_840), .B2(n_841), .C(n_842), .Y(n_839) );
OAI221xp5_ASAP7_75t_SL g919 ( .A1(n_424), .A2(n_720), .B1(n_920), .B2(n_921), .C(n_922), .Y(n_919) );
OAI221xp5_ASAP7_75t_SL g1100 ( .A1(n_424), .A2(n_563), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_426), .A2(n_654), .B(n_655), .Y(n_653) );
BUFx2_ASAP7_75t_L g775 ( .A(n_426), .Y(n_775) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g561 ( .A(n_427), .Y(n_561) );
BUFx3_ASAP7_75t_L g716 ( .A(n_427), .Y(n_716) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_427), .Y(n_874) );
INVx2_ASAP7_75t_L g965 ( .A(n_427), .Y(n_965) );
AND2x6_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g451 ( .A(n_428), .Y(n_451) );
AND2x4_ASAP7_75t_L g524 ( .A(n_428), .B(n_453), .Y(n_524) );
AND2x2_ASAP7_75t_L g487 ( .A(n_429), .B(n_464), .Y(n_487) );
AND2x6_ASAP7_75t_L g488 ( .A(n_429), .B(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_433), .Y(n_621) );
INVx1_ASAP7_75t_L g1023 ( .A(n_433), .Y(n_1023) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_434), .Y(n_509) );
BUFx2_ASAP7_75t_L g564 ( .A(n_434), .Y(n_564) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_434), .Y(n_594) );
BUFx4f_ASAP7_75t_SL g761 ( .A(n_434), .Y(n_761) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g447 ( .A(n_436), .Y(n_447) );
INVx1_ASAP7_75t_L g556 ( .A(n_437), .Y(n_556) );
AND2x4_ASAP7_75t_L g440 ( .A(n_438), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g446 ( .A(n_438), .B(n_447), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_438), .B(n_556), .Y(n_555) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g510 ( .A(n_440), .Y(n_510) );
BUFx2_ASAP7_75t_L g595 ( .A(n_440), .Y(n_595) );
INVx1_ASAP7_75t_L g759 ( .A(n_440), .Y(n_759) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g473 ( .A(n_442), .B(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_448), .B1(n_449), .B2(n_455), .Y(n_443) );
INVx1_ASAP7_75t_L g1070 ( .A(n_444), .Y(n_1070) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g567 ( .A(n_445), .Y(n_567) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx12f_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_446), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_449), .A2(n_553), .B1(n_625), .B2(n_626), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_449), .A2(n_722), .B1(n_824), .B2(n_825), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_449), .A2(n_722), .B1(n_894), .B2(n_895), .Y(n_893) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g559 ( .A(n_450), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_450), .A2(n_473), .B1(n_869), .B2(n_870), .Y(n_868) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND4x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_465), .C(n_475), .D(n_485), .Y(n_456) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
INVx2_ASAP7_75t_L g544 ( .A(n_459), .Y(n_544) );
INVx2_ASAP7_75t_L g598 ( .A(n_459), .Y(n_598) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx3_ASAP7_75t_L g791 ( .A(n_460), .Y(n_791) );
BUFx3_ASAP7_75t_L g809 ( .A(n_460), .Y(n_809) );
BUFx3_ASAP7_75t_L g902 ( .A(n_460), .Y(n_902) );
INVx1_ASAP7_75t_L g811 ( .A(n_461), .Y(n_811) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g515 ( .A(n_462), .Y(n_515) );
BUFx3_ASAP7_75t_L g602 ( .A(n_462), .Y(n_602) );
BUFx3_ASAP7_75t_L g691 ( .A(n_462), .Y(n_691) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_463), .B(n_464), .Y(n_739) );
AND2x4_ASAP7_75t_L g483 ( .A(n_464), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_468), .Y(n_548) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_468), .Y(n_1135) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g497 ( .A(n_469), .Y(n_497) );
INVx3_ASAP7_75t_L g666 ( .A(n_469), .Y(n_666) );
INVx1_ASAP7_75t_L g695 ( .A(n_469), .Y(n_695) );
INVx2_ASAP7_75t_L g752 ( .A(n_469), .Y(n_752) );
INVx5_ASAP7_75t_L g878 ( .A(n_469), .Y(n_878) );
INVx8_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
BUFx4f_ASAP7_75t_SL g549 ( .A(n_472), .Y(n_549) );
BUFx2_ASAP7_75t_L g753 ( .A(n_472), .Y(n_753) );
BUFx2_ASAP7_75t_L g813 ( .A(n_472), .Y(n_813) );
INVx6_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g786 ( .A(n_473), .Y(n_786) );
INVx1_ASAP7_75t_SL g980 ( .A(n_473), .Y(n_980) );
INVx1_ASAP7_75t_L g484 ( .A(n_474), .Y(n_484) );
INVx4_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g747 ( .A(n_477), .Y(n_747) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g499 ( .A(n_479), .Y(n_499) );
BUFx3_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
INVx2_ASAP7_75t_L g803 ( .A(n_479), .Y(n_803) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_479), .Y(n_1032) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_482), .Y(n_635) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g519 ( .A(n_483), .Y(n_519) );
BUFx3_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
BUFx2_ASAP7_75t_SL g605 ( .A(n_483), .Y(n_605) );
BUFx2_ASAP7_75t_L g663 ( .A(n_483), .Y(n_663) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_483), .Y(n_732) );
AND2x2_ASAP7_75t_L g944 ( .A(n_484), .B(n_556), .Y(n_944) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g518 ( .A(n_487), .Y(n_518) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
BUFx2_ASAP7_75t_SL g604 ( .A(n_487), .Y(n_604) );
INVx11_ASAP7_75t_L g514 ( .A(n_488), .Y(n_514) );
INVx11_ASAP7_75t_L g537 ( .A(n_488), .Y(n_537) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
XNOR2x2_ASAP7_75t_L g578 ( .A(n_491), .B(n_579), .Y(n_578) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_525), .Y(n_491) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .C(n_511), .D(n_520), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OA211x2_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .C(n_508), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_503), .A2(n_614), .B1(n_863), .B2(n_864), .Y(n_862) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx5_ASAP7_75t_L g592 ( .A(n_506), .Y(n_592) );
INVx2_ASAP7_75t_L g684 ( .A(n_506), .Y(n_684) );
INVx2_ASAP7_75t_L g970 ( .A(n_506), .Y(n_970) );
INVx4_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_509), .Y(n_720) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
INVx2_ASAP7_75t_L g734 ( .A(n_513), .Y(n_734) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g745 ( .A(n_514), .Y(n_745) );
INVx5_ASAP7_75t_SL g800 ( .A(n_514), .Y(n_800) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_514), .Y(n_997) );
INVx4_ASAP7_75t_L g1051 ( .A(n_514), .Y(n_1051) );
INVx1_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g942 ( .A(n_518), .Y(n_942) );
BUFx4f_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g677 ( .A(n_522), .Y(n_677) );
BUFx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_SL g585 ( .A(n_524), .Y(n_585) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_524), .Y(n_680) );
INVx1_ASAP7_75t_L g640 ( .A(n_526), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_608), .B1(n_609), .B2(n_638), .Y(n_526) );
INVx1_ASAP7_75t_L g638 ( .A(n_527), .Y(n_638) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_577), .B1(n_578), .B2(n_607), .Y(n_528) );
INVx1_ASAP7_75t_L g607 ( .A(n_529), .Y(n_607) );
INVx1_ASAP7_75t_SL g576 ( .A(n_530), .Y(n_576) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_531), .B(n_550), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .Y(n_532) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g630 ( .A(n_535), .Y(n_630) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_535), .Y(n_750) );
INVx4_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g689 ( .A(n_537), .Y(n_689) );
INVx2_ASAP7_75t_SL g789 ( .A(n_537), .Y(n_789) );
OAI21xp33_ASAP7_75t_SL g865 ( .A1(n_537), .A2(n_866), .B(n_867), .Y(n_865) );
INVx4_ASAP7_75t_L g929 ( .A(n_537), .Y(n_929) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g1003 ( .A(n_540), .Y(n_1003) );
BUFx2_ASAP7_75t_L g804 ( .A(n_541), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR3xp33_ASAP7_75t_SL g550 ( .A(n_551), .B(n_560), .C(n_568), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_557), .B2(n_558), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_553), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_553), .A2(n_558), .B1(n_924), .B2(n_925), .Y(n_923) );
INVx3_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_555), .A2(n_620), .B1(n_657), .B2(n_658), .Y(n_656) );
BUFx3_ASAP7_75t_L g722 ( .A(n_555), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_555), .A2(n_781), .B1(n_844), .B2(n_845), .Y(n_843) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_555), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_558), .A2(n_1105), .B1(n_1106), .B2(n_1107), .Y(n_1104) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g781 ( .A(n_559), .Y(n_781) );
OAI221xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_562), .B1(n_563), .B2(n_565), .C(n_566), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g582 ( .A1(n_561), .A2(n_583), .B(n_584), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_561), .A2(n_619), .B1(n_620), .B2(n_622), .C(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_572), .B2(n_573), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_570), .A2(n_616), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g710 ( .A(n_571), .Y(n_710) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g617 ( .A(n_574), .Y(n_617) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
XOR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_606), .Y(n_579) );
NAND3x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_596), .C(n_600), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .C(n_593), .Y(n_586) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g685 ( .A(n_589), .Y(n_685) );
INVx1_ASAP7_75t_SL g993 ( .A(n_589), .Y(n_993) );
BUFx4f_ASAP7_75t_L g1046 ( .A(n_589), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g777 ( .A(n_594), .Y(n_777) );
INVx2_ASAP7_75t_L g820 ( .A(n_594), .Y(n_820) );
INVx4_ASAP7_75t_L g1125 ( .A(n_594), .Y(n_1125) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
BUFx3_ASAP7_75t_L g903 ( .A(n_602), .Y(n_903) );
INVx1_ASAP7_75t_L g729 ( .A(n_604), .Y(n_729) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g637 ( .A(n_610), .Y(n_637) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_611), .B(n_627), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_618), .C(n_624), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_614), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
OAI22xp5_ASAP7_75t_SL g709 ( .A1(n_616), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_616), .A2(n_710), .B1(n_917), .B2(n_918), .Y(n_916) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g1072 ( .A(n_641), .Y(n_1072) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_830), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_699), .B2(n_829), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OA22x2_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_669), .B2(n_698), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g766 ( .A(n_646), .B(n_767), .Y(n_766) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_668), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_659), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .C(n_656), .Y(n_648) );
OA211x2_ASAP7_75t_L g754 ( .A1(n_652), .A2(n_755), .B(n_756), .C(n_757), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_652), .A2(n_710), .B1(n_837), .B2(n_838), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_652), .A2(n_710), .B1(n_885), .B2(n_886), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g698 ( .A(n_669), .Y(n_698) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_672), .B(n_686), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_681), .Y(n_672) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_693), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .Y(n_687) );
BUFx4f_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g829 ( .A(n_699), .Y(n_829) );
XOR2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_764), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_740), .B2(n_741), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_723), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_713), .C(n_718), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_717), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g952 ( .A1(n_715), .A2(n_953), .B(n_954), .Y(n_952) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_722), .A2(n_1022), .B1(n_1023), .B2(n_1024), .Y(n_1021) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .C(n_733), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND4xp75_ASAP7_75t_L g742 ( .A(n_743), .B(n_748), .C(n_754), .D(n_760), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_752), .Y(n_999) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g1065 ( .A(n_759), .Y(n_1065) );
INVx1_ASAP7_75t_L g890 ( .A(n_761), .Y(n_890) );
BUFx4f_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g1015 ( .A(n_763), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_793), .B2(n_828), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_792), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_782), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_773), .C(n_778), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_776), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g828 ( .A(n_793), .Y(n_828) );
INVx2_ASAP7_75t_L g827 ( .A(n_794), .Y(n_827) );
AND2x2_ASAP7_75t_SL g794 ( .A(n_795), .B(n_814), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_805), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_812), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .C(n_823), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_958), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_855), .B1(n_956), .B2(n_957), .Y(n_831) );
INVxp67_ASAP7_75t_L g956 ( .A(n_832), .Y(n_956) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_SL g853 ( .A(n_834), .Y(n_853) );
AND2x2_ASAP7_75t_SL g834 ( .A(n_835), .B(n_846), .Y(n_834) );
NOR3xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_839), .C(n_843), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_850), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g957 ( .A(n_855), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_910), .B1(n_911), .B2(n_955), .Y(n_855) );
INVx1_ASAP7_75t_L g955 ( .A(n_856), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_881), .B1(n_908), .B2(n_909), .Y(n_856) );
INVx1_ASAP7_75t_L g908 ( .A(n_857), .Y(n_908) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g880 ( .A(n_860), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_871), .Y(n_860) );
NOR3xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_865), .C(n_868), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_876), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_875), .Y(n_872) );
INVx2_ASAP7_75t_SL g888 ( .A(n_874), .Y(n_888) );
INVx2_ASAP7_75t_L g1013 ( .A(n_874), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_878), .Y(n_905) );
INVx2_ASAP7_75t_L g909 ( .A(n_881), .Y(n_909) );
INVx2_ASAP7_75t_SL g907 ( .A(n_882), .Y(n_907) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_896), .Y(n_882) );
NOR3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_887), .C(n_893), .Y(n_883) );
OAI221xp5_ASAP7_75t_SL g887 ( .A1(n_888), .A2(n_889), .B1(n_890), .B2(n_891), .C(n_892), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .Y(n_900) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OAI22xp5_ASAP7_75t_SL g911 ( .A1(n_912), .A2(n_913), .B1(n_936), .B2(n_937), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g935 ( .A(n_914), .Y(n_935) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_926), .Y(n_914) );
NOR3xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_919), .C(n_923), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_931), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_930), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .Y(n_931) );
INVx2_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
XNOR2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
NOR4xp75_ASAP7_75t_L g939 ( .A(n_940), .B(n_945), .C(n_948), .D(n_952), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g940 ( .A(n_941), .B(n_943), .Y(n_940) );
NAND2xp5_ASAP7_75t_SL g945 ( .A(n_946), .B(n_947), .Y(n_945) );
XNOR2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_1007), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_982), .B2(n_1006), .Y(n_959) );
INVx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_981), .Y(n_961) );
NAND2x1_ASAP7_75t_SL g962 ( .A(n_963), .B(n_973), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_968), .Y(n_963) );
OAI21xp5_ASAP7_75t_SL g964 ( .A1(n_965), .A2(n_966), .B(n_967), .Y(n_964) );
OAI21xp5_ASAP7_75t_SL g986 ( .A1(n_965), .A2(n_987), .B(n_988), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g968 ( .A(n_969), .B(n_971), .C(n_972), .Y(n_968) );
NOR2x1_ASAP7_75t_L g973 ( .A(n_974), .B(n_977), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g1006 ( .A(n_982), .Y(n_1006) );
INVx1_ASAP7_75t_SL g1005 ( .A(n_984), .Y(n_1005) );
NAND3x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_994), .C(n_1000), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
INVx1_ASAP7_75t_SL g992 ( .A(n_993), .Y(n_992) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_998), .Y(n_994) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .Y(n_1000) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B1(n_1034), .B2(n_1035), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
XOR2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1033), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1025), .Y(n_1010) );
NOR3xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1018), .C(n_1021), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .B1(n_1015), .B2(n_1016), .C(n_1017), .Y(n_1012) );
OAI21xp5_ASAP7_75t_L g1040 ( .A1(n_1013), .A2(n_1041), .B(n_1042), .Y(n_1040) );
OAI21xp5_ASAP7_75t_SL g1121 ( .A1(n_1013), .A2(n_1122), .B(n_1123), .Y(n_1121) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1029), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
INVx1_ASAP7_75t_SL g1034 ( .A(n_1035), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1057), .B2(n_1071), .Y(n_1035) );
INVx3_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
XOR2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1056), .Y(n_1037) );
NAND2xp5_ASAP7_75t_SL g1038 ( .A(n_1039), .B(n_1048), .Y(n_1038) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .C(n_1047), .Y(n_1043) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1046), .Y(n_1129) );
NOR2x1_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1053), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1052), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1057), .Y(n_1071) );
NAND4xp75_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1062), .C(n_1066), .D(n_1069), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
AND2x2_ASAP7_75t_SL g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
INVx1_ASAP7_75t_SL g1073 ( .A(n_1074), .Y(n_1073) );
NOR2x1_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1079), .Y(n_1074) );
OR2x2_ASAP7_75t_SL g1140 ( .A(n_1075), .B(n_1080), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1078), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g1111 ( .A(n_1076), .Y(n_1111) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1077), .B(n_1113), .Y(n_1116) );
CKINVDCx16_ASAP7_75t_R g1113 ( .A(n_1078), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_1080), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
OAI322xp33_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1110), .A3(n_1112), .B1(n_1114), .B2(n_1117), .C1(n_1118), .C2(n_1138), .Y(n_1086) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1088), .Y(n_1109) );
AND2x2_ASAP7_75t_SL g1088 ( .A(n_1089), .B(n_1096), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1093), .Y(n_1089) );
NAND2xp33_ASAP7_75t_SL g1090 ( .A(n_1091), .B(n_1092), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
NOR3xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1100), .C(n_1104), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_1115), .Y(n_1114) );
NAND4xp75_ASAP7_75t_SL g1119 ( .A(n_1120), .B(n_1132), .C(n_1136), .D(n_1137), .Y(n_1119) );
NOR2xp67_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1126), .Y(n_1120) );
INVx3_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1130), .C(n_1131), .Y(n_1126) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1134), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g1138 ( .A(n_1139), .Y(n_1138) );
CKINVDCx20_ASAP7_75t_R g1139 ( .A(n_1140), .Y(n_1139) );
endmodule