module real_jpeg_19267_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_41),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_1),
.B(n_101),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_10),
.B(n_23),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_145),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_1),
.A2(n_39),
.B(n_43),
.C(n_225),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_2),
.A2(n_34),
.B1(n_72),
.B2(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_72),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_3),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_106),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_106),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_189),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_9),
.B(n_72),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_22),
.B(n_31),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_10),
.B(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_130),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_129),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_109),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_109),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_81),
.B2(n_108),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_52),
.B1(n_79),
.B2(n_80),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_37),
.B(n_51),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_21),
.B(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_22),
.B(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_56),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_24),
.A2(n_27),
.B(n_30),
.C(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_26),
.B(n_35),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_26),
.Y(n_141)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_30),
.B(n_90),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_30),
.B(n_56),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_30),
.A2(n_31),
.B(n_44),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_32),
.A2(n_63),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_32),
.B(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_35),
.B(n_197),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_45),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_42),
.B(n_43),
.C(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_39),
.B(n_71),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_40),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_42),
.B(n_50),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_42),
.A2(n_47),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_42),
.Y(n_145)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_45),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_47),
.B(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_54),
.A2(n_61),
.B1(n_66),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_54),
.A2(n_66),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_54),
.B(n_224),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B(n_60),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_55),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_56),
.A2(n_86),
.B(n_118),
.Y(n_167)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_58),
.B(n_88),
.Y(n_119)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_61),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_62),
.A2(n_90),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_64),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_69),
.B(n_75),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_105),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_76),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.C(n_97),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_83),
.B(n_89),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_84),
.B(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_85),
.B(n_87),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_86),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_87),
.B(n_189),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_95),
.B(n_144),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_145),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_113),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_115),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_125),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_116),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_125),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_268),
.B(n_273),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_180),
.B(n_256),
.C(n_267),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_169),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_133),
.B(n_169),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_147),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_135),
.B(n_136),
.C(n_147),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_142),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_159),
.B1(n_160),
.B2(n_168),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_158),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_149),
.B(n_158),
.C(n_159),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2x1_ASAP7_75t_R g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_175),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_255),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_249),
.B(n_254),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_235),
.B(n_248),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_220),
.B(n_234),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_209),
.B(n_219),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_198),
.B(n_208),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_190),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_222),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_227),
.B1(n_228),
.B2(n_233),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_244),
.C(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);


endmodule