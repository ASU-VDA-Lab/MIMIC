module fake_jpeg_20451_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_50),
.B1(n_44),
.B2(n_51),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_35),
.B(n_27),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_21),
.B1(n_29),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_26),
.B1(n_32),
.B2(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_98),
.B1(n_65),
.B2(n_54),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_73),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_46),
.B1(n_51),
.B2(n_41),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_88),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_50),
.B1(n_44),
.B2(n_47),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_84),
.B1(n_87),
.B2(n_85),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_81),
.C(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_27),
.B(n_35),
.C(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_46),
.B1(n_41),
.B2(n_40),
.Y(n_84)
);

NAND2x1_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_36),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_36),
.B1(n_47),
.B2(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_94),
.Y(n_125)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_30),
.B1(n_28),
.B2(n_43),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_70),
.B(n_85),
.C(n_89),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_103),
.B(n_39),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_42),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_74),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_121),
.B1(n_126),
.B2(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_76),
.B(n_62),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_43),
.B1(n_52),
.B2(n_62),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_95),
.B1(n_96),
.B2(n_77),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_81),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_133),
.C(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_91),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_144),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_81),
.CI(n_83),
.CON(n_131),
.SN(n_131)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_132),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_138),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_71),
.B(n_73),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_137),
.B(n_143),
.Y(n_159)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_92),
.B(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_142),
.B1(n_48),
.B2(n_45),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_42),
.C(n_94),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_103),
.C(n_117),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_82),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_111),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_37),
.B(n_39),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_143),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_90),
.B1(n_78),
.B2(n_48),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_122),
.B1(n_105),
.B2(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_20),
.C(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_118),
.B(n_112),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_108),
.B1(n_111),
.B2(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_164),
.B1(n_168),
.B2(n_137),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_161),
.B(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_167),
.B1(n_173),
.B2(n_147),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_79),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_105),
.B1(n_107),
.B2(n_112),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_116),
.B1(n_39),
.B2(n_45),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_37),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_135),
.B1(n_129),
.B2(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_45),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_167),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_127),
.C(n_133),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_200),
.C(n_201),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_175),
.B1(n_156),
.B2(n_181),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_168),
.B1(n_155),
.B2(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_141),
.B1(n_131),
.B2(n_150),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_138),
.B1(n_48),
.B2(n_9),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_196),
.B1(n_180),
.B2(n_165),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_0),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_7),
.C(n_14),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_7),
.C(n_14),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_6),
.C(n_13),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.C(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_15),
.C(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_0),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_161),
.B(n_178),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_211),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_220),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_159),
.B(n_161),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_159),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.C(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_160),
.C(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_199),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_192),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_176),
.B(n_158),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_171),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_196),
.B1(n_197),
.B2(n_208),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_229),
.B1(n_232),
.B2(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_183),
.B1(n_195),
.B2(n_182),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_215),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_234),
.Y(n_250)
);

AO22x2_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_185),
.B1(n_186),
.B2(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_202),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_240),
.Y(n_245)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_212),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_226),
.B1(n_218),
.B2(n_242),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_249),
.B1(n_252),
.B2(n_245),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_233),
.B1(n_211),
.B2(n_239),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_254),
.C(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_209),
.C(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_198),
.B1(n_232),
.B2(n_231),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_204),
.C(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_231),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_261),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_253),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_265),
.Y(n_277)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_206),
.B1(n_223),
.B2(n_204),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_275),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_243),
.C(n_254),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_11),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_11),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_278),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_263),
.B(n_269),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_284),
.B(n_274),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_266),
.C(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_271),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_287),
.B(n_285),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.C(n_278),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_12),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_12),
.B(n_2),
.Y(n_300)
);


endmodule