module fake_jpeg_24559_n_282 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_38),
.B1(n_25),
.B2(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_32),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_49),
.Y(n_79)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_53),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_50),
.B1(n_38),
.B2(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_27),
.B1(n_32),
.B2(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_18),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_22),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_84),
.B1(n_90),
.B2(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_61),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_78),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_30),
.B(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_53),
.B1(n_20),
.B2(n_24),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_19),
.C(n_30),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_17),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_38),
.B1(n_35),
.B2(n_19),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_85),
.B1(n_51),
.B2(n_55),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_82),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_40),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_22),
.B1(n_16),
.B2(n_26),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_105),
.B1(n_117),
.B2(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_118),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_53),
.B1(n_51),
.B2(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_65),
.B1(n_59),
.B2(n_78),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_90),
.B1(n_88),
.B2(n_81),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_16),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_62),
.Y(n_124)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_114),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_16),
.B(n_17),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_116),
.B(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_48),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_87),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_60),
.A2(n_17),
.B(n_24),
.C(n_28),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_17),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_123),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_128),
.B(n_137),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_127),
.B1(n_131),
.B2(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_80),
.C(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_132),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_73),
.B(n_83),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_74),
.B1(n_62),
.B2(n_75),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_138),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_R g137 ( 
.A(n_109),
.B(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_77),
.B1(n_82),
.B2(n_29),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_95),
.B1(n_101),
.B2(n_116),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_21),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_17),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_65),
.B(n_71),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_144),
.B(n_128),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_98),
.A2(n_71),
.B(n_2),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_15),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_102),
.C(n_103),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_124),
.C(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_109),
.B(n_106),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_171),
.B(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_168),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OR2x4_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_95),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_129),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_100),
.B(n_91),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_3),
.B(n_4),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_1),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_122),
.A2(n_108),
.B1(n_15),
.B2(n_4),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_127),
.B1(n_139),
.B2(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_188),
.C(n_190),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_125),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_197),
.B(n_200),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_199),
.B(n_150),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_131),
.C(n_126),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_141),
.B1(n_136),
.B2(n_119),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_165),
.B1(n_152),
.B2(n_176),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_132),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_14),
.C(n_3),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_196),
.C(n_158),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_163),
.B(n_14),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_160),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_157),
.B(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_219),
.C(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_164),
.B(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_215),
.Y(n_234)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_149),
.C(n_173),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.C(n_183),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_152),
.C(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_224),
.C(n_229),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_231),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_190),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_223),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_196),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_177),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_235),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_180),
.C(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_191),
.B1(n_210),
.B2(n_206),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_243),
.B1(n_245),
.B2(n_168),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_211),
.B1(n_184),
.B2(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_204),
.B1(n_180),
.B2(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_203),
.B1(n_214),
.B2(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_189),
.B1(n_178),
.B2(n_161),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_228),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_235),
.B(n_200),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_243),
.C(n_220),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_169),
.C(n_150),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_170),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_257),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_265),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_239),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.C(n_266),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_209),
.C(n_248),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_255),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_272),
.B(n_5),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_161),
.B1(n_170),
.B2(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_276),
.Y(n_278)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_7),
.B(n_8),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_9),
.B(n_12),
.Y(n_277)
);

OA21x2_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_7),
.B(n_9),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_273),
.C(n_12),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_278),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_9),
.B(n_12),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_13),
.Y(n_282)
);


endmodule