module fake_jpeg_14413_n_401 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_47),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_58),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_72),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_12),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_88),
.Y(n_100)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_0),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_43),
.B(n_0),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_30),
.B1(n_41),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_102),
.B1(n_116),
.B2(n_126),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_43),
.B1(n_46),
.B2(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_107),
.B(n_119),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_54),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_41),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_19),
.B1(n_16),
.B2(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_138),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_85),
.B1(n_92),
.B2(n_87),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_134),
.B1(n_102),
.B2(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_36),
.Y(n_156)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_103),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_160),
.B1(n_183),
.B2(n_136),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_156),
.B(n_166),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_130),
.Y(n_157)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_58),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_174),
.C(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_16),
.B1(n_19),
.B2(n_84),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_168),
.Y(n_203)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_98),
.B(n_38),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_167),
.B(n_169),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_35),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_38),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_35),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_180),
.B(n_182),
.Y(n_212)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_206)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_116),
.A2(n_74),
.B1(n_86),
.B2(n_83),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_32),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_189),
.B1(n_120),
.B2(n_105),
.Y(n_209)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_175),
.B1(n_180),
.B2(n_124),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_137),
.B1(n_97),
.B2(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_199),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_109),
.B1(n_112),
.B2(n_96),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_222),
.B1(n_188),
.B2(n_184),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_47),
.B(n_32),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_25),
.B(n_39),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_110),
.B1(n_123),
.B2(n_115),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_64),
.B1(n_68),
.B2(n_82),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_61),
.C(n_135),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_154),
.C(n_187),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_163),
.A2(n_137),
.B1(n_122),
.B2(n_57),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_150),
.A2(n_152),
.B1(n_149),
.B2(n_157),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g222 ( 
.A1(n_164),
.A2(n_113),
.B1(n_135),
.B2(n_93),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_230),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_171),
.B1(n_170),
.B2(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_233),
.C(n_247),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_199),
.C(n_203),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_172),
.A3(n_173),
.B1(n_162),
.B2(n_181),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_170),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_198),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_214),
.B1(n_216),
.B2(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_179),
.B1(n_189),
.B2(n_154),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_246),
.Y(n_257)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_25),
.B(n_21),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_196),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_253),
.Y(n_276)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_46),
.B1(n_165),
.B2(n_158),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_250),
.B1(n_24),
.B2(n_200),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_21),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_24),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_196),
.C(n_28),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_192),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_40),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_201),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_261),
.C(n_262),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_201),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_211),
.B1(n_222),
.B2(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_231),
.B(n_211),
.C(n_206),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_240),
.B(n_246),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_198),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_225),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_275),
.B1(n_281),
.B2(n_44),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_200),
.B1(n_28),
.B2(n_40),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_249),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_220),
.B1(n_215),
.B2(n_36),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_232),
.B1(n_236),
.B2(n_227),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_284),
.B1(n_291),
.B2(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_234),
.B1(n_226),
.B2(n_240),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_243),
.B(n_226),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_286),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_241),
.B(n_238),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_266),
.C(n_278),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_274),
.B1(n_256),
.B2(n_261),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_255),
.A2(n_239),
.B1(n_237),
.B2(n_246),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_293),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_258),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_250),
.B1(n_244),
.B2(n_220),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_296),
.B1(n_300),
.B2(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_259),
.A2(n_73),
.B1(n_44),
.B2(n_182),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_257),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_257),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_266),
.A2(n_1),
.B(n_2),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_1),
.B(n_2),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_262),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_291),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_316),
.Y(n_329)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_311),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_283),
.A2(n_258),
.B1(n_276),
.B2(n_266),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_320),
.B1(n_326),
.B2(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_3),
.C(n_4),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_327),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_280),
.C(n_44),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_285),
.C(n_288),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_283),
.A2(n_280),
.B1(n_44),
.B2(n_7),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_289),
.B(n_5),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_322),
.A2(n_294),
.B1(n_293),
.B2(n_298),
.Y(n_340)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_312),
.A2(n_321),
.B1(n_306),
.B2(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_340),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_342),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_306),
.A2(n_287),
.B(n_286),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_323),
.B(n_307),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_296),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_285),
.C(n_289),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_339),
.C(n_309),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_305),
.C(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_341),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_312),
.B(n_282),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_314),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_350),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_313),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_337),
.C(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_351),
.B(n_352),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_311),
.C(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_317),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_356),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_336),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_321),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_284),
.C(n_320),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_303),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_325),
.C(n_338),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_347),
.C(n_350),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_367),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_346),
.A2(n_341),
.B1(n_343),
.B2(n_336),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_363),
.A2(n_366),
.B1(n_355),
.B2(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_365),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_343),
.B1(n_345),
.B2(n_307),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_342),
.C(n_335),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_353),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_368),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_370),
.B(n_316),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_374),
.B(n_376),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_358),
.C(n_335),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_377),
.A2(n_379),
.B(n_367),
.Y(n_384)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_378),
.A2(n_310),
.B1(n_315),
.B2(n_365),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_328),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_384),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_R g383 ( 
.A(n_375),
.B(n_360),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_383),
.A2(n_375),
.B(n_373),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_386),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_377),
.A2(n_369),
.B1(n_326),
.B2(n_300),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_371),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_391),
.Y(n_394)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_380),
.A2(n_301),
.B(n_8),
.C(n_9),
.Y(n_391)
);

AOI21x1_ASAP7_75t_L g392 ( 
.A1(n_390),
.A2(n_380),
.B(n_381),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_393),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_SL g397 ( 
.A(n_396),
.B(n_387),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_397),
.A2(n_394),
.B(n_395),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_391),
.B(n_6),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_399),
.B(n_6),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_8),
.Y(n_401)
);


endmodule