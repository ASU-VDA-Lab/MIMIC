module real_jpeg_20833_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_57;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_50;
wire n_29;
wire n_55;
wire n_58;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_49;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_60;
wire n_28;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_32;
wire n_16;
wire n_15;
wire n_13;

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_16),
.B1(n_17),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_21),
.B(n_33),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_43),
.B(n_45),
.C(n_46),
.D(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_43),
.Y(n_45)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_16),
.B1(n_17),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_24),
.B1(n_43),
.B2(n_44),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_5),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_38),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_31),
.B(n_37),
.Y(n_9)
);

NOR2xp67_ASAP7_75t_R g10 ( 
.A(n_11),
.B(n_25),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_11),
.B(n_25),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_15),
.B(n_19),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_28),
.Y(n_51)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2x1_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_28),
.B(n_44),
.C(n_47),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_61),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_55),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_55),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);


endmodule