module fake_jpeg_13484_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NAND4xp25_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_47),
.C(n_66),
.D(n_69),
.Y(n_89)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_71),
.Y(n_96)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_64),
.B1(n_57),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_94),
.B1(n_60),
.B2(n_55),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_93),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_53),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.C(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_52),
.B1(n_57),
.B2(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_71),
.C(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_107),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_110),
.B1(n_24),
.B2(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_117),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_75),
.B1(n_97),
.B2(n_62),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_55),
.B1(n_59),
.B2(n_54),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_68),
.B(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_75),
.B1(n_61),
.B2(n_67),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_118),
.C(n_10),
.Y(n_140)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_7),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_0),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_116),
.B(n_21),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_75),
.Y(n_117)
);

OA22x2_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_28),
.B1(n_45),
.B2(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_125),
.B1(n_138),
.B2(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_132),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_2),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_140),
.B(n_118),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_123),
.B(n_122),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_30),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_131),
.C(n_103),
.Y(n_142)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_29),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_139),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_128),
.B1(n_32),
.B2(n_33),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_118),
.C(n_36),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_131),
.C(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_11),
.B(n_12),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_136),
.B1(n_137),
.B2(n_134),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_40),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_14),
.B(n_140),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_149),
.C(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_157),
.B(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_163),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_154),
.A3(n_160),
.B1(n_143),
.B2(n_159),
.C1(n_158),
.C2(n_141),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_18),
.B(n_38),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_41),
.Y(n_169)
);


endmodule