module fake_aes_8647_n_1533 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1533);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1533;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_659;
wire n_386;
wire n_432;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1460;
wire n_1372;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx2_ASAP7_75t_L g331 ( .A(n_329), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_157), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_308), .Y(n_333) );
CKINVDCx14_ASAP7_75t_R g334 ( .A(n_226), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_264), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_113), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_134), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_251), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_104), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_244), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_267), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_325), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_137), .B(n_236), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_173), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_5), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_130), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_90), .Y(n_348) );
BUFx10_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_240), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_301), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_237), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_200), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_161), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_122), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_272), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_103), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_277), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_190), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_14), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_317), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_180), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_250), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_242), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_14), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_169), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_2), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_208), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_261), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_252), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_168), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_80), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_87), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_159), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_268), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_166), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_0), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_150), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_163), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_123), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_270), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_313), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_167), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_199), .Y(n_384) );
BUFx10_ASAP7_75t_L g385 ( .A(n_279), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_217), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_177), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_143), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_212), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_139), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_69), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_160), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_145), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_51), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_266), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_230), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_278), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_100), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_110), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_233), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_289), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_263), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_30), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_113), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_147), .Y(n_405) );
INVxp33_ASAP7_75t_L g406 ( .A(n_256), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_315), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_158), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_296), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_99), .Y(n_410) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_214), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_172), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_140), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_219), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_104), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_148), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_295), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_262), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_203), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_5), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_231), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_184), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_94), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_174), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_99), .Y(n_425) );
INVxp33_ASAP7_75t_SL g426 ( .A(n_165), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_291), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_207), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_307), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_80), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_114), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_229), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_171), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_9), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_45), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_117), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_324), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_222), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_245), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_58), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_186), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_98), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_243), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_70), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_192), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_93), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_211), .Y(n_447) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_151), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_101), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_282), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_293), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_202), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_35), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_6), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_11), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_239), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_311), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_204), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_187), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_56), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_292), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_40), .Y(n_462) );
NOR2xp67_ASAP7_75t_L g463 ( .A(n_55), .B(n_300), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_213), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_116), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_37), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_64), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_58), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_152), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_33), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_78), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_195), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_305), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_107), .Y(n_474) );
INVxp33_ASAP7_75t_L g475 ( .A(n_238), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_273), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_51), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_52), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_176), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_75), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_249), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_304), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_223), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_2), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_154), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_4), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_59), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_56), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_95), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_95), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_81), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_255), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_1), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_188), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_144), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_146), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_43), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_19), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_297), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_326), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_122), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_73), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_218), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_73), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_125), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_142), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_281), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_153), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_27), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_118), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_93), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_33), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_283), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_141), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_319), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_38), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_314), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_246), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_149), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_67), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_120), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_179), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_175), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_162), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_287), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_74), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_155), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_354), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_349), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_339), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_354), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_398), .Y(n_532) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_331), .A2(n_126), .B(n_124), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_440), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_373), .B(n_0), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_383), .B(n_1), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_354), .Y(n_537) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_373), .B(n_3), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_354), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_491), .B(n_3), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_388), .Y(n_541) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_331), .A2(n_128), .B(n_127), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_349), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_497), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_388), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_388), .Y(n_546) );
INVx5_ASAP7_75t_L g547 ( .A(n_388), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_377), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_474), .B(n_4), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_366), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_349), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_398), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_415), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_474), .B(n_7), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_415), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_338), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_377), .B(n_7), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_338), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_340), .B(n_8), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_402), .B(n_8), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_452), .Y(n_562) );
NAND2xp33_ASAP7_75t_L g563 ( .A(n_406), .B(n_129), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_452), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_343), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_452), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_434), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_435), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_465), .A2(n_13), .B1(n_10), .B2(n_12), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_452), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_434), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_531), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_555), .B(n_409), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_550), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_535), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_531), .Y(n_577) );
INVxp33_ASAP7_75t_L g578 ( .A(n_548), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_557), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_530), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_535), .A2(n_346), .B1(n_360), .B2(n_357), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_535), .B(n_343), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
BUFx10_ASAP7_75t_L g584 ( .A(n_535), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_549), .B(n_361), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_531), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_559), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_531), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_559), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_565), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_549), .B(n_361), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_543), .B(n_551), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_558), .A2(n_358), .B1(n_381), .B2(n_351), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_545), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_549), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_545), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_530), .B(n_534), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_554), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_545), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_543), .B(n_382), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_534), .B(n_406), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_565), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_543), .B(n_445), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_544), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_543), .B(n_551), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
INVx4_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
INVxp33_ASAP7_75t_L g612 ( .A(n_558), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_532), .A2(n_367), .B1(n_380), .B2(n_372), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_582), .A2(n_563), .B(n_533), .Y(n_614) );
INVx4_ASAP7_75t_L g615 ( .A(n_610), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_610), .B(n_551), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_578), .B(n_603), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_603), .B(n_529), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_606), .B(n_529), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_610), .A2(n_538), .B1(n_551), .B2(n_560), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_584), .B(n_376), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_610), .B(n_561), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_584), .B(n_447), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_584), .B(n_495), .Y(n_624) );
INVx4_ASAP7_75t_L g625 ( .A(n_610), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_606), .B(n_475), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_575), .A2(n_538), .B1(n_540), .B2(n_426), .Y(n_627) );
BUFx6f_ASAP7_75t_SL g628 ( .A(n_584), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_593), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_612), .B(n_426), .Y(n_630) );
NAND2xp33_ASAP7_75t_L g631 ( .A(n_609), .B(n_370), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_575), .A2(n_487), .B1(n_536), .B2(n_334), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_593), .Y(n_633) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_575), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_608), .B(n_475), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_608), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_579), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_580), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
OAI22xp5_ASAP7_75t_SL g640 ( .A1(n_595), .A2(n_486), .B1(n_490), .B2(n_470), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_604), .B(n_370), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_583), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_604), .B(n_352), .Y(n_643) );
OA22x2_ASAP7_75t_L g644 ( .A1(n_595), .A2(n_568), .B1(n_569), .B2(n_580), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_604), .B(n_464), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_573), .B(n_494), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_573), .B(n_494), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_599), .B(n_385), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_583), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_581), .B(n_334), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_599), .B(n_385), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_581), .B(n_609), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_599), .B(n_385), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_607), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_576), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_588), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_611), .B(n_532), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g658 ( .A(n_574), .B(n_569), .C(n_568), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_588), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_613), .B(n_493), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_590), .Y(n_661) );
AND2x6_ASAP7_75t_SL g662 ( .A(n_590), .B(n_399), .Y(n_662) );
NAND2x1_ASAP7_75t_L g663 ( .A(n_575), .B(n_542), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_586), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_586), .B(n_552), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_576), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_591), .Y(n_667) );
BUFx3_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_605), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_586), .B(n_571), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_605), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_613), .A2(n_351), .B1(n_381), .B2(n_358), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_597), .B(n_347), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_597), .A2(n_403), .B1(n_420), .B2(n_404), .Y(n_674) );
AOI22x1_ASAP7_75t_L g675 ( .A1(n_597), .A2(n_400), .B1(n_414), .B2(n_395), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_601), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_601), .B(n_542), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_582), .B(n_552), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_601), .A2(n_418), .B1(n_500), .B2(n_416), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_601), .B(n_416), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_585), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_585), .Y(n_682) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_592), .B(n_553), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_592), .B(n_345), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_572), .B(n_418), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_572), .A2(n_500), .B1(n_493), .B2(n_355), .Y(n_686) );
BUFx5_ASAP7_75t_L g687 ( .A(n_598), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_577), .B(n_336), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_577), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_577), .A2(n_486), .B1(n_490), .B2(n_470), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_587), .B(n_542), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_587), .B(n_391), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_587), .B(n_553), .Y(n_693) );
OR2x6_ASAP7_75t_L g694 ( .A(n_589), .B(n_411), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_589), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_598), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_602), .B(n_556), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_598), .B(n_353), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_617), .A2(n_410), .B(n_394), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_669), .Y(n_700) );
AOI21x1_ASAP7_75t_L g701 ( .A1(n_663), .A2(n_542), .B(n_344), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_626), .B(n_460), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_615), .B(n_356), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_629), .B(n_431), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_618), .A2(n_425), .B(n_430), .C(n_423), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_677), .A2(n_333), .B(n_332), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_633), .B(n_442), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_652), .A2(n_436), .B(n_455), .C(n_446), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_664), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_677), .A2(n_337), .B(n_335), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_614), .A2(n_342), .B(n_341), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_691), .A2(n_362), .B(n_350), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_615), .B(n_359), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_636), .B(n_444), .Y(n_714) );
INVx6_ASAP7_75t_L g715 ( .A(n_662), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_664), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_619), .A2(n_466), .B(n_471), .C(n_468), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_658), .B(n_651), .C(n_648), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_691), .A2(n_369), .B(n_363), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_668), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_638), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_685), .A2(n_511), .B1(n_520), .B2(n_504), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_SL g723 ( .A1(n_673), .A2(n_379), .B(n_384), .C(n_374), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_685), .A2(n_511), .B1(n_520), .B2(n_504), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_680), .A2(n_480), .B1(n_488), .B2(n_478), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_622), .A2(n_393), .B(n_392), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_672), .A2(n_449), .B1(n_454), .B2(n_453), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_641), .B(n_462), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_644), .A2(n_502), .B1(n_510), .B2(n_498), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_654), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_672), .B(n_477), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_660), .B(n_679), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_635), .B(n_484), .Y(n_733) );
NOR2xp33_ASAP7_75t_SL g734 ( .A(n_679), .B(n_489), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_634), .A2(n_628), .B1(n_627), .B2(n_650), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_616), .A2(n_408), .B(n_405), .Y(n_736) );
NAND2xp33_ASAP7_75t_SL g737 ( .A(n_628), .B(n_509), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_690), .B(n_365), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_676), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_647), .B(n_512), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_690), .B(n_567), .Y(n_741) );
BUFx8_ASAP7_75t_L g742 ( .A(n_681), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_665), .A2(n_413), .B(n_412), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_655), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_683), .A2(n_421), .B(n_419), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_640), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_686), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_625), .B(n_516), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_643), .B(n_521), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_670), .A2(n_428), .B(n_427), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_678), .A2(n_463), .B(n_467), .C(n_433), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_645), .B(n_467), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_625), .B(n_429), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_653), .B(n_450), .C(n_441), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_630), .A2(n_461), .B1(n_469), .B2(n_459), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_646), .B(n_364), .Y(n_756) );
NOR2xp33_ASAP7_75t_R g757 ( .A(n_631), .B(n_368), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_674), .B(n_375), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_644), .B(n_348), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_657), .A2(n_505), .B(n_496), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_620), .B(n_378), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_621), .A2(n_508), .B1(n_514), .B2(n_506), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_682), .A2(n_517), .B(n_515), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_639), .B(n_348), .Y(n_764) );
NOR2xp67_ASAP7_75t_L g765 ( .A(n_637), .B(n_131), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_661), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_642), .A2(n_523), .B(n_519), .C(n_395), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_SL g768 ( .A1(n_693), .A2(n_537), .B(n_539), .C(n_528), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_694), .Y(n_769) );
O2A1O1Ixp33_ASAP7_75t_L g770 ( .A1(n_649), .A2(n_414), .B(n_422), .C(n_400), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_656), .A2(n_437), .B(n_422), .Y(n_771) );
INVx5_ASAP7_75t_L g772 ( .A(n_666), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_L g773 ( .A1(n_659), .A2(n_438), .B(n_456), .C(n_437), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g774 ( .A1(n_667), .A2(n_456), .B(n_458), .C(n_438), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g775 ( .A(n_671), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_623), .B(n_386), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_624), .B(n_371), .Y(n_777) );
AOI33xp33_ASAP7_75t_L g778 ( .A1(n_632), .A2(n_482), .A3(n_492), .B1(n_524), .B2(n_527), .B3(n_570), .Y(n_778) );
A2O1A1Ixp33_ASAP7_75t_L g779 ( .A1(n_688), .A2(n_524), .B(n_492), .C(n_407), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_692), .B(n_387), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_697), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_697), .B(n_348), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_684), .B(n_389), .Y(n_783) );
AO22x1_ASAP7_75t_L g784 ( .A1(n_675), .A2(n_390), .B1(n_397), .B2(n_396), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_696), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_698), .A2(n_596), .B(n_594), .Y(n_786) );
A2O1A1Ixp33_ASAP7_75t_L g787 ( .A1(n_689), .A2(n_407), .B(n_472), .C(n_528), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_695), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_687), .B(n_401), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_687), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_638), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_617), .B(n_417), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_617), .B(n_424), .Y(n_793) );
O2A1O1Ixp5_ASAP7_75t_SL g794 ( .A1(n_698), .A2(n_448), .B(n_562), .C(n_546), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_677), .A2(n_472), .B(n_537), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_617), .B(n_432), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_618), .A2(n_566), .B(n_570), .C(n_541), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_615), .Y(n_798) );
BUFx3_ASAP7_75t_L g799 ( .A(n_638), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_617), .B(n_439), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_615), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_638), .B(n_348), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g803 ( .A1(n_618), .A2(n_566), .B(n_570), .C(n_541), .Y(n_803) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_655), .Y(n_804) );
AO21x1_ASAP7_75t_L g805 ( .A1(n_614), .A2(n_566), .B(n_562), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_618), .A2(n_526), .B(n_501), .C(n_451), .Y(n_806) );
OR2x6_ASAP7_75t_SL g807 ( .A(n_654), .B(n_443), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_677), .A2(n_547), .B(n_598), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_617), .B(n_457), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_617), .B(n_473), .Y(n_810) );
BUFx12f_ASAP7_75t_L g811 ( .A(n_654), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_638), .B(n_501), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_677), .A2(n_547), .B(n_598), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_664), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_617), .B(n_476), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_617), .B(n_479), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_617), .B(n_481), .Y(n_817) );
O2A1O1Ixp5_ASAP7_75t_L g818 ( .A1(n_663), .A2(n_485), .B(n_499), .C(n_483), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_617), .B(n_503), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_617), .B(n_507), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_629), .A2(n_526), .B1(n_501), .B2(n_518), .Y(n_821) );
BUFx8_ASAP7_75t_L g822 ( .A(n_628), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_629), .A2(n_526), .B1(n_501), .B2(n_522), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_690), .A2(n_526), .B1(n_525), .B2(n_513), .C(n_546), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_629), .A2(n_547), .B1(n_562), .B2(n_546), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_617), .B(n_12), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_617), .B(n_13), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_629), .A2(n_562), .B1(n_564), .B2(n_546), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_798), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_791), .B(n_15), .Y(n_830) );
NAND3x1_ASAP7_75t_L g831 ( .A(n_729), .B(n_15), .C(n_16), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_808), .A2(n_600), .B(n_562), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_700), .Y(n_833) );
OA21x2_ASAP7_75t_L g834 ( .A1(n_805), .A2(n_562), .B(n_546), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_721), .B(n_16), .Y(n_835) );
NOR2xp67_ASAP7_75t_SL g836 ( .A(n_811), .B(n_17), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_799), .B(n_17), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_718), .B(n_18), .Y(n_838) );
INVx5_ASAP7_75t_L g839 ( .A(n_772), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_732), .B(n_18), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_748), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_748), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_812), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_753), .Y(n_844) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_722), .Y(n_845) );
OAI22x1_ASAP7_75t_L g846 ( .A1(n_729), .A2(n_727), .B1(n_731), .B2(n_734), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_701), .A2(n_564), .B(n_132), .Y(n_847) );
CKINVDCx14_ASAP7_75t_R g848 ( .A(n_807), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_706), .A2(n_564), .B(n_133), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_813), .A2(n_600), .B(n_564), .Y(n_850) );
AND2x6_ASAP7_75t_L g851 ( .A(n_801), .B(n_564), .Y(n_851) );
AND2x4_ASAP7_75t_L g852 ( .A(n_720), .B(n_20), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g853 ( .A1(n_708), .A2(n_600), .B(n_22), .C(n_20), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_753), .Y(n_854) );
OAI21xp5_ASAP7_75t_L g855 ( .A1(n_710), .A2(n_21), .B(n_22), .Y(n_855) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_724), .A2(n_21), .B(n_23), .Y(n_856) );
OAI22x1_ASAP7_75t_L g857 ( .A1(n_730), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_741), .B(n_24), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_801), .B(n_25), .Y(n_859) );
OA21x2_ASAP7_75t_L g860 ( .A1(n_711), .A2(n_600), .B(n_135), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_802), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_712), .A2(n_138), .B(n_136), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_738), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_863) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_822), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_705), .B(n_28), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_759), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_782), .Y(n_867) );
AND2x2_ASAP7_75t_SL g868 ( .A(n_769), .B(n_29), .Y(n_868) );
NAND2xp33_ASAP7_75t_L g869 ( .A(n_744), .B(n_600), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_719), .A2(n_29), .B(n_30), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_772), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_822), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_802), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_766), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_795), .A2(n_31), .B(n_32), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_781), .A2(n_34), .B1(n_31), .B2(n_32), .Y(n_876) );
NOR4xp25_ASAP7_75t_L g877 ( .A(n_751), .B(n_36), .C(n_34), .D(n_35), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_826), .A2(n_38), .B1(n_36), .B2(n_37), .Y(n_878) );
AOI21xp33_ASAP7_75t_L g879 ( .A1(n_793), .A2(n_39), .B(n_40), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_717), .B(n_704), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g881 ( .A(n_757), .B(n_600), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_699), .B(n_39), .Y(n_882) );
BUFx2_ASAP7_75t_L g883 ( .A(n_742), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_707), .B(n_41), .Y(n_884) );
AO31x2_ASAP7_75t_L g885 ( .A1(n_774), .A2(n_43), .A3(n_41), .B(n_42), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_726), .A2(n_714), .B(n_789), .Y(n_886) );
INVx1_ASAP7_75t_SL g887 ( .A(n_775), .Y(n_887) );
OAI21xp33_ASAP7_75t_L g888 ( .A1(n_749), .A2(n_752), .B(n_702), .Y(n_888) );
AO31x2_ASAP7_75t_L g889 ( .A1(n_779), .A2(n_45), .A3(n_42), .B(n_44), .Y(n_889) );
OAI22x1_ASAP7_75t_L g890 ( .A1(n_762), .A2(n_47), .B1(n_44), .B2(n_46), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_739), .Y(n_891) );
INVx4_ASAP7_75t_L g892 ( .A(n_772), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_788), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_827), .A2(n_48), .B1(n_46), .B2(n_47), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_733), .B(n_48), .Y(n_895) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_744), .Y(n_896) );
OAI21x1_ASAP7_75t_L g897 ( .A1(n_794), .A2(n_164), .B(n_156), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_728), .B(n_725), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_764), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_709), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_778), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_786), .A2(n_178), .B(n_170), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_770), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_755), .B(n_49), .Y(n_904) );
OA21x2_ASAP7_75t_L g905 ( .A1(n_771), .A2(n_182), .B(n_181), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_715), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_740), .B(n_50), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_787), .A2(n_185), .B(n_183), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_773), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_792), .B(n_53), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_796), .B(n_53), .Y(n_911) );
NOR2xp33_ASAP7_75t_R g912 ( .A(n_737), .B(n_54), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_715), .B(n_54), .Y(n_913) );
AND3x4_ASAP7_75t_L g914 ( .A(n_746), .B(n_55), .C(n_57), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_723), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_765), .A2(n_191), .B(n_189), .Y(n_916) );
OAI21xp5_ASAP7_75t_L g917 ( .A1(n_736), .A2(n_57), .B(n_60), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_777), .B(n_60), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_756), .A2(n_194), .B(n_193), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_742), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g921 ( .A1(n_818), .A2(n_61), .B(n_62), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g922 ( .A1(n_806), .A2(n_197), .B(n_196), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_767), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_735), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g925 ( .A1(n_780), .A2(n_201), .B(n_198), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_800), .B(n_63), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_743), .A2(n_206), .B(n_205), .Y(n_927) );
OR2x2_ASAP7_75t_L g928 ( .A(n_809), .B(n_65), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_703), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_716), .Y(n_930) );
AOI221xp5_ASAP7_75t_SL g931 ( .A1(n_760), .A2(n_65), .B1(n_66), .B2(n_67), .C(n_68), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_828), .A2(n_210), .B(n_209), .Y(n_932) );
A2O1A1Ixp33_ASAP7_75t_L g933 ( .A1(n_750), .A2(n_68), .B(n_69), .C(n_70), .Y(n_933) );
OAI21x1_ASAP7_75t_L g934 ( .A1(n_825), .A2(n_216), .B(n_215), .Y(n_934) );
AND2x4_ASAP7_75t_L g935 ( .A(n_713), .B(n_71), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_810), .B(n_71), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_824), .B(n_72), .Y(n_937) );
AOI221x1_ASAP7_75t_L g938 ( .A1(n_797), .A2(n_72), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_814), .Y(n_939) );
BUFx3_ASAP7_75t_L g940 ( .A(n_790), .Y(n_940) );
OAI21xp5_ASAP7_75t_L g941 ( .A1(n_803), .A2(n_77), .B(n_78), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_815), .B(n_77), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_763), .A2(n_79), .B(n_81), .C(n_82), .Y(n_943) );
CKINVDCx14_ASAP7_75t_R g944 ( .A(n_821), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_754), .A2(n_79), .B(n_82), .C(n_83), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g946 ( .A1(n_745), .A2(n_259), .B(n_328), .Y(n_946) );
NAND3x1_ASAP7_75t_L g947 ( .A(n_776), .B(n_83), .C(n_84), .Y(n_947) );
AOI211x1_ASAP7_75t_L g948 ( .A1(n_823), .A2(n_84), .B(n_85), .C(n_86), .Y(n_948) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_804), .Y(n_949) );
BUFx4_ASAP7_75t_SL g950 ( .A(n_768), .Y(n_950) );
AO21x2_ASAP7_75t_L g951 ( .A1(n_761), .A2(n_260), .B(n_327), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_816), .B(n_85), .Y(n_952) );
AND2x4_ASAP7_75t_L g953 ( .A(n_790), .B(n_86), .Y(n_953) );
AOI21xp5_ASAP7_75t_L g954 ( .A1(n_817), .A2(n_258), .B(n_323), .Y(n_954) );
INVx2_ASAP7_75t_SL g955 ( .A(n_783), .Y(n_955) );
OAI21x1_ASAP7_75t_SL g956 ( .A1(n_819), .A2(n_87), .B(n_88), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_758), .Y(n_957) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_820), .A2(n_88), .B(n_89), .C(n_90), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_784), .B(n_89), .Y(n_959) );
INVx5_ASAP7_75t_L g960 ( .A(n_785), .Y(n_960) );
AO21x2_ASAP7_75t_L g961 ( .A1(n_785), .A2(n_265), .B(n_322), .Y(n_961) );
AOI21xp5_ASAP7_75t_L g962 ( .A1(n_808), .A2(n_257), .B(n_321), .Y(n_962) );
AO31x2_ASAP7_75t_L g963 ( .A1(n_805), .A2(n_91), .A3(n_92), .B(n_94), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_791), .B(n_91), .Y(n_964) );
OAI21x1_ASAP7_75t_L g965 ( .A1(n_701), .A2(n_269), .B(n_320), .Y(n_965) );
BUFx3_ASAP7_75t_L g966 ( .A(n_822), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_805), .A2(n_254), .B(n_318), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_700), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_791), .B(n_96), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_791), .B(n_96), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_799), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_811), .Y(n_972) );
NAND2xp5_ASAP7_75t_SL g973 ( .A(n_799), .B(n_97), .Y(n_973) );
NOR3xp33_ASAP7_75t_L g974 ( .A(n_718), .B(n_98), .C(n_100), .Y(n_974) );
NOR2xp67_ASAP7_75t_L g975 ( .A(n_772), .B(n_220), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_718), .B(n_101), .C(n_102), .Y(n_976) );
INVx2_ASAP7_75t_SL g977 ( .A(n_822), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_700), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_747), .B(n_102), .Y(n_979) );
OAI21x1_ASAP7_75t_L g980 ( .A1(n_701), .A2(n_271), .B(n_316), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_700), .Y(n_981) );
OA21x2_ASAP7_75t_L g982 ( .A1(n_805), .A2(n_253), .B(n_312), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_791), .B(n_103), .Y(n_983) );
OAI21xp5_ASAP7_75t_L g984 ( .A1(n_706), .A2(n_274), .B(n_310), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_833), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g986 ( .A1(n_886), .A2(n_105), .B(n_106), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_968), .Y(n_987) );
AO21x2_ASAP7_75t_L g988 ( .A1(n_875), .A2(n_248), .B(n_306), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_978), .Y(n_989) );
AO31x2_ASAP7_75t_L g990 ( .A1(n_938), .A2(n_106), .A3(n_107), .B(n_108), .Y(n_990) );
BUFx2_ASAP7_75t_SL g991 ( .A(n_966), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_845), .B(n_108), .Y(n_992) );
OR2x6_ASAP7_75t_L g993 ( .A(n_977), .B(n_109), .Y(n_993) );
BUFx4f_ASAP7_75t_SL g994 ( .A(n_887), .Y(n_994) );
AO21x1_ASAP7_75t_L g995 ( .A1(n_856), .A2(n_109), .B(n_110), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_888), .B(n_111), .Y(n_996) );
OAI21x1_ASAP7_75t_L g997 ( .A1(n_965), .A2(n_247), .B(n_303), .Y(n_997) );
AND2x4_ASAP7_75t_L g998 ( .A(n_839), .B(n_111), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_888), .B(n_112), .Y(n_999) );
AO31x2_ASAP7_75t_L g1000 ( .A1(n_846), .A2(n_112), .A3(n_114), .B(n_115), .Y(n_1000) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_834), .A2(n_275), .B(n_302), .Y(n_1001) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_971), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_891), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_868), .B(n_115), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_848), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_880), .B(n_116), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_981), .Y(n_1007) );
INVx4_ASAP7_75t_L g1008 ( .A(n_839), .Y(n_1008) );
OAI21x1_ASAP7_75t_L g1009 ( .A1(n_980), .A2(n_241), .B(n_299), .Y(n_1009) );
BUFx2_ASAP7_75t_R g1010 ( .A(n_906), .Y(n_1010) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_883), .Y(n_1011) );
AND2x6_ASAP7_75t_L g1012 ( .A(n_859), .B(n_117), .Y(n_1012) );
OAI21x1_ASAP7_75t_L g1013 ( .A1(n_916), .A2(n_276), .B(n_298), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_893), .B(n_901), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_866), .A2(n_118), .B(n_119), .Y(n_1015) );
AO21x2_ASAP7_75t_L g1016 ( .A1(n_875), .A2(n_235), .B(n_294), .Y(n_1016) );
AO31x2_ASAP7_75t_L g1017 ( .A1(n_853), .A2(n_120), .A3(n_121), .B(n_123), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_852), .Y(n_1018) );
OAI21x1_ASAP7_75t_L g1019 ( .A1(n_897), .A2(n_280), .B(n_221), .Y(n_1019) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_910), .A2(n_284), .B(n_224), .Y(n_1020) );
AO21x1_ASAP7_75t_L g1021 ( .A1(n_856), .A2(n_121), .B(n_225), .Y(n_1021) );
OAI21x1_ASAP7_75t_L g1022 ( .A1(n_902), .A2(n_227), .B(n_228), .Y(n_1022) );
INVxp67_ASAP7_75t_SL g1023 ( .A(n_852), .Y(n_1023) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_849), .A2(n_232), .B(n_234), .Y(n_1024) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_839), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_874), .Y(n_1026) );
AO31x2_ASAP7_75t_L g1027 ( .A1(n_915), .A2(n_285), .A3(n_286), .B(n_288), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_887), .B(n_330), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_912), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_920), .Y(n_1030) );
NAND2x1p5_ASAP7_75t_L g1031 ( .A(n_960), .B(n_892), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_903), .A2(n_909), .B1(n_923), .B2(n_840), .Y(n_1032) );
OAI21xp5_ASAP7_75t_L g1033 ( .A1(n_838), .A2(n_957), .B(n_858), .Y(n_1033) );
AO21x2_ASAP7_75t_L g1034 ( .A1(n_921), .A2(n_922), .B(n_946), .Y(n_1034) );
AO21x2_ASAP7_75t_L g1035 ( .A1(n_921), .A2(n_941), .B(n_862), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_830), .B(n_964), .Y(n_1036) );
INVx5_ASAP7_75t_L g1037 ( .A(n_851), .Y(n_1037) );
AO21x1_ASAP7_75t_L g1038 ( .A1(n_941), .A2(n_924), .B(n_959), .Y(n_1038) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_871), .Y(n_1039) );
AOI21x1_ASAP7_75t_L g1040 ( .A1(n_967), .A2(n_982), .B(n_860), .Y(n_1040) );
BUFx2_ASAP7_75t_R g1041 ( .A(n_898), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_859), .Y(n_1042) );
AO21x2_ASAP7_75t_L g1043 ( .A1(n_984), .A2(n_956), .B(n_951), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_865), .A2(n_882), .B1(n_914), .B2(n_918), .Y(n_1044) );
OAI21x1_ASAP7_75t_SL g1045 ( .A1(n_855), .A2(n_870), .B(n_917), .Y(n_1045) );
INVx3_ASAP7_75t_L g1046 ( .A(n_892), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_863), .A2(n_904), .B1(n_974), .B2(n_879), .Y(n_1047) );
OA21x2_ASAP7_75t_L g1048 ( .A1(n_931), .A2(n_927), .B(n_934), .Y(n_1048) );
AO21x2_ASAP7_75t_L g1049 ( .A1(n_951), .A2(n_976), .B(n_917), .Y(n_1049) );
NOR2xp67_ASAP7_75t_SL g1050 ( .A(n_960), .B(n_896), .Y(n_1050) );
OAI21xp5_ASAP7_75t_L g1051 ( .A1(n_937), .A2(n_925), .B(n_907), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_936), .B(n_867), .Y(n_1052) );
OA21x2_ASAP7_75t_L g1053 ( .A1(n_931), .A2(n_976), .B(n_932), .Y(n_1053) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_935), .Y(n_1054) );
AND2x4_ASAP7_75t_L g1055 ( .A(n_844), .B(n_854), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_843), .B(n_841), .Y(n_1056) );
CKINVDCx11_ASAP7_75t_R g1057 ( .A(n_935), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_842), .B(n_884), .Y(n_1058) );
OA21x2_ASAP7_75t_L g1059 ( .A1(n_962), .A2(n_954), .B(n_919), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_953), .Y(n_1060) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_940), .Y(n_1061) );
INVx8_ASAP7_75t_L g1062 ( .A(n_851), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_955), .B(n_928), .Y(n_1063) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_913), .Y(n_1064) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_864), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_835), .Y(n_1066) );
OAI21x1_ASAP7_75t_L g1067 ( .A1(n_905), .A2(n_908), .B(n_975), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_837), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_900), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_929), .Y(n_1070) );
AOI221xp5_ASAP7_75t_L g1071 ( .A1(n_877), .A2(n_979), .B1(n_878), .B2(n_857), .C(n_890), .Y(n_1071) );
AO31x2_ASAP7_75t_L g1072 ( .A1(n_943), .A2(n_958), .A3(n_933), .B(n_945), .Y(n_1072) );
OAI21x1_ASAP7_75t_L g1073 ( .A1(n_881), .A2(n_899), .B(n_829), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_930), .Y(n_1074) );
BUFx8_ASAP7_75t_L g1075 ( .A(n_872), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_895), .A2(n_944), .B1(n_894), .B2(n_942), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_969), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_973), .Y(n_1078) );
NAND2x1p5_ASAP7_75t_L g1079 ( .A(n_949), .B(n_873), .Y(n_1079) );
AO31x2_ASAP7_75t_L g1080 ( .A1(n_876), .A2(n_926), .A3(n_952), .B(n_911), .Y(n_1080) );
NAND2x1_ASAP7_75t_L g1081 ( .A(n_851), .B(n_939), .Y(n_1081) );
AO31x2_ASAP7_75t_L g1082 ( .A1(n_963), .A2(n_983), .A3(n_970), .B(n_948), .Y(n_1082) );
OA21x2_ASAP7_75t_L g1083 ( .A1(n_963), .A2(n_861), .B(n_948), .Y(n_1083) );
NOR2x1_ASAP7_75t_SL g1084 ( .A(n_961), .B(n_831), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_963), .Y(n_1085) );
OAI21x1_ASAP7_75t_L g1086 ( .A1(n_947), .A2(n_869), .B(n_950), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1087 ( .A(n_961), .Y(n_1087) );
NAND2x1p5_ASAP7_75t_L g1088 ( .A(n_836), .B(n_877), .Y(n_1088) );
OA21x2_ASAP7_75t_L g1089 ( .A1(n_889), .A2(n_805), .B(n_847), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_889), .Y(n_1090) );
OAI21xp5_ASAP7_75t_L g1091 ( .A1(n_885), .A2(n_710), .B(n_706), .Y(n_1091) );
OAI21x1_ASAP7_75t_SL g1092 ( .A1(n_885), .A2(n_946), .B(n_855), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_885), .Y(n_1093) );
NAND2x1p5_ASAP7_75t_L g1094 ( .A(n_839), .B(n_960), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_924), .A2(n_729), .B1(n_852), .B2(n_856), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_839), .B(n_799), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_839), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g1098 ( .A(n_839), .Y(n_1098) );
NAND2x1p5_ASAP7_75t_L g1099 ( .A(n_839), .B(n_960), .Y(n_1099) );
AND3x2_ASAP7_75t_L g1100 ( .A(n_883), .B(n_731), .C(n_734), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_839), .B(n_799), .Y(n_1101) );
AOI21x1_ASAP7_75t_L g1102 ( .A1(n_834), .A2(n_805), .B(n_701), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_891), .Y(n_1103) );
AOI21xp33_ASAP7_75t_SL g1104 ( .A1(n_914), .A2(n_868), .B(n_672), .Y(n_1104) );
AO21x2_ASAP7_75t_L g1105 ( .A1(n_875), .A2(n_805), .B(n_849), .Y(n_1105) );
NOR2x1_ASAP7_75t_SL g1106 ( .A(n_839), .B(n_960), .Y(n_1106) );
BUFx3_ASAP7_75t_L g1107 ( .A(n_966), .Y(n_1107) );
AOI21x1_ASAP7_75t_L g1108 ( .A1(n_834), .A2(n_805), .B(n_701), .Y(n_1108) );
OAI21xp5_ASAP7_75t_L g1109 ( .A1(n_886), .A2(n_710), .B(n_706), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_891), .Y(n_1110) );
CKINVDCx8_ASAP7_75t_R g1111 ( .A(n_972), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_839), .B(n_799), .Y(n_1112) );
AOI21xp5_ASAP7_75t_L g1113 ( .A1(n_832), .A2(n_711), .B(n_850), .Y(n_1113) );
NAND2x1p5_ASAP7_75t_L g1114 ( .A(n_839), .B(n_960), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_891), .Y(n_1115) );
CKINVDCx9p33_ASAP7_75t_R g1116 ( .A(n_883), .Y(n_1116) );
BUFx6f_ASAP7_75t_L g1117 ( .A(n_839), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_833), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_891), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_891), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_833), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_891), .Y(n_1122) );
OAI21x1_ASAP7_75t_SL g1123 ( .A1(n_946), .A2(n_855), .B(n_870), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_833), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_985), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1126 ( .A(n_1097), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_987), .Y(n_1127) );
INVx3_ASAP7_75t_L g1128 ( .A(n_1062), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_1037), .B(n_1023), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1003), .B(n_1103), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1110), .B(n_1115), .Y(n_1131) );
OAI21x1_ASAP7_75t_L g1132 ( .A1(n_1067), .A2(n_1108), .B(n_1102), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1096), .Y(n_1133) );
INVx3_ASAP7_75t_L g1134 ( .A(n_1062), .Y(n_1134) );
INVx3_ASAP7_75t_L g1135 ( .A(n_1062), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_989), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_1037), .B(n_1023), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1007), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1002), .B(n_1074), .Y(n_1139) );
NAND2x1_ASAP7_75t_L g1140 ( .A(n_1012), .B(n_1050), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1119), .B(n_1120), .Y(n_1141) );
AO21x2_ASAP7_75t_L g1142 ( .A1(n_1092), .A2(n_1123), .B(n_1045), .Y(n_1142) );
INVx3_ASAP7_75t_L g1143 ( .A(n_1037), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1122), .B(n_1026), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1032), .B(n_1033), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g1146 ( .A(n_1075), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_1096), .Y(n_1147) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_1094), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1085), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1101), .Y(n_1150) );
BUFx3_ASAP7_75t_L g1151 ( .A(n_1094), .Y(n_1151) );
OA21x2_ASAP7_75t_L g1152 ( .A1(n_1040), .A2(n_1093), .B(n_1090), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1118), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1044), .B(n_1121), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1089), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1032), .B(n_1033), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g1157 ( .A(n_1104), .B(n_1095), .Y(n_1157) );
OAI211xp5_ASAP7_75t_SL g1158 ( .A1(n_1057), .A2(n_1044), .B(n_1071), .C(n_1076), .Y(n_1158) );
OAI21xp5_ASAP7_75t_L g1159 ( .A1(n_1047), .A2(n_1051), .B(n_986), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_1099), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1069), .B(n_1124), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1014), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_1099), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1112), .B(n_1064), .Y(n_1164) );
INVx1_ASAP7_75t_SL g1165 ( .A(n_1116), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1056), .Y(n_1166) );
INVxp67_ASAP7_75t_L g1167 ( .A(n_1065), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1056), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_998), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_1114), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1042), .B(n_1015), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_998), .Y(n_1172) );
AOI21x1_ASAP7_75t_L g1173 ( .A1(n_1081), .A2(n_1053), .B(n_1048), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_1112), .Y(n_1174) );
INVx3_ASAP7_75t_L g1175 ( .A(n_1114), .Y(n_1175) );
AO21x2_ASAP7_75t_L g1176 ( .A1(n_1049), .A2(n_986), .B(n_1034), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1106), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_992), .B(n_1083), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1054), .B(n_1104), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1052), .Y(n_1180) );
NAND2xp5_ASAP7_75t_SL g1181 ( .A(n_1021), .B(n_1038), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1083), .B(n_1082), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_1098), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1055), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1185 ( .A(n_1075), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1055), .Y(n_1186) );
OR2x6_ASAP7_75t_L g1187 ( .A(n_1008), .B(n_1031), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1082), .B(n_1006), .Y(n_1188) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_1098), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1063), .B(n_1041), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1029), .B(n_1039), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1018), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1025), .Y(n_1193) );
AND2x4_ASAP7_75t_L g1194 ( .A(n_1060), .B(n_1025), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1006), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_996), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1082), .B(n_1066), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_996), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1199 ( .A(n_1098), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_999), .Y(n_1200) );
AO21x2_ASAP7_75t_L g1201 ( .A1(n_1049), .A2(n_1034), .B(n_1035), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1117), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_999), .Y(n_1203) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1046), .B(n_1008), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1117), .Y(n_1205) );
AO21x2_ASAP7_75t_L g1206 ( .A1(n_1035), .A2(n_1105), .B(n_1001), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1117), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_993), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1027), .Y(n_1209) );
CKINVDCx9p33_ASAP7_75t_R g1210 ( .A(n_1116), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1088), .B(n_1068), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_993), .Y(n_1212) );
HB1xp67_ASAP7_75t_L g1213 ( .A(n_1031), .Y(n_1213) );
OA21x2_ASAP7_75t_L g1214 ( .A1(n_1113), .A2(n_1087), .B(n_1001), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1058), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1004), .B(n_1036), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1058), .Y(n_1217) );
OR2x6_ASAP7_75t_L g1218 ( .A(n_1086), .B(n_1088), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1077), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1070), .Y(n_1220) );
INVx1_ASAP7_75t_SL g1221 ( .A(n_991), .Y(n_1221) );
INVx3_ASAP7_75t_L g1222 ( .A(n_1046), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_995), .Y(n_1223) );
AO21x1_ASAP7_75t_SL g1224 ( .A1(n_1100), .A2(n_1057), .B(n_1028), .Y(n_1224) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1061), .Y(n_1225) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_1011), .Y(n_1226) );
INVx1_ASAP7_75t_SL g1227 ( .A(n_1011), .Y(n_1227) );
OAI21xp5_ASAP7_75t_L g1228 ( .A1(n_1051), .A2(n_1091), .B(n_1109), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1017), .B(n_1080), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1017), .B(n_1080), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1197), .B(n_1000), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1180), .B(n_1100), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1145), .B(n_1000), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1149), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1178), .B(n_1017), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1145), .B(n_990), .Y(n_1236) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1155), .Y(n_1237) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1218), .B(n_1084), .Y(n_1238) );
AOI22xp33_ASAP7_75t_SL g1239 ( .A1(n_1157), .A2(n_994), .B1(n_1078), .B2(n_1016), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1125), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1156), .B(n_990), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1127), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1136), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1215), .B(n_1080), .Y(n_1244) );
NOR2x1_ASAP7_75t_L g1245 ( .A(n_1177), .B(n_1107), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1178), .B(n_990), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1138), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1156), .B(n_1072), .Y(n_1248) );
INVxp67_ASAP7_75t_SL g1249 ( .A(n_1126), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1217), .B(n_1030), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1154), .B(n_1072), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1229), .B(n_1105), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1152), .Y(n_1253) );
OAI31xp33_ASAP7_75t_L g1254 ( .A1(n_1158), .A2(n_1041), .A3(n_1020), .B(n_1079), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1229), .B(n_1043), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1230), .B(n_1091), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1182), .B(n_1072), .Y(n_1257) );
NAND2xp33_ASAP7_75t_R g1258 ( .A(n_1185), .B(n_1005), .Y(n_1258) );
OR2x2_ASAP7_75t_SL g1259 ( .A(n_1210), .B(n_1024), .Y(n_1259) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_1218), .B(n_1073), .Y(n_1260) );
BUFx3_ASAP7_75t_L g1261 ( .A(n_1151), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1188), .B(n_1161), .Y(n_1262) );
BUFx2_ASAP7_75t_L g1263 ( .A(n_1129), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1218), .B(n_1087), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1153), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_1218), .B(n_988), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1267 ( .A(n_1139), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1188), .B(n_1109), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1219), .Y(n_1269) );
INVxp67_ASAP7_75t_L g1270 ( .A(n_1226), .Y(n_1270) );
BUFx3_ASAP7_75t_L g1271 ( .A(n_1151), .Y(n_1271) );
AND2x4_ASAP7_75t_SL g1272 ( .A(n_1187), .B(n_1213), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1228), .B(n_1059), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1130), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1131), .Y(n_1275) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_1140), .Y(n_1276) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_1167), .Y(n_1277) );
INVxp67_ASAP7_75t_L g1278 ( .A(n_1225), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1202), .Y(n_1279) );
INVxp67_ASAP7_75t_SL g1280 ( .A(n_1129), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1141), .B(n_1013), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1148), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1144), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1159), .B(n_1022), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1211), .B(n_1009), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1216), .B(n_997), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1166), .Y(n_1287) );
INVxp67_ASAP7_75t_SL g1288 ( .A(n_1137), .Y(n_1288) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_1133), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_1137), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1196), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1168), .B(n_1111), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1211), .B(n_1019), .Y(n_1293) );
CKINVDCx20_ASAP7_75t_R g1294 ( .A(n_1146), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1171), .B(n_1010), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1192), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1162), .B(n_1195), .Y(n_1297) );
INVx3_ASAP7_75t_L g1298 ( .A(n_1143), .Y(n_1298) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_1238), .B(n_1142), .Y(n_1299) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1253), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_1238), .B(n_1142), .Y(n_1301) );
AND2x4_ASAP7_75t_SL g1302 ( .A(n_1279), .B(n_1187), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1262), .B(n_1176), .Y(n_1303) );
CKINVDCx20_ASAP7_75t_R g1304 ( .A(n_1294), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1269), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1267), .B(n_1164), .Y(n_1306) );
INVx1_ASAP7_75t_SL g1307 ( .A(n_1294), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1257), .B(n_1176), .Y(n_1308) );
HB1xp67_ASAP7_75t_L g1309 ( .A(n_1249), .Y(n_1309) );
INVx2_ASAP7_75t_SL g1310 ( .A(n_1272), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1240), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1242), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1257), .B(n_1176), .Y(n_1313) );
AND2x4_ASAP7_75t_L g1314 ( .A(n_1238), .B(n_1173), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1274), .B(n_1208), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1268), .B(n_1201), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1268), .B(n_1201), .Y(n_1317) );
AND2x4_ASAP7_75t_L g1318 ( .A(n_1260), .B(n_1132), .Y(n_1318) );
INVx3_ASAP7_75t_L g1319 ( .A(n_1260), .Y(n_1319) );
NAND2xp5_ASAP7_75t_SL g1320 ( .A(n_1239), .B(n_1165), .Y(n_1320) );
BUFx2_ASAP7_75t_SL g1321 ( .A(n_1261), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1256), .B(n_1201), .Y(n_1322) );
INVx1_ASAP7_75t_SL g1323 ( .A(n_1272), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1243), .Y(n_1324) );
INVx4_ASAP7_75t_L g1325 ( .A(n_1261), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1256), .B(n_1198), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1235), .B(n_1200), .Y(n_1327) );
BUFx3_ASAP7_75t_L g1328 ( .A(n_1271), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1275), .B(n_1212), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1235), .B(n_1203), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1247), .Y(n_1331) );
INVxp67_ASAP7_75t_SL g1332 ( .A(n_1289), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1292), .B(n_1227), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1246), .B(n_1206), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1248), .B(n_1223), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1248), .B(n_1179), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1246), .B(n_1206), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1231), .B(n_1206), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1265), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1231), .B(n_1209), .Y(n_1340) );
AND2x4_ASAP7_75t_SL g1341 ( .A(n_1298), .B(n_1187), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1244), .B(n_1181), .Y(n_1342) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1237), .Y(n_1343) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1233), .B(n_1181), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1296), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1297), .Y(n_1346) );
AND2x4_ASAP7_75t_L g1347 ( .A(n_1266), .B(n_1132), .Y(n_1347) );
INVx1_ASAP7_75t_SL g1348 ( .A(n_1271), .Y(n_1348) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_1234), .Y(n_1349) );
BUFx2_ASAP7_75t_L g1350 ( .A(n_1245), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1252), .B(n_1214), .Y(n_1351) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_1270), .B(n_1221), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1297), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1283), .B(n_1174), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1287), .Y(n_1355) );
HB1xp67_ASAP7_75t_L g1356 ( .A(n_1278), .Y(n_1356) );
INVx3_ASAP7_75t_R g1357 ( .A(n_1258), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1255), .B(n_1214), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1277), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1305), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1311), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1309), .B(n_1263), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1316), .B(n_1251), .Y(n_1363) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1300), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1312), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1324), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1326), .B(n_1263), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1331), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1326), .B(n_1290), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1339), .Y(n_1370) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_1320), .A2(n_1295), .B1(n_1190), .B2(n_1232), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1336), .B(n_1290), .Y(n_1372) );
OR2x6_ASAP7_75t_L g1373 ( .A(n_1321), .B(n_1266), .Y(n_1373) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1336), .B(n_1236), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1359), .B(n_1295), .Y(n_1375) );
AND2x4_ASAP7_75t_L g1376 ( .A(n_1299), .B(n_1264), .Y(n_1376) );
HB1xp67_ASAP7_75t_L g1377 ( .A(n_1349), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1345), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1316), .B(n_1291), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1355), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1332), .B(n_1236), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1317), .B(n_1291), .Y(n_1382) );
NAND2x1p5_ASAP7_75t_L g1383 ( .A(n_1325), .B(n_1163), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1384 ( .A(n_1346), .B(n_1353), .Y(n_1384) );
NAND2xp5_ASAP7_75t_SL g1385 ( .A(n_1325), .B(n_1276), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1327), .B(n_1280), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1327), .B(n_1288), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1343), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1317), .B(n_1241), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1330), .B(n_1285), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1356), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1315), .Y(n_1392) );
INVx1_ASAP7_75t_SL g1393 ( .A(n_1348), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1322), .B(n_1273), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1330), .B(n_1285), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1303), .B(n_1293), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1329), .Y(n_1397) );
AND2x4_ASAP7_75t_L g1398 ( .A(n_1299), .B(n_1264), .Y(n_1398) );
AND2x4_ASAP7_75t_L g1399 ( .A(n_1299), .B(n_1264), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1322), .B(n_1273), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1303), .B(n_1293), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1306), .B(n_1234), .Y(n_1402) );
INVx1_ASAP7_75t_SL g1403 ( .A(n_1328), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1350), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1354), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1340), .B(n_1255), .Y(n_1406) );
INVx5_ASAP7_75t_SL g1407 ( .A(n_1357), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1396), .B(n_1358), .Y(n_1408) );
NAND2xp5_ASAP7_75t_SL g1409 ( .A(n_1385), .B(n_1325), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1360), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1401), .B(n_1358), .Y(n_1411) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_1371), .A2(n_1310), .B1(n_1323), .B2(n_1320), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1392), .B(n_1308), .Y(n_1413) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_1376), .B(n_1301), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1361), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1394), .B(n_1344), .Y(n_1416) );
AND2x4_ASAP7_75t_SL g1417 ( .A(n_1373), .B(n_1310), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1397), .B(n_1313), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1405), .B(n_1313), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1365), .Y(n_1420) );
A2O1A1Ixp33_ASAP7_75t_L g1421 ( .A1(n_1385), .A2(n_1302), .B(n_1341), .C(n_1190), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1379), .B(n_1338), .Y(n_1422) );
INVx1_ASAP7_75t_SL g1423 ( .A(n_1393), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1366), .Y(n_1424) );
INVx2_ASAP7_75t_SL g1425 ( .A(n_1377), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1406), .B(n_1351), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1368), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1390), .B(n_1351), .Y(n_1428) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1394), .B(n_1344), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1379), .B(n_1338), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1370), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1378), .Y(n_1432) );
INVx2_ASAP7_75t_SL g1433 ( .A(n_1377), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1380), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1384), .Y(n_1435) );
INVx2_ASAP7_75t_SL g1436 ( .A(n_1403), .Y(n_1436) );
BUFx2_ASAP7_75t_L g1437 ( .A(n_1403), .Y(n_1437) );
INVx3_ASAP7_75t_L g1438 ( .A(n_1373), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1395), .B(n_1334), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1400), .B(n_1334), .Y(n_1440) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1364), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1400), .B(n_1337), .Y(n_1442) );
HB1xp67_ASAP7_75t_L g1443 ( .A(n_1388), .Y(n_1443) );
OAI21xp5_ASAP7_75t_L g1444 ( .A1(n_1421), .A2(n_1383), .B(n_1304), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_1412), .A2(n_1301), .B1(n_1404), .B2(n_1375), .Y(n_1445) );
OAI32xp33_ASAP7_75t_L g1446 ( .A1(n_1438), .A2(n_1383), .A3(n_1307), .B1(n_1362), .B2(n_1304), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1440), .B(n_1363), .Y(n_1447) );
NOR2xp33_ASAP7_75t_L g1448 ( .A(n_1423), .B(n_1391), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1410), .Y(n_1449) );
AOI211xp5_ASAP7_75t_L g1450 ( .A1(n_1409), .A2(n_1254), .B(n_1381), .C(n_1352), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1415), .Y(n_1451) );
OAI21xp33_ASAP7_75t_SL g1452 ( .A1(n_1409), .A2(n_1373), .B(n_1369), .Y(n_1452) );
OAI21xp33_ASAP7_75t_L g1453 ( .A1(n_1416), .A2(n_1382), .B(n_1389), .Y(n_1453) );
OAI21xp33_ASAP7_75t_L g1454 ( .A1(n_1416), .A2(n_1382), .B(n_1389), .Y(n_1454) );
INVx1_ASAP7_75t_SL g1455 ( .A(n_1437), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1420), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1424), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1427), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1428), .B(n_1376), .Y(n_1459) );
NOR2xp67_ASAP7_75t_L g1460 ( .A(n_1438), .B(n_1388), .Y(n_1460) );
AOI32xp33_ASAP7_75t_L g1461 ( .A1(n_1417), .A2(n_1302), .A3(n_1367), .B1(n_1387), .B2(n_1386), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1428), .B(n_1398), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1429), .B(n_1374), .Y(n_1463) );
INVxp67_ASAP7_75t_L g1464 ( .A(n_1425), .Y(n_1464) );
INVx3_ASAP7_75t_L g1465 ( .A(n_1417), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1453), .B(n_1440), .Y(n_1466) );
AOI21xp5_ASAP7_75t_L g1467 ( .A1(n_1444), .A2(n_1433), .B(n_1425), .Y(n_1467) );
INVxp67_ASAP7_75t_L g1468 ( .A(n_1455), .Y(n_1468) );
INVx1_ASAP7_75t_SL g1469 ( .A(n_1465), .Y(n_1469) );
OAI21xp5_ASAP7_75t_SL g1470 ( .A1(n_1444), .A2(n_1341), .B(n_1433), .Y(n_1470) );
OAI32xp33_ASAP7_75t_L g1471 ( .A1(n_1452), .A2(n_1429), .A3(n_1436), .B1(n_1443), .B2(n_1328), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1472 ( .A(n_1463), .B(n_1422), .Y(n_1472) );
AOI32xp33_ASAP7_75t_L g1473 ( .A1(n_1465), .A2(n_1414), .A3(n_1411), .B1(n_1408), .B2(n_1435), .Y(n_1473) );
O2A1O1Ixp33_ASAP7_75t_L g1474 ( .A1(n_1446), .A2(n_1333), .B(n_1250), .C(n_1220), .Y(n_1474) );
AOI221xp5_ASAP7_75t_L g1475 ( .A1(n_1454), .A2(n_1419), .B1(n_1432), .B2(n_1434), .C(n_1431), .Y(n_1475) );
O2A1O1Ixp33_ASAP7_75t_L g1476 ( .A1(n_1464), .A2(n_1282), .B(n_1418), .C(n_1413), .Y(n_1476) );
O2A1O1Ixp33_ASAP7_75t_L g1477 ( .A1(n_1464), .A2(n_1172), .B(n_1169), .C(n_1191), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1449), .Y(n_1478) );
AOI221xp5_ASAP7_75t_SL g1479 ( .A1(n_1445), .A2(n_1442), .B1(n_1430), .B2(n_1439), .C(n_1411), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_1447), .B(n_1442), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1451), .Y(n_1481) );
OAI21xp5_ASAP7_75t_L g1482 ( .A1(n_1460), .A2(n_1170), .B(n_1160), .Y(n_1482) );
AOI22xp5_ASAP7_75t_L g1483 ( .A1(n_1469), .A2(n_1450), .B1(n_1448), .B2(n_1407), .Y(n_1483) );
OAI31xp33_ASAP7_75t_L g1484 ( .A1(n_1470), .A2(n_1459), .A3(n_1462), .B(n_1456), .Y(n_1484) );
AOI211xp5_ASAP7_75t_L g1485 ( .A1(n_1471), .A2(n_1414), .B(n_1458), .C(n_1457), .Y(n_1485) );
AOI221x1_ASAP7_75t_L g1486 ( .A1(n_1467), .A2(n_1447), .B1(n_1193), .B2(n_1205), .C(n_1207), .Y(n_1486) );
AOI22xp33_ASAP7_75t_SL g1487 ( .A1(n_1482), .A2(n_1319), .B1(n_1398), .B2(n_1399), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1479), .B(n_1439), .Y(n_1488) );
AOI22xp33_ASAP7_75t_SL g1489 ( .A1(n_1482), .A2(n_1319), .B1(n_1399), .B2(n_1301), .Y(n_1489) );
NOR2xp33_ASAP7_75t_L g1490 ( .A(n_1468), .B(n_1408), .Y(n_1490) );
NOR3xp33_ASAP7_75t_SL g1491 ( .A(n_1474), .B(n_1210), .C(n_1224), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1478), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1493 ( .A(n_1475), .B(n_1426), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1494 ( .A(n_1480), .B(n_1402), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1483), .B(n_1466), .Y(n_1495) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_1492), .Y(n_1496) );
NAND3xp33_ASAP7_75t_L g1497 ( .A(n_1485), .B(n_1473), .C(n_1476), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1488), .B(n_1481), .Y(n_1498) );
NAND4xp25_ASAP7_75t_SL g1499 ( .A(n_1484), .B(n_1461), .C(n_1477), .D(n_1472), .Y(n_1499) );
NAND2xp5_ASAP7_75t_SL g1500 ( .A(n_1491), .B(n_1314), .Y(n_1500) );
OAI21xp33_ASAP7_75t_L g1501 ( .A1(n_1493), .A2(n_1335), .B(n_1372), .Y(n_1501) );
NOR2x1_ASAP7_75t_L g1502 ( .A(n_1490), .B(n_1187), .Y(n_1502) );
OAI211xp5_ASAP7_75t_L g1503 ( .A1(n_1487), .A2(n_1150), .B(n_1147), .C(n_1286), .Y(n_1503) );
AOI211xp5_ASAP7_75t_L g1504 ( .A1(n_1499), .A2(n_1497), .B(n_1500), .C(n_1503), .Y(n_1504) );
AND2x2_ASAP7_75t_SL g1505 ( .A(n_1495), .B(n_1486), .Y(n_1505) );
NOR3x1_ASAP7_75t_L g1506 ( .A(n_1498), .B(n_1489), .C(n_1170), .Y(n_1506) );
NOR2xp33_ASAP7_75t_L g1507 ( .A(n_1501), .B(n_1494), .Y(n_1507) );
NOR2x1_ASAP7_75t_L g1508 ( .A(n_1502), .B(n_1175), .Y(n_1508) );
NOR2xp33_ASAP7_75t_SL g1509 ( .A(n_1496), .B(n_1160), .Y(n_1509) );
NOR2x1p5_ASAP7_75t_L g1510 ( .A(n_1504), .B(n_1175), .Y(n_1510) );
NAND4xp75_ASAP7_75t_L g1511 ( .A(n_1506), .B(n_1183), .C(n_1199), .D(n_1189), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1507), .B(n_1441), .Y(n_1512) );
NAND5xp2_ASAP7_75t_L g1513 ( .A(n_1509), .B(n_1284), .C(n_1184), .D(n_1186), .E(n_1281), .Y(n_1513) );
AOI22xp5_ASAP7_75t_L g1514 ( .A1(n_1505), .A2(n_1318), .B1(n_1266), .B2(n_1347), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1510), .B(n_1508), .Y(n_1515) );
INVx2_ASAP7_75t_L g1516 ( .A(n_1512), .Y(n_1516) );
INVx2_ASAP7_75t_L g1517 ( .A(n_1511), .Y(n_1517) );
INVx2_ASAP7_75t_L g1518 ( .A(n_1514), .Y(n_1518) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1513), .Y(n_1519) );
INVx4_ASAP7_75t_L g1520 ( .A(n_1517), .Y(n_1520) );
AOI31xp33_ASAP7_75t_L g1521 ( .A1(n_1519), .A2(n_1516), .A3(n_1518), .B(n_1515), .Y(n_1521) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1516), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_1521), .A2(n_1259), .B1(n_1342), .B2(n_1335), .Y(n_1523) );
AO22x2_ASAP7_75t_L g1524 ( .A1(n_1520), .A2(n_1175), .B1(n_1204), .B2(n_1199), .Y(n_1524) );
OAI21xp5_ASAP7_75t_L g1525 ( .A1(n_1522), .A2(n_1204), .B(n_1183), .Y(n_1525) );
O2A1O1Ixp33_ASAP7_75t_L g1526 ( .A1(n_1525), .A2(n_1520), .B(n_1134), .C(n_1135), .Y(n_1526) );
NOR3xp33_ASAP7_75t_L g1527 ( .A(n_1523), .B(n_1128), .C(n_1134), .Y(n_1527) );
OAI21xp5_ASAP7_75t_L g1528 ( .A1(n_1526), .A2(n_1524), .B(n_1204), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1527), .B(n_1222), .Y(n_1529) );
OR2x6_ASAP7_75t_L g1530 ( .A(n_1528), .B(n_1128), .Y(n_1530) );
AO21x2_ASAP7_75t_L g1531 ( .A1(n_1529), .A2(n_1194), .B(n_1441), .Y(n_1531) );
AOI21xp5_ASAP7_75t_L g1532 ( .A1(n_1530), .A2(n_1135), .B(n_1143), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_1532), .A2(n_1531), .B1(n_1318), .B2(n_1314), .Y(n_1533) );
endmodule