module fake_jpeg_9324_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_31;
wire n_17;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_4),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_1),
.B1(n_4),
.B2(n_7),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_12),
.B1(n_10),
.B2(n_14),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_22),
.B(n_27),
.C(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_23),
.Y(n_32)
);

FAx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_23),
.CI(n_9),
.CON(n_35),
.SN(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_22),
.C(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_34),
.B(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_49),
.B(n_50),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.C(n_35),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_44),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_31),
.B(n_35),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_41),
.C(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_27),
.Y(n_61)
);


endmodule