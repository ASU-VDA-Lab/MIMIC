module fake_ariane_3360_n_1764 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1764);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1764;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_18),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_44),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_41),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_59),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_57),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_43),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_16),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_34),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_83),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_25),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_77),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_39),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_128),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_69),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_72),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_50),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_12),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_23),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_5),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_130),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_38),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_87),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_112),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_86),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_38),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_66),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_20),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_45),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_41),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_28),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_46),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_17),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_92),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_99),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_45),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_144),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_96),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_73),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_88),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_48),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_113),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_28),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_12),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_81),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_51),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_71),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_135),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_37),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_121),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_50),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_60),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_103),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_124),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_9),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_48),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_139),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_7),
.Y(n_268)
);

BUFx8_ASAP7_75t_SL g269 ( 
.A(n_148),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_82),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_9),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_20),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_5),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_44),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_109),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_19),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_125),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_39),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_126),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_11),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_0),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_94),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_17),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_141),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_118),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_115),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_26),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_140),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_102),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_111),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_49),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_91),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_52),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_133),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_79),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_75),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_117),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_137),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_127),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_129),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_123),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_156),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_156),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_228),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_166),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_173),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_173),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_181),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_219),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_202),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_192),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_241),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_242),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_237),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_163),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_165),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_255),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_219),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_198),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_198),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_213),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_162),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_219),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_200),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_157),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_205),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_269),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_205),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_253),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_263),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_209),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_253),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_303),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_221),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_227),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_230),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_158),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_230),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_231),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_241),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_159),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_231),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_168),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_241),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_211),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_176),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_178),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_180),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_246),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_246),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_183),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_193),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_241),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_248),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_248),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_196),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_241),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_165),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_249),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_197),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_204),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_170),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_265),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_170),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_355),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_265),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_314),
.B(n_172),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_333),
.B(n_160),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_384),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_336),
.B(n_160),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_382),
.B1(n_344),
.B2(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

BUFx8_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_361),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_334),
.B(n_172),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_318),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_326),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_388),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_339),
.B(n_164),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_380),
.A2(n_251),
.B1(n_268),
.B2(n_273),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_343),
.B(n_195),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_282),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_322),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_336),
.B(n_174),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_358),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_359),
.B(n_304),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_317),
.B(n_195),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_366),
.B(n_203),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_374),
.A2(n_223),
.B(n_203),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_375),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

INVx6_ASAP7_75t_L g459 ( 
.A(n_349),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_355),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_328),
.A2(n_233),
.B(n_223),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_342),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_402),
.A2(n_382),
.B1(n_344),
.B2(n_282),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_405),
.A2(n_327),
.B1(n_330),
.B2(n_335),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_433),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_413),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_433),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_399),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_462),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_462),
.B(n_327),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_330),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_396),
.B(n_324),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_462),
.B(n_335),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_414),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

NOR2x1p5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_347),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_462),
.B(n_370),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_440),
.B(n_315),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_371),
.C(n_370),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_462),
.B(n_371),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_452),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_399),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

NOR2x1p5_ASAP7_75t_L g511 ( 
.A(n_463),
.B(n_347),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_460),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_396),
.B(n_372),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_457),
.B(n_372),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_414),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_R g525 ( 
.A(n_460),
.B(n_340),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_409),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_390),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_457),
.B(n_373),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_440),
.B(n_373),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_459),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_398),
.B(n_376),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_439),
.B(n_346),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_398),
.B(n_404),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_458),
.B(n_377),
.C(n_376),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_406),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_390),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_442),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_390),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_439),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_390),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_407),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_426),
.Y(n_547)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_463),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_402),
.A2(n_458),
.B1(n_457),
.B2(n_422),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_457),
.B(n_377),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_402),
.A2(n_283),
.B1(n_276),
.B2(n_164),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_407),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_394),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_408),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_404),
.B(n_386),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_463),
.B(n_338),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_408),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_430),
.B(n_253),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_422),
.B(n_208),
.C(n_207),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_397),
.A2(n_289),
.B1(n_258),
.B2(n_256),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_427),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_421),
.A2(n_235),
.B(n_233),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

OAI21xp33_ASAP7_75t_SL g566 ( 
.A1(n_420),
.A2(n_283),
.B(n_268),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_459),
.B(n_167),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_427),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_443),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_443),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_463),
.B(n_217),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_461),
.A2(n_276),
.B1(n_167),
.B2(n_187),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_443),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_443),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_453),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_409),
.B(n_369),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_461),
.A2(n_187),
.B1(n_186),
.B2(n_296),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_453),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_393),
.B(n_235),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_415),
.B(n_350),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_415),
.B(n_218),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_453),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_394),
.B(n_243),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_461),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_433),
.B(n_251),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_453),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_416),
.B(n_243),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_456),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_456),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_393),
.B(n_254),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_417),
.B(n_222),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_461),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_393),
.B(n_254),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_393),
.B(n_186),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_393),
.B(n_259),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_456),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_456),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_400),
.B(n_259),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_487),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_559),
.B(n_400),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_549),
.B(n_417),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_L g616 ( 
.A(n_474),
.B(n_436),
.C(n_419),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_419),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_606),
.A2(n_434),
.B1(n_412),
.B2(n_401),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_522),
.B(n_412),
.Y(n_619)
);

O2A1O1Ixp5_ASAP7_75t_L g620 ( 
.A1(n_576),
.A2(n_403),
.B(n_423),
.C(n_411),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_533),
.B(n_412),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_559),
.B(n_400),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_400),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_525),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_466),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_468),
.B(n_400),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_556),
.B(n_412),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_531),
.B(n_412),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_464),
.A2(n_420),
.B1(n_459),
.B2(n_449),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_468),
.B(n_397),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_499),
.A2(n_459),
.B1(n_455),
.B2(n_442),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_589),
.B(n_459),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_588),
.A2(n_401),
.B1(n_450),
.B2(n_448),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_434),
.Y(n_635)
);

AOI22x1_ASAP7_75t_L g636 ( 
.A1(n_504),
.A2(n_421),
.B1(n_416),
.B2(n_418),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_523),
.B(n_450),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_531),
.B(n_437),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_531),
.B(n_437),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_532),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_416),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_596),
.A2(n_496),
.B(n_473),
.C(n_557),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_532),
.B(n_437),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_473),
.B(n_455),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_550),
.B(n_416),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_474),
.B(n_352),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_513),
.B(n_445),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_515),
.B(n_445),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_521),
.B(n_448),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_532),
.B(n_437),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_584),
.B(n_437),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_467),
.B(n_449),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_538),
.B(n_418),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_495),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_540),
.B(n_418),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_520),
.B(n_429),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_465),
.B(n_418),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_494),
.B(n_435),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_489),
.B(n_429),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_535),
.B(n_418),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_471),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_588),
.B(n_424),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_588),
.B(n_607),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_588),
.B(n_424),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_588),
.A2(n_454),
.B1(n_431),
.B2(n_447),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_561),
.B(n_451),
.C(n_435),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_584),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_544),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_588),
.B(n_424),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_607),
.B(n_424),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_558),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_607),
.B(n_424),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_607),
.B(n_431),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_607),
.B(n_431),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_482),
.B(n_403),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_558),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_542),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_484),
.B(n_403),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_548),
.A2(n_292),
.B1(n_264),
.B2(n_271),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_534),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_477),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_611),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_610),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_552),
.A2(n_454),
.B1(n_432),
.B2(n_447),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_511),
.B(n_432),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_536),
.B(n_411),
.Y(n_688)
);

NOR2x1p5_ASAP7_75t_L g689 ( 
.A(n_520),
.B(n_451),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_555),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_611),
.B(n_432),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_577),
.A2(n_454),
.B1(n_447),
.B2(n_444),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_492),
.B(n_411),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_548),
.B(n_502),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_548),
.B(n_438),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_611),
.B(n_438),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_477),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_509),
.B(n_438),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_611),
.B(n_441),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_611),
.B(n_441),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_498),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_611),
.A2(n_441),
.B1(n_444),
.B2(n_266),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_594),
.B(n_444),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_594),
.B(n_423),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_568),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_479),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_599),
.B(n_423),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_480),
.B(n_224),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_479),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_603),
.B(n_296),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_600),
.B(n_287),
.C(n_288),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_483),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_484),
.B(n_262),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_483),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_504),
.B(n_262),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_484),
.B(n_266),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_504),
.B(n_275),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_596),
.A2(n_481),
.B1(n_486),
.B2(n_568),
.Y(n_720)
);

NAND2x1p5_ASAP7_75t_L g721 ( 
.A(n_519),
.B(n_275),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_495),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_542),
.B(n_560),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_568),
.B(n_273),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_509),
.B(n_229),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_490),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_545),
.B(n_277),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_546),
.B(n_277),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_590),
.B(n_236),
.Y(n_729)
);

O2A1O1Ixp5_ASAP7_75t_L g730 ( 
.A1(n_546),
.A2(n_299),
.B(n_310),
.C(n_280),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_551),
.B(n_280),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_568),
.B(n_252),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_519),
.B(n_274),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_586),
.A2(n_274),
.B1(n_287),
.B2(n_288),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_490),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_554),
.B(n_272),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_500),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_551),
.B(n_278),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_498),
.A2(n_310),
.B1(n_189),
.B2(n_279),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_475),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_553),
.B(n_294),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_300),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_554),
.B(n_305),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_500),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_562),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_493),
.B(n_174),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_493),
.B(n_161),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_506),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_503),
.B(n_169),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_503),
.B(n_171),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_565),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_212),
.C(n_214),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_507),
.B(n_510),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_497),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_497),
.B(n_1),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_506),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_514),
.Y(n_757)
);

OAI221xp5_ASAP7_75t_L g758 ( 
.A1(n_507),
.A2(n_279),
.B1(n_220),
.B2(n_162),
.C(n_175),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_493),
.B(n_179),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_510),
.A2(n_220),
.B(n_175),
.C(n_307),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_469),
.A2(n_307),
.B(n_3),
.C(n_4),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_493),
.B(n_182),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_493),
.B(n_505),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_514),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_505),
.B(n_304),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_518),
.B(n_185),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_470),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_565),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_518),
.B(n_188),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_497),
.B(n_2),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_501),
.B(n_190),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_593),
.B(n_191),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_501),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_526),
.A2(n_446),
.B1(n_304),
.B2(n_311),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_571),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_571),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_740),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_640),
.B(n_526),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_617),
.B(n_593),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_740),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_740),
.Y(n_783)
);

BUFx4f_ASAP7_75t_L g784 ( 
.A(n_646),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_661),
.B(n_687),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_618),
.A2(n_602),
.B1(n_572),
.B2(n_573),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_622),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_SL g788 ( 
.A(n_725),
.B(n_199),
.C(n_194),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_501),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_617),
.A2(n_475),
.B1(n_602),
.B2(n_595),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_669),
.B(n_508),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_626),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_640),
.B(n_505),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_631),
.B(n_470),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_677),
.B(n_650),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_655),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_652),
.B(n_508),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_640),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_677),
.B(n_472),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_655),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_670),
.B(n_673),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_678),
.B(n_472),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_663),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_640),
.B(n_505),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_685),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_612),
.B(n_512),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_637),
.B(n_478),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_658),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_637),
.B(n_478),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_512),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_706),
.B(n_485),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_690),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_660),
.B(n_485),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_698),
.B(n_505),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_627),
.B(n_488),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_619),
.B(n_621),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_625),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_616),
.B(n_724),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_619),
.B(n_488),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_663),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_683),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_618),
.A2(n_475),
.B1(n_512),
.B2(n_547),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_661),
.B(n_547),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_614),
.B(n_547),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_689),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_687),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_621),
.B(n_491),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_R g828 ( 
.A(n_628),
.B(n_563),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_723),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_733),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_691),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_705),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_698),
.B(n_581),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_647),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_628),
.B(n_491),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_624),
.B(n_569),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_648),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_613),
.B(n_581),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_721),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_683),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_734),
.A2(n_575),
.B1(n_572),
.B2(n_573),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_733),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_700),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_649),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_653),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_707),
.B(n_569),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_644),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_623),
.B(n_581),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_754),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_699),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_713),
.B(n_595),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_684),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_708),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_662),
.B(n_595),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_634),
.B(n_753),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_735),
.Y(n_856)
);

INVx3_ASAP7_75t_SL g857 ( 
.A(n_736),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_720),
.B(n_581),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_744),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_703),
.B(n_597),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_742),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_679),
.B(n_597),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_754),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_SL g864 ( 
.A(n_682),
.B(n_597),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_756),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_708),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_764),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_773),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_711),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_773),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_703),
.B(n_562),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_564),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_729),
.B(n_732),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_767),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_711),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_732),
.B(n_575),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_SL g877 ( 
.A(n_681),
.B(n_244),
.C(n_210),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_751),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_714),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_656),
.A2(n_722),
.B(n_680),
.Y(n_880)
);

INVx5_ASAP7_75t_L g881 ( 
.A(n_770),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_695),
.B(n_581),
.Y(n_882)
);

AND2x6_ASAP7_75t_L g883 ( 
.A(n_664),
.B(n_666),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_714),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_668),
.B(n_578),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_680),
.A2(n_585),
.B(n_608),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_630),
.A2(n_585),
.B1(n_608),
.B2(n_605),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_703),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_716),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_629),
.B(n_609),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_703),
.B(n_564),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_703),
.B(n_567),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_688),
.B(n_567),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_710),
.A2(n_574),
.B1(n_605),
.B2(n_570),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_688),
.B(n_570),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_729),
.B(n_578),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_710),
.A2(n_574),
.B1(n_580),
.B2(n_582),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_726),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_642),
.B(n_609),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_737),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_737),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_675),
.B(n_579),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_748),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_748),
.B(n_580),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_757),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_R g908 ( 
.A(n_755),
.B(n_563),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_757),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_638),
.B(n_579),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_632),
.B(n_609),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_775),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_775),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_709),
.B(n_582),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_734),
.A2(n_604),
.B1(n_601),
.B2(n_598),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_738),
.A2(n_591),
.B1(n_604),
.B2(n_601),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_712),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_641),
.B(n_591),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_755),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_641),
.B(n_583),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_645),
.B(n_583),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_738),
.B(n_587),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_776),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_741),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_645),
.B(n_587),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_727),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_728),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_671),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_654),
.B(n_598),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_SL g931 ( 
.A1(n_758),
.A2(n_206),
.B1(n_201),
.B2(n_312),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_768),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_686),
.B(n_516),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_657),
.B(n_659),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_743),
.B(n_609),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_761),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_739),
.A2(n_609),
.B1(n_543),
.B2(n_541),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_745),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_639),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_731),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_715),
.A2(n_543),
.B(n_541),
.C(n_539),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_704),
.B(n_516),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_739),
.A2(n_539),
.B1(n_530),
.B2(n_527),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_715),
.Y(n_944)
);

INVx3_ASAP7_75t_SL g945 ( 
.A(n_718),
.Y(n_945)
);

BUFx4f_ASAP7_75t_L g946 ( 
.A(n_718),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_686),
.B(n_517),
.Y(n_947)
);

NOR2x2_ASAP7_75t_L g948 ( 
.A(n_774),
.B(n_2),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_643),
.B(n_530),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_752),
.A2(n_281),
.B1(n_225),
.B2(n_226),
.C(n_309),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_696),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_667),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_717),
.B(n_517),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_676),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_692),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_774),
.B(n_527),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_651),
.B(n_215),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_697),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_719),
.B(n_232),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_701),
.A2(n_446),
.B1(n_476),
.B2(n_308),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_702),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_808),
.B(n_749),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_778),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_817),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_785),
.B(n_672),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_873),
.A2(n_620),
.B(n_747),
.C(n_762),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_808),
.B(n_693),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_834),
.B(n_693),
.Y(n_968)
);

AND2x4_ASAP7_75t_SL g969 ( 
.A(n_782),
.B(n_694),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_795),
.A2(n_674),
.B(n_763),
.Y(n_970)
);

INVx6_ASAP7_75t_L g971 ( 
.A(n_782),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_795),
.A2(n_694),
.B(n_636),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_784),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_816),
.A2(n_772),
.B(n_750),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_782),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_783),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_R g977 ( 
.A(n_783),
.B(n_766),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_787),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_837),
.B(n_844),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_816),
.A2(n_769),
.B(n_759),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_889),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_919),
.A2(n_847),
.B(n_925),
.C(n_801),
.Y(n_982)
);

NOR2x1p5_ASAP7_75t_SL g983 ( 
.A(n_885),
.B(n_730),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_777),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_784),
.B(n_771),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_783),
.Y(n_986)
);

OR2x6_ASAP7_75t_SL g987 ( 
.A(n_948),
.B(n_234),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_830),
.B(n_746),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_959),
.B(n_760),
.C(n_746),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_845),
.A2(n_765),
.B(n_285),
.C(n_306),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_799),
.A2(n_765),
.B(n_284),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_798),
.B(n_476),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_886),
.A2(n_476),
.B(n_304),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_829),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_880),
.A2(n_476),
.B(n_304),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_944),
.B(n_238),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_842),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_832),
.B(n_3),
.Y(n_998)
);

AO31x2_ASAP7_75t_L g999 ( 
.A1(n_941),
.A2(n_446),
.A3(n_476),
.B(n_114),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_785),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_798),
.Y(n_1001)
);

BUFx8_ASAP7_75t_L g1002 ( 
.A(n_818),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_799),
.A2(n_239),
.B(n_302),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_781),
.A2(n_240),
.B1(n_245),
.B2(n_250),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_855),
.A2(n_257),
.B(n_298),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_874),
.Y(n_1006)
);

AO22x1_ASAP7_75t_L g1007 ( 
.A1(n_857),
.A2(n_290),
.B1(n_297),
.B2(n_295),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_826),
.B(n_6),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_781),
.A2(n_260),
.B(n_261),
.C(n_267),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_798),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_SL g1011 ( 
.A1(n_861),
.A2(n_270),
.B1(n_291),
.B2(n_293),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_789),
.B(n_6),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_860),
.A2(n_56),
.B(n_152),
.Y(n_1013)
);

AO21x1_ASAP7_75t_L g1014 ( 
.A1(n_855),
.A2(n_827),
.B(n_819),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_945),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_805),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_812),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_8),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_R g1019 ( 
.A(n_779),
.B(n_58),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_780),
.B(n_10),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_839),
.B(n_13),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_798),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_831),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_801),
.A2(n_13),
.B(n_14),
.C(n_18),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_938),
.B(n_14),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_850),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_825),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_779),
.B(n_80),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_792),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_863),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_864),
.B(n_90),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_934),
.A2(n_95),
.B(n_147),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_863),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_823),
.B(n_24),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_856),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_946),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_863),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_881),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_934),
.A2(n_827),
.B(n_819),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_859),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_823),
.B(n_30),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_843),
.B(n_31),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_889),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_878),
.B(n_939),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_835),
.A2(n_105),
.B(n_146),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_936),
.A2(n_446),
.B1(n_33),
.B2(n_35),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_917),
.B(n_32),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_878),
.B(n_33),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_828),
.A2(n_908),
.B(n_835),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_806),
.B(n_40),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_SL g1051 ( 
.A(n_881),
.B(n_40),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_807),
.B(n_42),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_862),
.B(n_49),
.C(n_446),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_936),
.A2(n_446),
.B(n_62),
.C(n_98),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_791),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_876),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_939),
.B(n_54),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_807),
.B(n_809),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_796),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_788),
.Y(n_1061)
);

BUFx5_ASAP7_75t_L g1062 ( 
.A(n_852),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_809),
.B(n_446),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_932),
.B(n_446),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_881),
.A2(n_794),
.B1(n_797),
.B2(n_802),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_868),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_868),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_794),
.B(n_927),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_878),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_867),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_875),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_901),
.A2(n_132),
.B(n_142),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_849),
.B(n_143),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_846),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_860),
.A2(n_893),
.B(n_871),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_846),
.B(n_851),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_928),
.B(n_940),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_898),
.B(n_810),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_957),
.B(n_950),
.C(n_877),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_813),
.B(n_935),
.C(n_838),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_923),
.B(n_952),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_813),
.B(n_848),
.C(n_802),
.Y(n_1083)
);

BUFx4f_ASAP7_75t_L g1084 ( 
.A(n_851),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_871),
.A2(n_893),
.B(n_872),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_904),
.B(n_836),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_910),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_815),
.B(n_954),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_824),
.A2(n_790),
.B(n_899),
.C(n_896),
.Y(n_1089)
);

BUFx8_ASAP7_75t_SL g1090 ( 
.A(n_870),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_910),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_815),
.A2(n_811),
.B(n_836),
.C(n_918),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_951),
.Y(n_1093)
);

INVx11_ASAP7_75t_L g1094 ( 
.A(n_852),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_884),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_955),
.B(n_958),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_961),
.B(n_895),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_922),
.B(n_924),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_895),
.B(n_897),
.Y(n_1099)
);

INVx3_ASAP7_75t_SL g1100 ( 
.A(n_949),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_897),
.B(n_933),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_911),
.A2(n_858),
.B(n_926),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_872),
.A2(n_894),
.B(n_914),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_920),
.A2(n_926),
.B(n_921),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_800),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_888),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_922),
.B(n_924),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_879),
.B(n_903),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_879),
.B(n_903),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_894),
.A2(n_914),
.B(n_811),
.Y(n_1110)
);

AOI221x1_ASAP7_75t_L g1111 ( 
.A1(n_1036),
.A2(n_882),
.B1(n_913),
.B2(n_920),
.C(n_921),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_974),
.A2(n_918),
.B(n_887),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_997),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_971),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_993),
.A2(n_953),
.B(n_906),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_973),
.B(n_951),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1039),
.A2(n_881),
.B(n_854),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_971),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1103),
.A2(n_916),
.B(n_930),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1110),
.A2(n_942),
.B(n_947),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1092),
.A2(n_1076),
.B(n_972),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1102),
.A2(n_892),
.B(n_793),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1073),
.A2(n_892),
.B(n_804),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1080),
.A2(n_931),
.B(n_929),
.C(n_822),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1099),
.A2(n_786),
.B1(n_951),
.B2(n_937),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_L g1126 ( 
.A(n_1001),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1057),
.B(n_909),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_SL g1128 ( 
.A(n_1061),
.B(n_960),
.C(n_814),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1013),
.A2(n_912),
.B(n_907),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1014),
.A2(n_833),
.B(n_956),
.Y(n_1130)
);

CKINVDCx11_ASAP7_75t_R g1131 ( 
.A(n_987),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_SL g1132 ( 
.A(n_964),
.B(n_951),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1085),
.A2(n_905),
.B(n_902),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1104),
.A2(n_900),
.B(n_890),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_984),
.Y(n_1135)
);

XOR2xp5_ASAP7_75t_L g1136 ( 
.A(n_994),
.B(n_1027),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_1090),
.Y(n_1137)
);

INVxp67_ASAP7_75t_SL g1138 ( 
.A(n_1079),
.Y(n_1138)
);

BUFx2_ASAP7_75t_R g1139 ( 
.A(n_1100),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1089),
.A2(n_949),
.B(n_943),
.C(n_915),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1059),
.A2(n_904),
.B(n_820),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_980),
.A2(n_904),
.B(n_821),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1069),
.A2(n_803),
.B(n_840),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_1053),
.A2(n_853),
.B(n_866),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_982),
.A2(n_1020),
.B(n_979),
.C(n_1042),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_970),
.A2(n_869),
.B(n_891),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1078),
.B(n_883),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_989),
.A2(n_841),
.B(n_883),
.C(n_852),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1101),
.A2(n_883),
.B(n_852),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1088),
.B(n_883),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1084),
.B(n_981),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1046),
.A2(n_1084),
.B1(n_967),
.B2(n_1077),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1063),
.A2(n_1066),
.B(n_998),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1097),
.A2(n_966),
.B(n_1049),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1034),
.B(n_996),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_963),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1041),
.B(n_1002),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1049),
.A2(n_1045),
.B(n_1032),
.Y(n_1158)
);

AO21x1_ASAP7_75t_L g1159 ( 
.A1(n_1046),
.A2(n_968),
.B(n_1024),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_1038),
.A2(n_1082),
.B1(n_991),
.B2(n_1055),
.C(n_1018),
.Y(n_1160)
);

AO22x2_ASAP7_75t_L g1161 ( 
.A1(n_1087),
.A2(n_962),
.B1(n_1072),
.B2(n_1106),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1096),
.A2(n_1095),
.A3(n_978),
.B(n_1029),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1074),
.A2(n_1086),
.B(n_1005),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_SL g1164 ( 
.A(n_1086),
.B(n_1001),
.Y(n_1164)
);

NAND2xp33_ASAP7_75t_R g1165 ( 
.A(n_977),
.B(n_1031),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1109),
.A2(n_1023),
.B(n_1071),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1041),
.A2(n_1034),
.B1(n_1008),
.B2(n_1016),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1017),
.A2(n_1035),
.B(n_1052),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_965),
.B(n_1006),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1026),
.A2(n_1040),
.B(n_985),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1083),
.A2(n_1081),
.B(n_1009),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1015),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_1041),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1011),
.B(n_1070),
.Y(n_1174)
);

AND2x2_ASAP7_75t_SL g1175 ( 
.A(n_1058),
.B(n_1091),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1056),
.B(n_1000),
.Y(n_1176)
);

NOR4xp25_ASAP7_75t_L g1177 ( 
.A(n_1048),
.B(n_1012),
.C(n_1021),
.D(n_1025),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_1098),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1003),
.A2(n_990),
.B(n_1054),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1043),
.A2(n_1044),
.B(n_1108),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_1060),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1001),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1051),
.A2(n_1086),
.B(n_1047),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_SL g1184 ( 
.A(n_1010),
.B(n_1022),
.Y(n_1184)
);

O2A1O1Ixp5_ASAP7_75t_L g1185 ( 
.A1(n_1004),
.A2(n_1050),
.B(n_1007),
.C(n_975),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1062),
.A2(n_992),
.B(n_975),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1010),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_969),
.A2(n_965),
.B(n_1093),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_999),
.A2(n_983),
.A3(n_1062),
.B(n_1094),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1075),
.B(n_976),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1062),
.A2(n_992),
.B(n_986),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1062),
.A2(n_976),
.B(n_986),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1030),
.B(n_1033),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1030),
.A2(n_1033),
.B(n_1068),
.Y(n_1194)
);

BUFx4_ASAP7_75t_SL g1195 ( 
.A(n_1008),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1030),
.A2(n_1033),
.B(n_1068),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1037),
.B(n_1068),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1010),
.B(n_1022),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_988),
.A2(n_1064),
.B(n_1062),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_999),
.A2(n_1011),
.B(n_1037),
.C(n_1067),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_999),
.A2(n_988),
.B(n_1022),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_988),
.A2(n_1037),
.B(n_1067),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1065),
.A2(n_1067),
.B(n_1008),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1065),
.A2(n_1075),
.B(n_1019),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1075),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1065),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_R g1207 ( 
.A(n_1028),
.B(n_1002),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1014),
.A2(n_1104),
.B(n_974),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1014),
.A2(n_1110),
.A3(n_1103),
.B(n_974),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1015),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1015),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_979),
.B(n_617),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_979),
.B(n_617),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1066),
.A2(n_816),
.B(n_873),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1084),
.B(n_873),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_SL g1225 ( 
.A1(n_1014),
.A2(n_1092),
.B(n_1069),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_963),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1041),
.B(n_1034),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1001),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_963),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1069),
.B(n_1099),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1080),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1099),
.A2(n_873),
.B1(n_618),
.B2(n_617),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_987),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1080),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_995),
.A2(n_993),
.B(n_1102),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_984),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1014),
.A2(n_1110),
.A3(n_1103),
.B(n_974),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_984),
.Y(n_1243)
);

OA22x2_ASAP7_75t_L g1244 ( 
.A1(n_1008),
.A2(n_542),
.B1(n_409),
.B2(n_434),
.Y(n_1244)
);

AO32x2_ASAP7_75t_L g1245 ( 
.A1(n_1066),
.A2(n_1036),
.A3(n_434),
.B1(n_1038),
.B2(n_845),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_974),
.A2(n_816),
.B(n_781),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1001),
.B(n_1010),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1014),
.A2(n_1110),
.A3(n_1103),
.B(n_974),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1057),
.B(n_829),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1080),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1092),
.A2(n_1099),
.B(n_816),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1092),
.A2(n_1099),
.B(n_816),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1039),
.A2(n_816),
.B(n_1110),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1080),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1080),
.A2(n_873),
.B(n_617),
.C(n_816),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_984),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1219),
.B(n_1220),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_SL g1259 ( 
.A(n_1175),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1166),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1236),
.A2(n_1238),
.B1(n_1235),
.B2(n_1250),
.C(n_1255),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1155),
.B(n_1176),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1229),
.A2(n_1240),
.B(n_1239),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1126),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1121),
.A2(n_1154),
.B(n_1209),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1187),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1211),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1216),
.A2(n_1227),
.B(n_1221),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1171),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1256),
.A2(n_1236),
.B(n_1145),
.C(n_1206),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1168),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1115),
.A2(n_1117),
.B(n_1129),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1244),
.A2(n_1167),
.B1(n_1138),
.B2(n_1157),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1230),
.A2(n_1254),
.B(n_1142),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1164),
.B(n_1202),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1135),
.Y(n_1277)
);

AO222x2_ASAP7_75t_L g1278 ( 
.A1(n_1195),
.A2(n_1131),
.B1(n_1245),
.B2(n_1157),
.C1(n_1173),
.C2(n_1237),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1249),
.B(n_1127),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1252),
.A2(n_1253),
.B(n_1246),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1231),
.A2(n_1234),
.B1(n_1223),
.B2(n_1171),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1144),
.A2(n_1153),
.B(n_1119),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1234),
.B(n_1178),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1152),
.B1(n_1124),
.B2(n_1140),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1184),
.B(n_1132),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1126),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1133),
.A2(n_1123),
.B(n_1146),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1207),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1122),
.A2(n_1201),
.B(n_1134),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1177),
.B(n_1185),
.C(n_1160),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1141),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1165),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1136),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1210),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1172),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1190),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1217),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1174),
.B(n_1210),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1162),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1120),
.A2(n_1130),
.B(n_1163),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1241),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1200),
.A2(n_1222),
.B(n_1111),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1199),
.B(n_1152),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1151),
.B(n_1169),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1187),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1162),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1112),
.A2(n_1186),
.B(n_1191),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1243),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1125),
.A2(n_1161),
.B1(n_1169),
.B2(n_1245),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1181),
.A2(n_1148),
.B(n_1150),
.Y(n_1310)
);

XOR2xp5_ASAP7_75t_L g1311 ( 
.A(n_1139),
.B(n_1161),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1257),
.B(n_1113),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1218),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1177),
.A2(n_1150),
.B(n_1125),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1192),
.A2(n_1183),
.B(n_1149),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1156),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1182),
.B(n_1232),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1149),
.A2(n_1147),
.B(n_1143),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1151),
.A2(n_1128),
.B1(n_1213),
.B2(n_1251),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_1212),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1170),
.A2(n_1179),
.B(n_1180),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1212),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1247),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1193),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1190),
.B(n_1197),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1194),
.A2(n_1196),
.B(n_1203),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1114),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1205),
.B(n_1204),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1118),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1179),
.A2(n_1245),
.B(n_1188),
.C(n_1116),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1197),
.B(n_1247),
.Y(n_1332)
);

OAI221xp5_ASAP7_75t_L g1333 ( 
.A1(n_1198),
.A2(n_1182),
.B1(n_1232),
.B2(n_1228),
.C(n_1233),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1215),
.A2(n_1242),
.B(n_1248),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1189),
.A2(n_1215),
.B(n_1242),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1189),
.B(n_1215),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1189),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1166),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1154),
.A2(n_1014),
.A3(n_1222),
.B(n_1158),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1231),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1168),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1155),
.B(n_987),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1168),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1171),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1236),
.A2(n_1244),
.B1(n_434),
.B2(n_1167),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1168),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1215),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1236),
.A2(n_873),
.B1(n_617),
.B2(n_618),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1139),
.B(n_487),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1121),
.A2(n_1154),
.B(n_1209),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1166),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1219),
.B(n_1220),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1235),
.A2(n_1238),
.B1(n_1255),
.B2(n_1250),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1235),
.A2(n_1238),
.B1(n_1255),
.B2(n_1250),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1137),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1126),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1235),
.B(n_873),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_SL g1359 ( 
.A(n_1139),
.B(n_487),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1171),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1154),
.A2(n_1158),
.B(n_1144),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1223),
.B(n_1043),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1168),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1168),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1121),
.A2(n_1154),
.B(n_1209),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1236),
.A2(n_873),
.B1(n_617),
.B2(n_618),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1168),
.Y(n_1369)
);

AOI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_617),
.B1(n_873),
.B2(n_434),
.C(n_618),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1236),
.A2(n_873),
.B(n_1238),
.C(n_1235),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1121),
.A2(n_1154),
.B(n_1209),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1219),
.B(n_1220),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1168),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1236),
.A2(n_618),
.B1(n_1244),
.B2(n_873),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1236),
.A2(n_618),
.B1(n_1244),
.B2(n_873),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1231),
.B(n_1167),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1249),
.B(n_1176),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1154),
.A2(n_1014),
.A3(n_1222),
.B(n_1158),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1208),
.A2(n_1226),
.B(n_1224),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1236),
.A2(n_617),
.B(n_873),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1312),
.Y(n_1383)
);

NOR2x1_ASAP7_75t_SL g1384 ( 
.A(n_1378),
.B(n_1284),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1330),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1358),
.A2(n_1382),
.B(n_1372),
.C(n_1355),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1370),
.A2(n_1368),
.B(n_1349),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1330),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1277),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1356),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1358),
.A2(n_1372),
.B(n_1354),
.C(n_1271),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1263),
.B(n_1298),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1353),
.B(n_1374),
.Y(n_1394)
);

NAND4xp25_ASAP7_75t_L g1395 ( 
.A(n_1261),
.B(n_1271),
.C(n_1345),
.D(n_1376),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1279),
.B(n_1313),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1376),
.A2(n_1377),
.B1(n_1345),
.B2(n_1274),
.Y(n_1397)
);

OAI22x1_ASAP7_75t_L g1398 ( 
.A1(n_1311),
.A2(n_1278),
.B1(n_1320),
.B2(n_1292),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1379),
.B(n_1301),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1270),
.A2(n_1360),
.B(n_1344),
.C(n_1377),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1290),
.B(n_1281),
.C(n_1363),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1274),
.A2(n_1259),
.B1(n_1309),
.B2(n_1295),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1326),
.B(n_1325),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1308),
.B(n_1304),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_1309),
.B1(n_1295),
.B2(n_1278),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1317),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1331),
.A2(n_1336),
.B(n_1321),
.C(n_1304),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1331),
.A2(n_1303),
.B(n_1336),
.C(n_1292),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1314),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1340),
.A2(n_1285),
.B1(n_1302),
.B2(n_1373),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1314),
.B(n_1347),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1285),
.A2(n_1329),
.B(n_1303),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1303),
.A2(n_1291),
.B(n_1300),
.C(n_1342),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1302),
.A2(n_1351),
.B1(n_1367),
.B2(n_1373),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1265),
.A2(n_1286),
.B(n_1347),
.C(n_1359),
.Y(n_1415)
);

OA22x2_ASAP7_75t_L g1416 ( 
.A1(n_1288),
.A2(n_1276),
.B1(n_1328),
.B2(n_1332),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1321),
.A2(n_1323),
.B1(n_1350),
.B2(n_1369),
.C(n_1365),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1282),
.B(n_1334),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1328),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1305),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1302),
.A2(n_1351),
.B1(n_1266),
.B2(n_1367),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1333),
.A2(n_1319),
.B(n_1316),
.C(n_1307),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1297),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1318),
.A2(n_1315),
.B(n_1267),
.C(n_1323),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1318),
.A2(n_1315),
.B(n_1351),
.C(n_1266),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1296),
.B(n_1276),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1272),
.Y(n_1427)
);

O2A1O1Ixp5_ASAP7_75t_L g1428 ( 
.A1(n_1341),
.A2(n_1343),
.B(n_1346),
.C(n_1375),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1305),
.B(n_1297),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1322),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1327),
.C(n_1289),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1357),
.A2(n_1310),
.B(n_1322),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1357),
.A2(n_1299),
.B(n_1306),
.C(n_1352),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1268),
.A2(n_1294),
.B1(n_1293),
.B2(n_1364),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1262),
.A2(n_1381),
.B(n_1264),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1324),
.B(n_1322),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1334),
.B(n_1268),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1260),
.A2(n_1338),
.B(n_1352),
.C(n_1362),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1260),
.A2(n_1338),
.B(n_1362),
.C(n_1335),
.Y(n_1439)
);

INVx5_ASAP7_75t_L g1440 ( 
.A(n_1306),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1337),
.B(n_1310),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1348),
.A2(n_1361),
.B(n_1366),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1339),
.B(n_1380),
.Y(n_1443)
);

OA22x2_ASAP7_75t_L g1444 ( 
.A1(n_1287),
.A2(n_1273),
.B1(n_1371),
.B2(n_1339),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1269),
.A2(n_1382),
.B(n_816),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1382),
.A2(n_816),
.B(n_1280),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1382),
.A2(n_816),
.B(n_1280),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1312),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1295),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_SL g1452 ( 
.A(n_1378),
.B(n_1231),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1378),
.B(n_1340),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1349),
.A2(n_1368),
.B1(n_1370),
.B2(n_1382),
.Y(n_1454)
);

AOI221x1_ASAP7_75t_SL g1455 ( 
.A1(n_1358),
.A2(n_1355),
.B1(n_1354),
.B2(n_184),
.C(n_192),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1378),
.B(n_1340),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1349),
.A2(n_1368),
.B1(n_1370),
.B2(n_1382),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1263),
.B(n_1298),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1382),
.A2(n_816),
.B(n_1280),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1409),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1443),
.B(n_1437),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1441),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1383),
.B(n_1450),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1430),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1435),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1427),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1414),
.B(n_1421),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1428),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1397),
.A2(n_1395),
.B1(n_1454),
.B2(n_1458),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1414),
.B(n_1421),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1389),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1411),
.B(n_1418),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1447),
.B(n_1457),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1431),
.B(n_1436),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1444),
.B(n_1407),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1454),
.A2(n_1458),
.B(n_1387),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1426),
.B(n_1413),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1445),
.A2(n_1410),
.B(n_1460),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1397),
.A2(n_1395),
.B1(n_1405),
.B2(n_1402),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1439),
.A2(n_1448),
.B(n_1446),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1426),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1438),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1406),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1410),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1422),
.A2(n_1402),
.B(n_1434),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1434),
.A2(n_1432),
.B(n_1433),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1404),
.B(n_1399),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1416),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1417),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1412),
.B(n_1453),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1393),
.B(n_1459),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1425),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1440),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1408),
.A2(n_1401),
.B(n_1386),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1392),
.A2(n_1449),
.B(n_1390),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1424),
.A2(n_1405),
.B(n_1400),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1464),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1486),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1465),
.Y(n_1505)
);

INVx3_ASAP7_75t_SL g1506 ( 
.A(n_1477),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1465),
.Y(n_1507)
);

OR2x2_ASAP7_75t_SL g1508 ( 
.A(n_1487),
.B(n_1385),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1472),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1472),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1470),
.A2(n_1398),
.B1(n_1455),
.B2(n_1394),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1462),
.B(n_1429),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1462),
.B(n_1396),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1462),
.B(n_1384),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_1394),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1467),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1480),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1468),
.B(n_1452),
.Y(n_1520)
);

AOI322xp5_ASAP7_75t_L g1521 ( 
.A1(n_1470),
.A2(n_1482),
.A3(n_1492),
.B1(n_1479),
.B2(n_1455),
.C1(n_1478),
.C2(n_1491),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1468),
.B(n_1456),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1461),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1468),
.B(n_1471),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1499),
.B(n_1420),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1415),
.C(n_1419),
.Y(n_1527)
);

OAI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1521),
.A2(n_1482),
.B(n_1471),
.C(n_1468),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1527),
.A2(n_1492),
.B1(n_1491),
.B2(n_1478),
.Y(n_1529)
);

AOI31xp33_ASAP7_75t_L g1530 ( 
.A1(n_1527),
.A2(n_1478),
.A3(n_1487),
.B(n_1471),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1508),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1504),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1523),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1523),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1506),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1513),
.A2(n_1488),
.B1(n_1497),
.B2(n_1500),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1512),
.A2(n_1497),
.B(n_1488),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1513),
.A2(n_1488),
.B1(n_1497),
.B2(n_1500),
.Y(n_1540)
);

AOI33xp33_ASAP7_75t_L g1541 ( 
.A1(n_1524),
.A2(n_1478),
.A3(n_1471),
.B1(n_1498),
.B2(n_1495),
.B3(n_1469),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1503),
.B(n_1423),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1526),
.A2(n_1485),
.B(n_1517),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1512),
.B(n_1480),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1503),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1506),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1506),
.Y(n_1548)
);

OAI21xp33_ASAP7_75t_L g1549 ( 
.A1(n_1521),
.A2(n_1481),
.B(n_1495),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1517),
.A2(n_1495),
.B1(n_1488),
.B2(n_1499),
.C(n_1497),
.Y(n_1550)
);

AND4x1_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1497),
.C(n_1469),
.D(n_1385),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1512),
.A2(n_1488),
.B1(n_1491),
.B2(n_1497),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1506),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1494),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1494),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1512),
.A2(n_1519),
.B1(n_1491),
.B2(n_1480),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1502),
.B(n_1490),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1526),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_L g1559 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1499),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1501),
.A2(n_1485),
.B(n_1476),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1519),
.A2(n_1493),
.B1(n_1481),
.B2(n_1480),
.Y(n_1563)
);

NOR2xp67_ASAP7_75t_SL g1564 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_1391),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1519),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1561),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1557),
.Y(n_1568)
);

AND4x1_ASAP7_75t_L g1569 ( 
.A(n_1537),
.B(n_1520),
.C(n_1516),
.D(n_1522),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1538),
.A2(n_1559),
.B(n_1509),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1550),
.B(n_1469),
.C(n_1498),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1538),
.A2(n_1510),
.B(n_1509),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1557),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1553),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1531),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1565),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1532),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1551),
.Y(n_1579)
);

INVx3_ASAP7_75t_SL g1580 ( 
.A(n_1547),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1530),
.A2(n_1483),
.B(n_1481),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1534),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1388),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1531),
.Y(n_1585)
);

NOR2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1559),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1543),
.Y(n_1589)
);

AO21x1_ASAP7_75t_SL g1590 ( 
.A1(n_1540),
.A2(n_1518),
.B(n_1525),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1553),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

AOI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1549),
.A2(n_1488),
.B(n_1500),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1541),
.B(n_1520),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_SL g1595 ( 
.A(n_1549),
.B(n_1451),
.C(n_1507),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1533),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1587),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1528),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1593),
.A2(n_1529),
.B1(n_1500),
.B2(n_1552),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1576),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1572),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1586),
.B(n_1580),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1579),
.A2(n_1556),
.B1(n_1500),
.B2(n_1489),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1570),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1594),
.B(n_1546),
.Y(n_1607)
);

AOI322xp5_ASAP7_75t_L g1608 ( 
.A1(n_1595),
.A2(n_1563),
.A3(n_1558),
.B1(n_1515),
.B2(n_1520),
.C1(n_1545),
.C2(n_1475),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1581),
.A2(n_1556),
.B(n_1545),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1568),
.B(n_1544),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1545),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1580),
.B(n_1547),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1575),
.B(n_1545),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1576),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1580),
.B(n_1536),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1578),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1578),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_1574),
.B(n_1548),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1570),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1592),
.B(n_1539),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1585),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1575),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1569),
.B(n_1562),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1567),
.Y(n_1628)
);

NAND4xp25_ASAP7_75t_L g1629 ( 
.A(n_1596),
.B(n_1507),
.C(n_1505),
.D(n_1466),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1569),
.B(n_1566),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1574),
.B(n_1564),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1602),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1598),
.B(n_1592),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1602),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1615),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1627),
.B(n_1574),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1627),
.B(n_1574),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1615),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1626),
.B(n_1564),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1625),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1577),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1603),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1600),
.B(n_1589),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1623),
.B(n_1494),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1618),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1601),
.A2(n_1607),
.B1(n_1606),
.B2(n_1621),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1597),
.B(n_1574),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1597),
.B(n_1591),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1614),
.B(n_1483),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1603),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1611),
.B(n_1591),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1613),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1604),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1605),
.A2(n_1584),
.B(n_1500),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1619),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1617),
.Y(n_1664)
);

CKINVDCx16_ASAP7_75t_R g1665 ( 
.A(n_1642),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1601),
.C(n_1608),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1645),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1599),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1637),
.B(n_1600),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1658),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1653),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1653),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1652),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1629),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1641),
.B(n_1608),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1641),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1635),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1635),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1636),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1638),
.B(n_1604),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1639),
.B(n_1616),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1651),
.A2(n_1590),
.B1(n_1617),
.B2(n_1629),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1634),
.B(n_1612),
.C(n_1610),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1659),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1657),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1672),
.Y(n_1691)
);

AOI322xp5_ASAP7_75t_L g1692 ( 
.A1(n_1679),
.A2(n_1665),
.A3(n_1687),
.B1(n_1678),
.B2(n_1689),
.C1(n_1667),
.C2(n_1666),
.Y(n_1692)
);

OAI32xp33_ASAP7_75t_L g1693 ( 
.A1(n_1665),
.A2(n_1639),
.A3(n_1641),
.B1(n_1606),
.B2(n_1621),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1672),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1676),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1676),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1649),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1686),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1671),
.B(n_1655),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1682),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1681),
.B(n_1636),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1682),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1686),
.B(n_1655),
.Y(n_1703)
);

AOI21xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1690),
.A2(n_1663),
.B(n_1657),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1690),
.A2(n_1663),
.B(n_1657),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1681),
.B(n_1640),
.Y(n_1706)
);

OAI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1680),
.A2(n_1678),
.B1(n_1654),
.B2(n_1609),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1688),
.A2(n_1664),
.B1(n_1647),
.B2(n_1644),
.Y(n_1708)
);

CKINVDCx14_ASAP7_75t_R g1709 ( 
.A(n_1685),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_R g1711 ( 
.A(n_1668),
.B(n_1616),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1698),
.B(n_1671),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1710),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1711),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1691),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1707),
.A2(n_1673),
.B1(n_1680),
.B2(n_1675),
.Y(n_1718)
);

BUFx12f_ASAP7_75t_L g1719 ( 
.A(n_1704),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1705),
.B(n_1674),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1694),
.Y(n_1721)
);

AOI32xp33_ASAP7_75t_L g1722 ( 
.A1(n_1718),
.A2(n_1692),
.A3(n_1710),
.B1(n_1706),
.B2(n_1701),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1716),
.A2(n_1699),
.B1(n_1677),
.B2(n_1674),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1677),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1712),
.A2(n_1697),
.B1(n_1669),
.B2(n_1611),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1719),
.A2(n_1708),
.B1(n_1688),
.B2(n_1644),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1714),
.A2(n_1706),
.B(n_1701),
.Y(n_1727)
);

NAND4xp75_ASAP7_75t_L g1728 ( 
.A(n_1720),
.B(n_1702),
.C(n_1700),
.D(n_1696),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1669),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1719),
.A2(n_1647),
.B1(n_1656),
.B2(n_1664),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1722),
.A2(n_1720),
.B1(n_1715),
.B2(n_1614),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1729),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1724),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1728),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1727),
.A2(n_1693),
.B(n_1715),
.C(n_1717),
.Y(n_1735)
);

OAI32xp33_ASAP7_75t_L g1736 ( 
.A1(n_1731),
.A2(n_1725),
.A3(n_1723),
.B1(n_1721),
.B2(n_1695),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1732),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1734),
.B(n_1726),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1734),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1735),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1740),
.B(n_1683),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1730),
.B1(n_1684),
.B2(n_1683),
.C(n_1656),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1741),
.A2(n_1684),
.B(n_1631),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1738),
.A2(n_1740),
.B1(n_1737),
.B2(n_1739),
.Y(n_1745)
);

NOR2x1_ASAP7_75t_L g1746 ( 
.A(n_1738),
.B(n_1640),
.Y(n_1746)
);

NOR2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1745),
.B(n_1736),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1746),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1744),
.A2(n_1650),
.B(n_1646),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1747),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1751),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1751),
.Y(n_1753)
);

INVx4_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

OAI22x1_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1748),
.B1(n_1742),
.B2(n_1743),
.Y(n_1755)
);

OR3x2_ASAP7_75t_L g1756 ( 
.A(n_1754),
.B(n_1755),
.C(n_1749),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1754),
.B(n_1646),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_R g1758 ( 
.A(n_1757),
.B(n_1606),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1756),
.A2(n_1661),
.B(n_1650),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1759),
.B(n_1661),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1758),
.B(n_1662),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1662),
.B1(n_1643),
.B2(n_1648),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1762),
.A2(n_1621),
.B1(n_1606),
.B2(n_1628),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1621),
.B(n_1620),
.C(n_1643),
.Y(n_1764)
);


endmodule