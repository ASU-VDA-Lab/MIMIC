module real_jpeg_32888_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g168 ( 
.A(n_0),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_0),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_0),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_1),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_105),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_105),
.B1(n_219),
.B2(n_223),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_1),
.A2(n_105),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_4),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_5),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_5),
.A2(n_174),
.B1(n_394),
.B2(n_399),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22x1_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_25),
.B1(n_90),
.B2(n_94),
.Y(n_89)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_25),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22x1_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_25),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_6),
.B(n_278),
.Y(n_277)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_6),
.A2(n_302),
.A3(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_6),
.B(n_143),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_7),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_54),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_9),
.A2(n_54),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_9),
.A2(n_54),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_375),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_245),
.B(n_373),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_208),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_17),
.B(n_209),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.C(n_188),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_18),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.Y(n_18)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_19),
.B(n_61),
.C(n_98),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_49),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_25),
.B(n_26),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_27),
.Y(n_26)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_25),
.B(n_196),
.Y(n_195)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_25),
.A2(n_272),
.A3(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_25),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_R g346 ( 
.A(n_25),
.B(n_77),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_25),
.B(n_180),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_26),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_29),
.B(n_50),
.Y(n_237)
);

NAND2x1p5_ASAP7_75t_L g385 ( 
.A(n_29),
.B(n_231),
.Y(n_385)
);

NOR2x1p5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_36),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_41),
.Y(n_196)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_45),
.Y(n_161)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NAND2x1p5_ASAP7_75t_L g384 ( 
.A(n_49),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_51),
.Y(n_154)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_97),
.B1(n_98),
.B2(n_145),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_61),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_88),
.B(n_89),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_62),
.B(n_89),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_62),
.B(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_62),
.B(n_254),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_77),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_87),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_80),
.Y(n_316)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2x1p5_ASAP7_75t_L g217 ( 
.A(n_88),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_88),
.B(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_88),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_88),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_89),
.B(n_293),
.Y(n_292)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_93),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_93),
.Y(n_274)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_96),
.Y(n_400)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_135),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_100),
.B(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_104),
.Y(n_243)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_136),
.Y(n_191)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_110),
.B(n_241),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_110),
.A2(n_241),
.B(n_387),
.Y(n_386)
);

AO21x2_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_117),
.B(n_126),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_112),
.Y(n_275)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_131),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_132),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_135),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_144),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g369 ( 
.A(n_146),
.B(n_189),
.Y(n_369)
);

XNOR2x1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_163),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_147),
.B(n_163),
.Y(n_227)
);

OAI31xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_151),
.A3(n_154),
.B(n_155),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_169),
.B(n_178),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_168),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_169),
.A2(n_205),
.B(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_172),
.Y(n_329)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_173),
.Y(n_328)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_173),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_178),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_178),
.B(n_321),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_179),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.C(n_197),
.Y(n_189)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_190),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_195),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_199),
.Y(n_350)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_200),
.B(n_322),
.Y(n_321)
);

BUFx4f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_205),
.B(n_325),
.Y(n_347)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_226),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_211),
.B(n_226),
.C(n_404),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_212),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_213),
.B(n_215),
.Y(n_388)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_214),
.A2(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_216),
.B(n_253),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_217),
.B(n_294),
.Y(n_332)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_227),
.B(n_229),
.C(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_238),
.Y(n_380)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_367),
.B(n_371),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_296),
.B(n_366),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_283),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_249),
.B(n_283),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_261),
.C(n_264),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_251),
.B(n_261),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_252),
.B(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_265),
.B(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_282),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_271),
.Y(n_295)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_291),
.C(n_295),
.Y(n_370)
);

OAI22x1_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_359),
.B(n_365),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_335),
.B(n_358),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_319),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_319),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_317),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_301),
.B1(n_317),
.B2(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_330),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_320),
.Y(n_362)
);

AND2x4_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_361),
.C(n_362),
.Y(n_360)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_344),
.B(n_357),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_338),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI21x1_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_348),
.B(n_356),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_347),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_363),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_370),
.Y(n_372)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_405),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_403),
.Y(n_377)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_389),
.B1(n_390),
.B2(n_402),
.Y(n_381)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

XOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_401),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_403),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);


endmodule