module fake_ariane_329_n_2016 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2016);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2016;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_50),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_117),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_49),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_28),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_116),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_57),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_171),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_41),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_133),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_12),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_86),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_68),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_103),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_136),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_56),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_56),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_34),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_162),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_51),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_139),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_159),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_74),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_130),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_27),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_106),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_147),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_57),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_82),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_45),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_152),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_156),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_43),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_71),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_35),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_28),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_43),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_37),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_4),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_115),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_123),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_88),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_104),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_174),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_164),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_24),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_59),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_26),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_122),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_141),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_99),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_97),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_148),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_127),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_121),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_178),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_158),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_41),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_160),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_89),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_55),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_128),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_93),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_79),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_9),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_113),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_188),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_75),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_169),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_19),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_177),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_107),
.Y(n_307)
);

BUFx8_ASAP7_75t_SL g308 ( 
.A(n_48),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_12),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_101),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_5),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_48),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_95),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_181),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_109),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_40),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_60),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_25),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_175),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_0),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_26),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_108),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_25),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_135),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_61),
.Y(n_329)
);

INVxp33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_114),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_44),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_45),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_16),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_60),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_6),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_31),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_38),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_145),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_55),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_102),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_24),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_98),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_144),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_62),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_13),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_29),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_168),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_63),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_49),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_70),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_73),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_92),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_80),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_110),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_173),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_77),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_35),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_180),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_23),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_76),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_34),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_65),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_62),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_125),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_53),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_8),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_87),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_193),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_22),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_5),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_126),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_8),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_1),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_151),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_189),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_21),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_46),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_16),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_84),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_170),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_91),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_185),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_190),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_54),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_30),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_229),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_375),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_268),
.B(n_1),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_378),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_201),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_211),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_219),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_308),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_220),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_209),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_204),
.B(n_7),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_221),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_252),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_206),
.B(n_7),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_195),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_270),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_268),
.B(n_9),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_195),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_270),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_289),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_295),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_10),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_270),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_209),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_195),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_195),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_240),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_388),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_388),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_246),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_264),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_388),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_241),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_290),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_304),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_317),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_196),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_258),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_318),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_196),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_289),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_319),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_213),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_197),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_197),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_261),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_198),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_198),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_337),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_199),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_286),
.B(n_10),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_199),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_203),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_316),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_328),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_253),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_200),
.B(n_11),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_253),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_203),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_278),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_204),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_278),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_334),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_356),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_376),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_294),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_205),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_205),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_208),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_277),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_334),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_213),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_224),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_294),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_210),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_202),
.B(n_11),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_343),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_277),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_347),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_277),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_277),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_207),
.B(n_13),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_301),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_286),
.B(n_14),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_286),
.B(n_15),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_301),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_210),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_212),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_392),
.A2(n_236),
.B(n_225),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_399),
.B(n_331),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_342),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_449),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_407),
.B(n_374),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_301),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_407),
.B(n_393),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_414),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_301),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_243),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_479),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_301),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_458),
.A2(n_302),
.B(n_281),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_480),
.A2(n_251),
.B(n_249),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_480),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_396),
.B(n_371),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_405),
.B(n_216),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_482),
.A2(n_283),
.B(n_255),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_397),
.B(n_371),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_413),
.B(n_371),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_485),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_433),
.Y(n_527)
);

AND2x2_ASAP7_75t_SL g528 ( 
.A(n_418),
.B(n_281),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_477),
.A2(n_302),
.B(n_293),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_488),
.B(n_291),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_310),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_457),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_459),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_461),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_326),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_401),
.B(n_353),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_408),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_416),
.B(n_371),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

AND3x2_ASAP7_75t_L g546 ( 
.A(n_395),
.B(n_330),
.C(n_370),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_431),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_432),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_410),
.B(n_371),
.Y(n_549)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_435),
.B(n_295),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_437),
.B(n_389),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_412),
.B(n_389),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_445),
.B(n_358),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_412),
.B(n_389),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_456),
.A2(n_373),
.B(n_372),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_490),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

NOR2x1_ASAP7_75t_L g566 ( 
.A(n_391),
.B(n_384),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_415),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_409),
.B(n_389),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_500),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_462),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_567),
.B(n_436),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_527),
.B(n_419),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_494),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_567),
.B(n_441),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_491),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_503),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_567),
.B(n_441),
.Y(n_583)
);

BUFx4f_ASAP7_75t_L g584 ( 
.A(n_549),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_517),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_497),
.Y(n_588)
);

BUFx6f_ASAP7_75t_SL g589 ( 
.A(n_567),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_503),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_499),
.B(n_374),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_494),
.B(n_385),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_567),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_513),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_503),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_513),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_494),
.B(n_273),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_527),
.B(n_419),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_547),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_539),
.B(n_424),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_517),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_539),
.B(n_424),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_539),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_556),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_517),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_556),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_547),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_517),
.Y(n_617)
);

BUFx4f_ASAP7_75t_L g618 ( 
.A(n_549),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_567),
.B(n_442),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_503),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_505),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_567),
.B(n_274),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_505),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_496),
.B(n_425),
.Y(n_625)
);

INVxp33_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_505),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_564),
.B(n_565),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_500),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_505),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_528),
.A2(n_440),
.B1(n_420),
.B2(n_469),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_525),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_505),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_564),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_398),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_498),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_512),
.B(n_425),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_321),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_547),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_526),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_528),
.A2(n_428),
.B1(n_377),
.B2(n_390),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_506),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_496),
.B(n_428),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_526),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_512),
.B(n_442),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_565),
.B(n_444),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_569),
.B(n_231),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_498),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_565),
.B(n_444),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_506),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_506),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_500),
.Y(n_660)
);

BUFx4f_ASAP7_75t_L g661 ( 
.A(n_549),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_569),
.B(n_570),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_528),
.B(n_520),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_512),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_509),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_547),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_547),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_551),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_500),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_509),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_528),
.B(n_446),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_549),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_569),
.B(n_231),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_528),
.A2(n_489),
.B1(n_476),
.B2(n_469),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_569),
.B(n_389),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_510),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_569),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_547),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_510),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_549),
.A2(n_489),
.B1(n_476),
.B2(n_468),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_511),
.Y(n_687)
);

BUFx4f_ASAP7_75t_L g688 ( 
.A(n_569),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_520),
.B(n_446),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_499),
.A2(n_448),
.B1(n_468),
.B2(n_451),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_511),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_511),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_570),
.Y(n_694)
);

BUFx10_ASAP7_75t_L g695 ( 
.A(n_569),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_511),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_515),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_501),
.B(n_448),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_570),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_570),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_501),
.B(n_451),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_554),
.B(n_452),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_501),
.B(n_452),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_515),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_547),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_501),
.B(n_544),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_501),
.B(n_460),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_460),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_502),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_569),
.B(n_568),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_499),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_515),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_499),
.A2(n_204),
.B1(n_232),
.B2(n_216),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_500),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_569),
.B(n_212),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_R g716 ( 
.A(n_546),
.B(n_403),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_500),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_515),
.Y(n_718)
);

AND2x6_ASAP7_75t_L g719 ( 
.A(n_568),
.B(n_232),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_519),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_628),
.B(n_568),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_584),
.A2(n_618),
.B1(n_661),
.B2(n_674),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_611),
.B(n_568),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_577),
.B(n_568),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_584),
.A2(n_568),
.B1(n_499),
.B2(n_507),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_572),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_612),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_612),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_584),
.A2(n_618),
.B1(n_661),
.B2(n_592),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_578),
.B(n_501),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_605),
.B(n_560),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_654),
.B(n_657),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_643),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_571),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_618),
.A2(n_499),
.B1(n_561),
.B2(n_507),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_578),
.B(n_499),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_643),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_625),
.B(n_651),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_694),
.B(n_592),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_686),
.B(n_563),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_666),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_563),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_592),
.B(n_563),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_637),
.B(n_563),
.C(n_562),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_592),
.B(n_560),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_661),
.B(n_541),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_592),
.B(n_542),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_592),
.B(n_542),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_699),
.B(n_542),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_699),
.B(n_542),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_581),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_599),
.B(n_562),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_700),
.B(n_495),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_688),
.B(n_541),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_607),
.B(n_495),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_595),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_673),
.A2(n_524),
.B1(n_523),
.B2(n_540),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_614),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_675),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_571),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_700),
.B(n_541),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_630),
.B(n_523),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_664),
.B(n_523),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_680),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_609),
.B(n_566),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_588),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_663),
.A2(n_531),
.B(n_543),
.C(n_540),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_664),
.B(n_523),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_689),
.B(n_698),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_707),
.B(n_702),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_708),
.B(n_566),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_523),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_674),
.A2(n_529),
.B(n_514),
.C(n_524),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_681),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_626),
.B(n_566),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_599),
.B(n_403),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_610),
.B(n_523),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_684),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_629),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_677),
.B(n_553),
.C(n_544),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_604),
.B(n_524),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_575),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_688),
.B(n_524),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_684),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_594),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_604),
.B(n_524),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_604),
.B(n_524),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_662),
.B(n_540),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_594),
.Y(n_794)
);

BUFx5_ASAP7_75t_L g795 ( 
.A(n_593),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_688),
.B(n_529),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_630),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_596),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_597),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_597),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_604),
.Y(n_802)
);

AND2x4_ASAP7_75t_SL g803 ( 
.A(n_575),
.B(n_404),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_603),
.B(n_544),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_601),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_616),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_616),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_711),
.B(n_529),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_595),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_685),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_632),
.B(n_653),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_L g813 ( 
.A1(n_690),
.A2(n_545),
.B(n_543),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_711),
.B(n_543),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_603),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_604),
.B(n_545),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_653),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_629),
.B(n_552),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_604),
.B(n_545),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_716),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_591),
.A2(n_333),
.B1(n_332),
.B2(n_215),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_614),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_701),
.B(n_703),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_660),
.Y(n_825)
);

BUFx8_ASAP7_75t_L g826 ( 
.A(n_701),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_719),
.B(n_548),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_624),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_719),
.B(n_548),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_634),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_703),
.B(n_531),
.C(n_548),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_719),
.B(n_591),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_685),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_636),
.B(n_546),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_593),
.B(n_529),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_719),
.B(n_557),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_706),
.B(n_544),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_719),
.B(n_557),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_636),
.B(n_423),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_706),
.B(n_557),
.C(n_533),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_634),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_693),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_591),
.B(n_660),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_719),
.B(n_518),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_648),
.B(n_553),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_640),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_719),
.B(n_518),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_595),
.B(n_535),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_679),
.B(n_518),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_640),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_679),
.B(n_518),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_642),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_642),
.Y(n_853)
);

OAI221xp5_ASAP7_75t_L g854 ( 
.A1(n_713),
.A2(n_535),
.B1(n_537),
.B2(n_555),
.C(n_332),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_679),
.B(n_692),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_622),
.A2(n_550),
.B1(n_559),
.B2(n_558),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_693),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_622),
.A2(n_550),
.B1(n_559),
.B2(n_558),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_692),
.B(n_537),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_647),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_692),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_696),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_670),
.B(n_553),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_670),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_593),
.B(n_552),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_714),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_714),
.B(n_553),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_717),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_717),
.B(n_555),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_662),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_585),
.B(n_550),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_585),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_587),
.B(n_429),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_576),
.A2(n_215),
.B1(n_333),
.B2(n_335),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_585),
.B(n_552),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_647),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_586),
.B(n_558),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_580),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_598),
.B(n_558),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_652),
.B(n_559),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_579),
.B(n_338),
.C(n_335),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_658),
.A2(n_514),
.B(n_559),
.C(n_533),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_583),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_710),
.A2(n_715),
.B(n_619),
.C(n_667),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_SL g885 ( 
.A(n_586),
.B(n_338),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_586),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_835),
.A2(n_676),
.B(n_655),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_835),
.A2(n_676),
.B(n_655),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_843),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_760),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_824),
.B(n_434),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_843),
.B(n_443),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_777),
.A2(n_659),
.B(n_658),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_732),
.B(n_662),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_773),
.B(n_662),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_774),
.B(n_665),
.C(n_659),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_662),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_839),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_723),
.B(n_598),
.Y(n_900)
);

AO21x2_ASAP7_75t_L g901 ( 
.A1(n_796),
.A2(n_809),
.B(n_817),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_757),
.B(n_662),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_757),
.B(n_662),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_839),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_796),
.A2(n_859),
.B(n_848),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_775),
.A2(n_645),
.B1(n_622),
.B2(n_454),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_SL g907 ( 
.A1(n_721),
.A2(n_665),
.B(n_652),
.C(n_582),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_823),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_812),
.A2(n_574),
.B(n_590),
.C(n_582),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_882),
.A2(n_671),
.B(n_669),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_774),
.B(n_608),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_738),
.B(n_608),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_884),
.A2(n_590),
.B(n_574),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_727),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_855),
.A2(n_682),
.B(n_598),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_731),
.A2(n_602),
.B(n_620),
.C(n_600),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_855),
.A2(n_695),
.B(n_682),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_812),
.A2(n_600),
.B(n_620),
.C(n_602),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_734),
.B(n_682),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_728),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_775),
.B(n_608),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_826),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_803),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_848),
.A2(n_695),
.B(n_589),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_859),
.A2(n_623),
.B(n_621),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_804),
.B(n_455),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_821),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_747),
.A2(n_623),
.B(n_621),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_869),
.B(n_613),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_756),
.A2(n_695),
.B(n_589),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_747),
.A2(n_589),
.B(n_613),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_733),
.A2(n_631),
.B(n_635),
.C(n_627),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_734),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_734),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_877),
.A2(n_617),
.B(n_613),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_815),
.B(n_465),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_730),
.B(n_466),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_865),
.A2(n_633),
.B(n_617),
.Y(n_938)
);

CKINVDCx10_ASAP7_75t_R g939 ( 
.A(n_826),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_730),
.B(n_837),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_734),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_731),
.A2(n_622),
.B1(n_645),
.B2(n_633),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_865),
.A2(n_633),
.B(n_617),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_879),
.A2(n_631),
.B(n_627),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_869),
.B(n_767),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_879),
.A2(n_639),
.B(n_635),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_762),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_875),
.A2(n_644),
.B(n_639),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_793),
.A2(n_649),
.B(n_644),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_780),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_849),
.A2(n_667),
.B(n_646),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_767),
.B(n_622),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_851),
.A2(n_667),
.B(n_646),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_724),
.B(n_622),
.Y(n_954)
);

OAI321xp33_ASAP7_75t_L g955 ( 
.A1(n_854),
.A2(n_534),
.A3(n_530),
.B1(n_271),
.B2(n_297),
.C(n_280),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_724),
.B(n_622),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_762),
.B(n_580),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_733),
.B(n_470),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_871),
.A2(n_646),
.B(n_649),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_737),
.A2(n_650),
.B(n_718),
.C(n_712),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_798),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_831),
.B(n_645),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_875),
.A2(n_650),
.B(n_709),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_880),
.A2(n_514),
.B(n_672),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_762),
.B(n_580),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_831),
.B(n_645),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_779),
.B(n_645),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_779),
.B(n_645),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_741),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_754),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_874),
.A2(n_341),
.B(n_339),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_725),
.A2(n_709),
.B(n_687),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_755),
.B(n_645),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_776),
.B(n_672),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_781),
.B(n_687),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_737),
.B(n_691),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_809),
.A2(n_829),
.B(n_827),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_761),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_786),
.B(n_474),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_836),
.A2(n_709),
.B(n_697),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_845),
.B(n_691),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_873),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_863),
.B(n_697),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_739),
.A2(n_718),
.B(n_712),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_838),
.A2(n_704),
.B(n_696),
.Y(n_985)
);

AO21x1_ASAP7_75t_L g986 ( 
.A1(n_820),
.A2(n_514),
.B(n_530),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_766),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_818),
.B(n_478),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_762),
.B(n_580),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_788),
.A2(n_720),
.B(n_704),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_867),
.B(n_533),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_783),
.B(n_580),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_746),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_840),
.B(n_533),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_750),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_783),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_783),
.B(n_606),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_753),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_783),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_763),
.A2(n_788),
.B(n_770),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_751),
.A2(n_720),
.B(n_615),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_798),
.B(n_481),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_744),
.B(n_606),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_735),
.A2(n_561),
.B1(n_516),
.B2(n_521),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_735),
.A2(n_705),
.B1(n_683),
.B2(n_668),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_868),
.B(n_606),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_840),
.A2(n_678),
.B1(n_683),
.B2(n_705),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_868),
.B(n_606),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_883),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_752),
.A2(n_615),
.B(n_606),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_769),
.A2(n_638),
.B(n_615),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_787),
.A2(n_638),
.B(n_615),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_740),
.B(n_533),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_881),
.B(n_533),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_825),
.B(n_534),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_790),
.A2(n_797),
.B(n_794),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_799),
.A2(n_638),
.B(n_615),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_813),
.B(n_504),
.Y(n_1019)
);

AO21x1_ASAP7_75t_L g1020 ( 
.A1(n_844),
.A2(n_847),
.B(n_745),
.Y(n_1020)
);

NAND3xp33_ASAP7_75t_L g1021 ( 
.A(n_759),
.B(n_341),
.C(n_339),
.Y(n_1021)
);

OAI22x1_ASAP7_75t_L g1022 ( 
.A1(n_834),
.A2(n_267),
.B1(n_309),
.B2(n_298),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_742),
.B(n_504),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_743),
.B(n_866),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_822),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_866),
.B(n_504),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_825),
.B(n_638),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_736),
.B(n_504),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_764),
.B(n_534),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_825),
.B(n_504),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_800),
.Y(n_1031)
);

BUFx4f_ASAP7_75t_L g1032 ( 
.A(n_864),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_771),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_795),
.B(n_678),
.Y(n_1034)
);

CKINVDCx10_ASAP7_75t_R g1035 ( 
.A(n_784),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_864),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_638),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_801),
.A2(n_683),
.B(n_668),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_805),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_806),
.A2(n_683),
.B(n_668),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_872),
.B(n_504),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_807),
.A2(n_705),
.B(n_683),
.C(n_668),
.Y(n_1042)
);

AO21x1_ASAP7_75t_L g1043 ( 
.A1(n_729),
.A2(n_522),
.B(n_519),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_808),
.A2(n_705),
.B(n_668),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_814),
.A2(n_678),
.B1(n_705),
.B2(n_344),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_872),
.B(n_678),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_816),
.A2(n_656),
.B(n_641),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_864),
.B(n_214),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_785),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_778),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_791),
.B(n_561),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_886),
.B(n_678),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_SL g1053 ( 
.A(n_768),
.B(n_232),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_886),
.B(n_226),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_878),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_828),
.A2(n_656),
.B(n_641),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_830),
.A2(n_233),
.B(n_230),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_765),
.A2(n_678),
.B(n_656),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_841),
.A2(n_656),
.B(n_641),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_846),
.B(n_678),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_850),
.B(n_532),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_852),
.A2(n_656),
.B(n_641),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_853),
.B(n_532),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_860),
.A2(n_641),
.B(n_561),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_876),
.A2(n_561),
.B(n_516),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_792),
.B(n_561),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_772),
.A2(n_538),
.B(n_536),
.C(n_532),
.Y(n_1067)
);

INVx11_ASAP7_75t_L g1068 ( 
.A(n_819),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_885),
.A2(n_235),
.B(n_234),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_878),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_758),
.B(n_532),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_819),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_945),
.B(n_722),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_SL g1074 ( 
.A(n_950),
.B(n_239),
.C(n_238),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_921),
.B(n_912),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_911),
.A2(n_905),
.B(n_929),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_892),
.B(n_536),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_958),
.B(n_247),
.C(n_242),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_905),
.A2(n_832),
.B(n_810),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1025),
.A2(n_722),
.B1(n_870),
.B2(n_748),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_902),
.B(n_758),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_896),
.A2(n_861),
.B(n_810),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_971),
.A2(n_903),
.B(n_898),
.C(n_961),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_891),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1054),
.A2(n_976),
.B(n_895),
.C(n_994),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_924),
.A2(n_861),
.B(n_878),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1017),
.B(n_782),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_SL g1088 ( 
.A(n_904),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1017),
.B(n_789),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1003),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_970),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_926),
.B(n_536),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_993),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_915),
.A2(n_878),
.B(n_749),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1064),
.A2(n_833),
.B(n_811),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_942),
.A2(n_955),
.B(n_918),
.C(n_909),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_920),
.A2(n_768),
.B1(n_802),
.B2(n_858),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_995),
.A2(n_802),
.B1(n_856),
.B2(n_857),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_917),
.A2(n_795),
.B(n_842),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_998),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_SL g1101 ( 
.A1(n_952),
.A2(n_862),
.B(n_561),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_981),
.B(n_795),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_937),
.B(n_795),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_795),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1002),
.B(n_988),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_937),
.A2(n_936),
.B1(n_979),
.B2(n_940),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_954),
.A2(n_795),
.B(n_280),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_975),
.B(n_1031),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_956),
.A2(n_297),
.B(n_271),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_899),
.B(n_927),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_914),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1039),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1034),
.A2(n_516),
.B(n_492),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_906),
.A2(n_538),
.B1(n_536),
.B2(n_263),
.Y(n_1114)
);

OAI22x1_ASAP7_75t_L g1115 ( 
.A1(n_893),
.A2(n_538),
.B1(n_262),
.B2(n_313),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1029),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_969),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_887),
.A2(n_492),
.B(n_516),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_887),
.A2(n_492),
.B(n_516),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_893),
.B(n_923),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_978),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1032),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1057),
.A2(n_538),
.B(n_522),
.C(n_519),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_940),
.B(n_214),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1008),
.A2(n_522),
.B(n_519),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_987),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_888),
.A2(n_492),
.B(n_521),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_890),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_983),
.B(n_492),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1033),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_982),
.A2(n_1022),
.B1(n_1021),
.B2(n_923),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_1068),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_933),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_889),
.B(n_217),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1000),
.B(n_492),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1050),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1064),
.A2(n_521),
.B(n_516),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1010),
.B(n_922),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_939),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_960),
.A2(n_522),
.B(n_493),
.C(n_516),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_964),
.A2(n_521),
.B(n_492),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_933),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_SL g1143 ( 
.A(n_1069),
.B(n_257),
.C(n_327),
.Y(n_1143)
);

INVx3_ASAP7_75t_SL g1144 ( 
.A(n_933),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1061),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1000),
.B(n_521),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_SL g1147 ( 
.A(n_1048),
.B(n_322),
.C(n_320),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_889),
.B(n_250),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1011),
.A2(n_1013),
.B(n_1012),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1032),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_908),
.B(n_254),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1016),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_888),
.A2(n_521),
.B(n_340),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1072),
.A2(n_260),
.B1(n_349),
.B2(n_383),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_977),
.A2(n_521),
.B(n_245),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_977),
.A2(n_244),
.B(n_222),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1035),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_L g1159 ( 
.A(n_1055),
.B(n_276),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1065),
.A2(n_894),
.B(n_1011),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1030),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_941),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_999),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1063),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_962),
.A2(n_348),
.B(n_311),
.C(n_324),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_1007),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_931),
.A2(n_315),
.B(n_314),
.Y(n_1167)
);

AO32x1_ASAP7_75t_L g1168 ( 
.A1(n_1006),
.A2(n_493),
.A3(n_498),
.B1(n_18),
.B2(n_21),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_941),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1049),
.B(n_312),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_941),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1026),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_999),
.Y(n_1173)
);

BUFx8_ASAP7_75t_SL g1174 ( 
.A(n_947),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_966),
.A2(n_365),
.B(n_323),
.C(n_352),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_947),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1043),
.A2(n_493),
.B(n_502),
.C(n_18),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_SL g1178 ( 
.A(n_947),
.B(n_382),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_934),
.B(n_1036),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_996),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_991),
.B(n_502),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_996),
.B(n_217),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1041),
.Y(n_1183)
);

INVx3_ASAP7_75t_SL g1184 ( 
.A(n_996),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_935),
.A2(n_223),
.B(n_227),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1014),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1036),
.B(n_498),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_910),
.A2(n_305),
.B(n_237),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_972),
.A2(n_306),
.B(n_228),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_897),
.A2(n_218),
.B1(n_344),
.B2(n_387),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_R g1191 ( 
.A(n_1053),
.B(n_218),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1028),
.A2(n_345),
.B1(n_387),
.B2(n_366),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_967),
.B(n_502),
.Y(n_1193)
);

CKINVDCx14_ASAP7_75t_R g1194 ( 
.A(n_1055),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_345),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1024),
.B(n_366),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_972),
.A2(n_1013),
.B(n_1012),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_968),
.B(n_1009),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_913),
.A2(n_15),
.B(n_17),
.C(n_22),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_SL g1201 ( 
.A(n_932),
.B(n_354),
.C(n_275),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1018),
.A2(n_300),
.B(n_259),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_990),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1015),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1037),
.B(n_498),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1023),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1018),
.A2(n_303),
.B(n_265),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_957),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1020),
.A2(n_498),
.B1(n_502),
.B2(n_380),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_965),
.B(n_248),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_901),
.Y(n_1211)
);

OR2x6_ASAP7_75t_SL g1212 ( 
.A(n_1019),
.B(n_266),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_925),
.B(n_502),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_984),
.B(n_948),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1071),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1005),
.A2(n_502),
.B1(n_325),
.B2(n_379),
.Y(n_1216)
);

OA22x2_ASAP7_75t_L g1217 ( 
.A1(n_1045),
.A2(n_362),
.B1(n_269),
.B2(n_272),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_916),
.B(n_502),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_901),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1047),
.B(n_498),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1038),
.A2(n_307),
.B(n_282),
.Y(n_1221)
);

BUFx2_ASAP7_75t_SL g1222 ( 
.A(n_989),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1065),
.A2(n_299),
.B(n_279),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_963),
.B(n_502),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_992),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1051),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1066),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1038),
.A2(n_498),
.B(n_368),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1004),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1105),
.B(n_17),
.Y(n_1230)
);

AO32x2_ASAP7_75t_L g1231 ( 
.A1(n_1211),
.A2(n_986),
.A3(n_907),
.B1(n_1042),
.B2(n_1044),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1139),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1106),
.B(n_997),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1211),
.A2(n_1040),
.A3(n_1044),
.B(n_973),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1078),
.A2(n_1067),
.B(n_1027),
.C(n_900),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_L g1236 ( 
.A1(n_1223),
.A2(n_919),
.B(n_1040),
.C(n_930),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1200),
.A2(n_1046),
.B(n_1052),
.C(n_928),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1191),
.B(n_963),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1108),
.A2(n_943),
.B1(n_938),
.B2(n_1060),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1132),
.B(n_944),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1223),
.A2(n_951),
.B(n_953),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1092),
.B(n_23),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1103),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1104),
.A2(n_1058),
.B(n_1059),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_1062),
.B(n_1059),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1076),
.A2(n_985),
.B(n_951),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1075),
.A2(n_1062),
.B(n_1056),
.Y(n_1248)
);

AOI31xp67_ASAP7_75t_L g1249 ( 
.A1(n_1203),
.A2(n_1001),
.A3(n_985),
.B(n_1056),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1116),
.B(n_1108),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1206),
.B(n_1047),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1074),
.A2(n_1192),
.B(n_1170),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1075),
.A2(n_949),
.B(n_946),
.C(n_980),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1077),
.B(n_959),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1122),
.B(n_953),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1161),
.B(n_1229),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1162),
.B(n_959),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1149),
.A2(n_231),
.B(n_256),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1149),
.A2(n_231),
.B(n_256),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1111),
.B(n_30),
.Y(n_1260)
);

AO21x2_ASAP7_75t_L g1261 ( 
.A1(n_1101),
.A2(n_231),
.B(n_256),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1102),
.A2(n_1146),
.B(n_1135),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1088),
.Y(n_1263)
);

BUFx5_ASAP7_75t_L g1264 ( 
.A(n_1205),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1102),
.A2(n_364),
.B(n_360),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1228),
.A2(n_1198),
.A3(n_1214),
.B(n_1226),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1166),
.B(n_31),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1095),
.A2(n_231),
.B(n_256),
.Y(n_1268)
);

AOI221x1_ASAP7_75t_L g1269 ( 
.A1(n_1228),
.A2(n_231),
.B1(n_256),
.B2(n_36),
.C(n_37),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1085),
.A2(n_357),
.B(n_355),
.C(n_351),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1083),
.A2(n_350),
.B(n_346),
.C(n_296),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1073),
.A2(n_292),
.B1(n_288),
.B2(n_256),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1073),
.A2(n_256),
.B(n_231),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1160),
.A2(n_1099),
.B(n_1086),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1079),
.A2(n_256),
.B(n_90),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1199),
.A2(n_32),
.B(n_33),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1080),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1183),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1212),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1162),
.B(n_131),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1080),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1135),
.A2(n_140),
.B(n_192),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1146),
.A2(n_119),
.B(n_191),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1122),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1124),
.A2(n_1112),
.B1(n_1100),
.B2(n_1093),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1094),
.A2(n_105),
.B(n_183),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1082),
.A2(n_100),
.B(n_172),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1081),
.A2(n_85),
.B(n_166),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1128),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1165),
.A2(n_58),
.B(n_59),
.C(n_61),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1081),
.A2(n_64),
.B(n_69),
.Y(n_1291)
);

AOI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1217),
.A2(n_72),
.B(n_78),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1121),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1192),
.A2(n_83),
.B1(n_142),
.B2(n_149),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1126),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1129),
.A2(n_1107),
.B(n_1089),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1137),
.A2(n_153),
.B(n_155),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1174),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1122),
.B(n_194),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1224),
.A2(n_1119),
.B(n_1118),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1091),
.A2(n_1217),
.B1(n_1190),
.B2(n_1115),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1120),
.B(n_1158),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1130),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1190),
.B2(n_1159),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1150),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1117),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1175),
.A2(n_1096),
.B(n_1134),
.C(n_1151),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1194),
.B(n_1132),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1150),
.Y(n_1310)
);

NAND2xp33_ASAP7_75t_L g1311 ( 
.A(n_1150),
.B(n_1110),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1131),
.B(n_1090),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1090),
.B(n_1147),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1129),
.A2(n_1087),
.B(n_1089),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1090),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1162),
.B(n_1179),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1144),
.B(n_1184),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1214),
.A2(n_1227),
.A3(n_1156),
.B(n_1113),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1172),
.B(n_1164),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1137),
.A2(n_1127),
.B(n_1154),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1136),
.B(n_1169),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1186),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1097),
.B(n_1162),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1171),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1163),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1087),
.A2(n_1213),
.B(n_1220),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1143),
.A2(n_1188),
.B(n_1157),
.C(n_1209),
.Y(n_1327)
);

AOI221xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1189),
.A2(n_1145),
.B1(n_1185),
.B2(n_1196),
.C(n_1216),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1176),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1213),
.A2(n_1220),
.B(n_1181),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1141),
.A2(n_1218),
.B(n_1219),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1195),
.B(n_1215),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1220),
.A2(n_1181),
.B(n_1193),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1193),
.A2(n_1109),
.B(n_1218),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1133),
.B(n_1142),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_SL g1336 ( 
.A1(n_1182),
.A2(n_1201),
.B(n_1098),
.C(n_1210),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1178),
.A2(n_1177),
.B(n_1125),
.C(n_1221),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1219),
.A2(n_1140),
.B(n_1098),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1123),
.A2(n_1216),
.B(n_1207),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1168),
.A2(n_1205),
.B(n_1202),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1167),
.A2(n_1173),
.B(n_1180),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1114),
.A2(n_1225),
.A3(n_1168),
.B(n_1197),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1208),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1114),
.A2(n_1225),
.A3(n_1168),
.B(n_1197),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1222),
.A2(n_1208),
.A3(n_1204),
.B(n_1187),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1179),
.A2(n_1208),
.B(n_1187),
.C(n_1176),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1176),
.A2(n_945),
.B(n_905),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1155),
.A2(n_945),
.B(n_589),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1105),
.A2(n_775),
.B(n_774),
.C(n_732),
.Y(n_1349)
);

INVx5_ASAP7_75t_L g1350 ( 
.A(n_1174),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1105),
.A2(n_839),
.B1(n_926),
.B2(n_604),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1105),
.A2(n_812),
.B(n_732),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1128),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1105),
.A2(n_812),
.B1(n_636),
.B2(n_732),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1111),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1174),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1359)
);

NOR2xp67_ASAP7_75t_L g1360 ( 
.A(n_1162),
.B(n_1197),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1105),
.A2(n_732),
.B1(n_812),
.B2(n_945),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1122),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1105),
.B(n_732),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1365)
);

NOR2x1p5_ASAP7_75t_SL g1366 ( 
.A(n_1203),
.B(n_990),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1075),
.A2(n_732),
.B(n_945),
.C(n_903),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1105),
.B(n_892),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1105),
.B(n_892),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1075),
.A2(n_732),
.B(n_945),
.C(n_903),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1139),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1160),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1105),
.A2(n_839),
.B1(n_926),
.B2(n_604),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1105),
.A2(n_775),
.B(n_774),
.C(n_732),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1149),
.A2(n_1198),
.B(n_1095),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1229),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1084),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1104),
.A2(n_688),
.B(n_945),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_SL g1386 ( 
.A(n_1110),
.B(n_1191),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1105),
.B(n_892),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1139),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1122),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1084),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1105),
.B(n_732),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1232),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1354),
.A2(n_1377),
.B1(n_1351),
.B2(n_1361),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1353),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1383),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1354),
.A2(n_1276),
.B1(n_1281),
.B2(n_1277),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1363),
.A2(n_1391),
.B1(n_1304),
.B2(n_1277),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1355),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1244),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1375),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1358),
.Y(n_1401)
);

BUFx10_ASAP7_75t_L g1402 ( 
.A(n_1388),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1298),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1324),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1386),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1369),
.B(n_1373),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1352),
.A2(n_1379),
.B1(n_1349),
.B2(n_1252),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1315),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1352),
.A2(n_1252),
.B1(n_1304),
.B2(n_1230),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1281),
.A2(n_1267),
.B1(n_1387),
.B2(n_1308),
.Y(n_1410)
);

CKINVDCx6p67_ASAP7_75t_R g1411 ( 
.A(n_1298),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1307),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1312),
.A2(n_1233),
.B1(n_1242),
.B2(n_1273),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1317),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1279),
.A2(n_1301),
.B1(n_1292),
.B2(n_1332),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1298),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1272),
.A2(n_1270),
.B1(n_1289),
.B2(n_1327),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1272),
.A2(n_1278),
.B1(n_1285),
.B2(n_1250),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1273),
.A2(n_1339),
.B1(n_1283),
.B2(n_1322),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1350),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1293),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1384),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1350),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1260),
.A2(n_1337),
.B1(n_1271),
.B2(n_1348),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1339),
.A2(n_1283),
.B1(n_1319),
.B2(n_1297),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1295),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1297),
.A2(n_1256),
.B1(n_1383),
.B2(n_1390),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1347),
.B2(n_1313),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1325),
.Y(n_1429)
);

INVx4_ASAP7_75t_SL g1430 ( 
.A(n_1345),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1238),
.A2(n_1323),
.B1(n_1321),
.B2(n_1343),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1305),
.A2(n_1254),
.B1(n_1302),
.B2(n_1241),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1335),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1350),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1347),
.A2(n_1290),
.B1(n_1309),
.B2(n_1240),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1311),
.A2(n_1336),
.B1(n_1264),
.B2(n_1362),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1269),
.A2(n_1326),
.B1(n_1316),
.B2(n_1362),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1329),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1241),
.A2(n_1264),
.B1(n_1320),
.B2(n_1251),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1264),
.A2(n_1320),
.B1(n_1243),
.B2(n_1262),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_L g1441 ( 
.A(n_1315),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1345),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1240),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1345),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1284),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1310),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1310),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1266),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1310),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1284),
.B(n_1389),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1264),
.Y(n_1451)
);

NAND2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1360),
.B(n_1306),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1264),
.A2(n_1314),
.B1(n_1340),
.B2(n_1389),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1306),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1239),
.A2(n_1333),
.B1(n_1261),
.B2(n_1282),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1261),
.A2(n_1341),
.B1(n_1330),
.B2(n_1291),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1265),
.A2(n_1255),
.B(n_1247),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1299),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1338),
.A2(n_1288),
.B1(n_1328),
.B2(n_1357),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1235),
.A2(n_1360),
.B1(n_1381),
.B2(n_1364),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1346),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1356),
.A2(n_1385),
.B1(n_1372),
.B2(n_1367),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1342),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1368),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1280),
.A2(n_1248),
.B1(n_1296),
.B2(n_1257),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1342),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1374),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1344),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1344),
.B(n_1280),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1328),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1376),
.Y(n_1471)
);

BUFx10_ASAP7_75t_L g1472 ( 
.A(n_1344),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1334),
.A2(n_1247),
.B1(n_1245),
.B2(n_1287),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1246),
.A2(n_1237),
.B1(n_1286),
.B2(n_1376),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1253),
.A2(n_1231),
.B1(n_1318),
.B2(n_1236),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1300),
.A2(n_1331),
.B1(n_1275),
.B2(n_1259),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1274),
.B(n_1268),
.Y(n_1477)
);

INVx6_ASAP7_75t_L g1478 ( 
.A(n_1366),
.Y(n_1478)
);

CKINVDCx6p67_ASAP7_75t_R g1479 ( 
.A(n_1231),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1258),
.A2(n_1365),
.B1(n_1380),
.B2(n_1378),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1234),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1359),
.A2(n_1370),
.B1(n_1371),
.B2(n_1382),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1231),
.A2(n_1354),
.B1(n_1105),
.B2(n_1391),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1249),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1234),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1244),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1244),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1298),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1266),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1314),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1375),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1354),
.A2(n_1105),
.B1(n_599),
.B2(n_603),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1310),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1363),
.A2(n_1391),
.B(n_1354),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1383),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1316),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1375),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1504)
);

OAI21xp33_ASAP7_75t_L g1505 ( 
.A1(n_1352),
.A2(n_1354),
.B(n_1349),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1363),
.B(n_1391),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1354),
.A2(n_1105),
.B1(n_599),
.B2(n_603),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1244),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1263),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1354),
.A2(n_1105),
.B1(n_599),
.B2(n_603),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1353),
.Y(n_1511)
);

CKINVDCx6p67_ASAP7_75t_R g1512 ( 
.A(n_1298),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1363),
.B(n_1391),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1354),
.A2(n_775),
.B1(n_1361),
.B2(n_812),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1244),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1244),
.Y(n_1516)
);

BUFx12f_ASAP7_75t_L g1517 ( 
.A(n_1375),
.Y(n_1517)
);

BUFx8_ASAP7_75t_L g1518 ( 
.A(n_1232),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1232),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1361),
.A2(n_839),
.B1(n_812),
.B2(n_423),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1266),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1354),
.A2(n_839),
.B1(n_604),
.B2(n_1105),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1361),
.A2(n_839),
.B1(n_812),
.B2(n_423),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1353),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1263),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1383),
.B(n_1310),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1244),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1354),
.A2(n_839),
.B1(n_604),
.B2(n_1105),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1399),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1395),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1448),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1430),
.B(n_1442),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1506),
.B(n_1513),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1422),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1416),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1394),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1492),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1478),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1524),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1443),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1397),
.A2(n_1526),
.B1(n_1521),
.B2(n_1396),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1495),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1488),
.A2(n_1494),
.B1(n_1493),
.B2(n_1491),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1447),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1495),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1449),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1499),
.B(n_1398),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1474),
.A2(n_1473),
.B(n_1462),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1473),
.A2(n_1462),
.B(n_1456),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1486),
.Y(n_1557)
);

AND2x2_ASAP7_75t_SL g1558 ( 
.A(n_1396),
.B(n_1488),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1505),
.B(n_1500),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1487),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1404),
.B(n_1489),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1508),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1515),
.B(n_1516),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1531),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1443),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

BUFx2_ASAP7_75t_SL g1567 ( 
.A(n_1490),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1421),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1426),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1491),
.A2(n_1514),
.B1(n_1493),
.B2(n_1504),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1520),
.B(n_1522),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1481),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1407),
.A2(n_1523),
.B(n_1527),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1430),
.B(n_1444),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1412),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1451),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1468),
.B(n_1433),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1511),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1392),
.Y(n_1579)
);

AO21x2_ASAP7_75t_L g1580 ( 
.A1(n_1475),
.A2(n_1465),
.B(n_1469),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1463),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1466),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1432),
.B(n_1406),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1529),
.B(n_1528),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1438),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1432),
.B(n_1439),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1439),
.B(n_1472),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1485),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1423),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1472),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1455),
.A2(n_1453),
.B(n_1457),
.Y(n_1591)
);

AOI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1424),
.A2(n_1460),
.B(n_1464),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1471),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1429),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1403),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1451),
.B(n_1409),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1441),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1456),
.A2(n_1482),
.B(n_1477),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1521),
.A2(n_1526),
.B1(n_1483),
.B2(n_1494),
.Y(n_1599)
);

AO31x2_ASAP7_75t_L g1600 ( 
.A1(n_1417),
.A2(n_1467),
.A3(n_1435),
.B(n_1410),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1471),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1482),
.A2(n_1477),
.B(n_1455),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1490),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1414),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1450),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1471),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1484),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1497),
.A2(n_1507),
.B1(n_1510),
.B2(n_1436),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1430),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1461),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1453),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1425),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1465),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1470),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1480),
.A2(n_1476),
.B(n_1440),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1445),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1476),
.A2(n_1480),
.B(n_1440),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1425),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1419),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1437),
.A2(n_1419),
.B(n_1427),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1501),
.B(n_1514),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1427),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_R g1623 ( 
.A(n_1519),
.B(n_1517),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1437),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1413),
.B(n_1504),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1431),
.A2(n_1452),
.B(n_1502),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1413),
.B(n_1501),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1458),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1498),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1459),
.A2(n_1428),
.B(n_1418),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1459),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1405),
.Y(n_1632)
);

AO21x2_ASAP7_75t_L g1633 ( 
.A1(n_1428),
.A2(n_1418),
.B(n_1415),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1509),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1502),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1454),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1434),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1446),
.B(n_1393),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1411),
.Y(n_1639)
);

CKINVDCx8_ASAP7_75t_R g1640 ( 
.A(n_1503),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1420),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1557),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1628),
.B(n_1415),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1573),
.B(n_1533),
.C(n_1525),
.Y(n_1644)
);

NOR2xp67_ASAP7_75t_L g1645 ( 
.A(n_1614),
.B(n_1530),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1557),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1599),
.A2(n_1512),
.B(n_1408),
.C(n_1496),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1571),
.A2(n_1400),
.B(n_1408),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1623),
.B(n_1401),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1605),
.B(n_1402),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1558),
.B(n_1402),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1548),
.A2(n_1401),
.B(n_1518),
.C(n_1625),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1564),
.B(n_1518),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1558),
.A2(n_1550),
.B1(n_1570),
.B2(n_1621),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1583),
.Y(n_1655)
);

AO21x2_ASAP7_75t_L g1656 ( 
.A1(n_1612),
.A2(n_1618),
.B(n_1620),
.Y(n_1656)
);

AO32x2_ASAP7_75t_L g1657 ( 
.A1(n_1545),
.A2(n_1576),
.A3(n_1603),
.B1(n_1629),
.B2(n_1547),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1583),
.B(n_1542),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1578),
.B(n_1534),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1539),
.B(n_1559),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1555),
.A2(n_1556),
.B(n_1615),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1534),
.B(n_1585),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1563),
.B(n_1607),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1560),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1563),
.B(n_1607),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1625),
.A2(n_1608),
.B1(n_1627),
.B2(n_1584),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1565),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1549),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1551),
.B(n_1553),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1613),
.A2(n_1555),
.B(n_1552),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1561),
.B(n_1554),
.Y(n_1671)
);

AO32x2_ASAP7_75t_L g1672 ( 
.A1(n_1545),
.A2(n_1576),
.A3(n_1603),
.B1(n_1629),
.B2(n_1547),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1564),
.B(n_1577),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1535),
.B(n_1566),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_SL g1675 ( 
.A(n_1565),
.B(n_1567),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1579),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1562),
.Y(n_1677)
);

BUFx2_ASAP7_75t_R g1678 ( 
.A(n_1541),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1627),
.B(n_1596),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1551),
.B(n_1553),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1624),
.A2(n_1633),
.B1(n_1631),
.B2(n_1630),
.C(n_1619),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1588),
.B(n_1616),
.Y(n_1682)
);

AO21x2_ASAP7_75t_L g1683 ( 
.A1(n_1612),
.A2(n_1618),
.B(n_1620),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1613),
.A2(n_1624),
.B(n_1614),
.C(n_1631),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_L g1685 ( 
.A(n_1595),
.B(n_1541),
.Y(n_1685)
);

NOR4xp25_ASAP7_75t_SL g1686 ( 
.A(n_1595),
.B(n_1589),
.C(n_1590),
.D(n_1538),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1687)
);

AO21x1_ASAP7_75t_L g1688 ( 
.A1(n_1622),
.A2(n_1611),
.B(n_1586),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1586),
.A2(n_1622),
.B(n_1611),
.C(n_1638),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1637),
.Y(n_1690)
);

AOI211xp5_ASAP7_75t_L g1691 ( 
.A1(n_1556),
.A2(n_1587),
.B(n_1615),
.C(n_1638),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1602),
.A2(n_1598),
.B(n_1592),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1568),
.B(n_1569),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1592),
.A2(n_1638),
.B(n_1552),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1549),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1634),
.A2(n_1597),
.B1(n_1632),
.B2(n_1591),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1633),
.A2(n_1630),
.B1(n_1591),
.B2(n_1580),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1597),
.A2(n_1591),
.B1(n_1639),
.B2(n_1641),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1633),
.A2(n_1610),
.B(n_1600),
.C(n_1630),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_SL g1700 ( 
.A1(n_1579),
.A2(n_1641),
.B(n_1639),
.C(n_1636),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1597),
.Y(n_1701)
);

CKINVDCx11_ASAP7_75t_R g1702 ( 
.A(n_1640),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1594),
.B(n_1575),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1581),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1597),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1537),
.B(n_1574),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1591),
.A2(n_1626),
.B(n_1546),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1602),
.A2(n_1598),
.B(n_1581),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1667),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1708),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1655),
.B(n_1580),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1668),
.B(n_1695),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1658),
.B(n_1580),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1661),
.B(n_1617),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1653),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1708),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1668),
.B(n_1544),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1654),
.A2(n_1635),
.B1(n_1617),
.B2(n_1600),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1642),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1671),
.B(n_1651),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1646),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1695),
.B(n_1671),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1708),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1692),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1664),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1670),
.B(n_1544),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1666),
.A2(n_1681),
.B1(n_1697),
.B2(n_1688),
.Y(n_1727)
);

INVx5_ASAP7_75t_L g1728 ( 
.A(n_1706),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1670),
.B(n_1543),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1704),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1653),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1704),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1677),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1663),
.B(n_1617),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1681),
.A2(n_1590),
.B1(n_1600),
.B2(n_1536),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1665),
.B(n_1662),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1694),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1687),
.B(n_1593),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1659),
.B(n_1593),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1673),
.B(n_1606),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1691),
.B(n_1601),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1657),
.B(n_1582),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1728),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1715),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1730),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1717),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1674),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1722),
.B(n_1690),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1728),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1734),
.B(n_1736),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1712),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1712),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1650),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1728),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1730),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1716),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1727),
.B(n_1647),
.C(n_1697),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1727),
.A2(n_1683),
.B1(n_1656),
.B2(n_1643),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1710),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1737),
.B(n_1699),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1719),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1736),
.B(n_1657),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1736),
.B(n_1657),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1735),
.A2(n_1644),
.B1(n_1656),
.B2(n_1683),
.Y(n_1768)
);

OAI33xp33_ASAP7_75t_L g1769 ( 
.A1(n_1726),
.A2(n_1696),
.A3(n_1660),
.B1(n_1698),
.B2(n_1703),
.B3(n_1693),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1713),
.B(n_1699),
.Y(n_1770)
);

NAND4xp25_ASAP7_75t_L g1771 ( 
.A(n_1735),
.B(n_1647),
.C(n_1652),
.D(n_1648),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1718),
.A2(n_1652),
.B1(n_1684),
.B2(n_1689),
.C(n_1679),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1721),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1716),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1711),
.B(n_1657),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1713),
.B(n_1679),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1737),
.A2(n_1685),
.B(n_1702),
.C(n_1640),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1725),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1711),
.B(n_1672),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1718),
.A2(n_1572),
.B1(n_1707),
.B2(n_1609),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1672),
.Y(n_1782)
);

OAI31xp33_ASAP7_75t_L g1783 ( 
.A1(n_1720),
.A2(n_1684),
.A3(n_1689),
.B(n_1741),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1709),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1728),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1739),
.B(n_1672),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1732),
.B(n_1726),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1725),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1763),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1765),
.B(n_1742),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1763),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1771),
.B(n_1720),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1767),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1744),
.B(n_1732),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1765),
.B(n_1742),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1767),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1773),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1771),
.B(n_1676),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1773),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1774),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1766),
.B(n_1742),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1758),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1758),
.Y(n_1804)
);

INVx4_ASAP7_75t_L g1805 ( 
.A(n_1743),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1758),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1756),
.A2(n_1723),
.B(n_1724),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1744),
.B(n_1725),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1766),
.B(n_1709),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1784),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1752),
.B(n_1728),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1743),
.B(n_1728),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1752),
.B(n_1738),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1747),
.B(n_1733),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1764),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1764),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1784),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1764),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1782),
.B(n_1738),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1782),
.B(n_1738),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1779),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1779),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1676),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1747),
.B(n_1733),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1789),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1792),
.B(n_1753),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1792),
.B(n_1753),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1813),
.B(n_1824),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1803),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1799),
.A2(n_1759),
.B(n_1762),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1791),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1813),
.B(n_1745),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1803),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_L g1837 ( 
.A(n_1799),
.B(n_1778),
.C(n_1759),
.D(n_1783),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1812),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1791),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1794),
.Y(n_1840)
);

INVxp67_ASAP7_75t_L g1841 ( 
.A(n_1825),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1805),
.B(n_1743),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1803),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1794),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1813),
.B(n_1745),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1797),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1817),
.B(n_1776),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1797),
.Y(n_1850)
);

NAND4xp25_ASAP7_75t_L g1851 ( 
.A(n_1825),
.B(n_1783),
.C(n_1750),
.D(n_1762),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1795),
.B(n_1787),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1776),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1798),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1798),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1745),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1795),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1815),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1800),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1800),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1815),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1809),
.B(n_1780),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1809),
.B(n_1780),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1801),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1808),
.B(n_1787),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1801),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1805),
.B(n_1756),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1793),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1824),
.B(n_1786),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1812),
.B(n_1805),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1815),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1827),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1828),
.B(n_1808),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1833),
.B(n_1809),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1827),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1842),
.B(n_1812),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1829),
.B(n_1814),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1857),
.B(n_1819),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1841),
.Y(n_1880)
);

NAND2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_SL g1882 ( 
.A(n_1837),
.B(n_1678),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1830),
.B(n_1790),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1830),
.B(n_1790),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1838),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_1814),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1852),
.B(n_1826),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1835),
.B(n_1796),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1831),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1847),
.B(n_1796),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1845),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1834),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1851),
.B(n_1819),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1847),
.B(n_1796),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1834),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1839),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1870),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1856),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1865),
.B(n_1820),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1838),
.B(n_1649),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1856),
.B(n_1802),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1869),
.B(n_1838),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1849),
.A2(n_1769),
.B1(n_1772),
.B2(n_1760),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1865),
.B(n_1826),
.Y(n_1906)
);

OAI211xp5_ASAP7_75t_L g1907 ( 
.A1(n_1868),
.A2(n_1805),
.B(n_1853),
.C(n_1863),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1862),
.B(n_1748),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1882),
.B(n_1874),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1880),
.B(n_1869),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1905),
.A2(n_1769),
.B1(n_1768),
.B2(n_1772),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1886),
.B(n_1820),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1872),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1895),
.A2(n_1770),
.B1(n_1802),
.B2(n_1811),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1893),
.A2(n_1770),
.B(n_1859),
.C(n_1866),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1902),
.A2(n_1768),
.B1(n_1781),
.B2(n_1714),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1872),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1878),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1885),
.A2(n_1713),
.B1(n_1710),
.B2(n_1729),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1878),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1907),
.A2(n_1839),
.B(n_1840),
.C(n_1866),
.Y(n_1921)
);

NOR3xp33_ASAP7_75t_L g1922 ( 
.A(n_1875),
.B(n_1850),
.C(n_1840),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1886),
.B(n_1820),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1891),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1900),
.B(n_1802),
.Y(n_1925)
);

OAI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1873),
.A2(n_1871),
.B1(n_1832),
.B2(n_1861),
.C(n_1836),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1873),
.A2(n_1871),
.B1(n_1843),
.B2(n_1861),
.C(n_1836),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1900),
.B(n_1702),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1890),
.B(n_1842),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1877),
.B(n_1685),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1876),
.A2(n_1700),
.B(n_1867),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1890),
.B(n_1846),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1894),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1892),
.B(n_1867),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1892),
.B(n_1848),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1913),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1934),
.B(n_1896),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1929),
.B(n_1896),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1917),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1909),
.A2(n_1899),
.B(n_1887),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1918),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1920),
.Y(n_1942)
);

INVxp33_ASAP7_75t_L g1943 ( 
.A(n_1909),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1910),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1911),
.A2(n_1877),
.B1(n_1879),
.B2(n_1901),
.C(n_1908),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1915),
.B(n_1903),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1925),
.B(n_1908),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1912),
.B(n_1903),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_SL g1949 ( 
.A(n_1928),
.B(n_1589),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1924),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1923),
.B(n_1883),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1933),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1932),
.Y(n_1953)
);

NAND5xp2_ASAP7_75t_SL g1954 ( 
.A(n_1931),
.B(n_1904),
.C(n_1884),
.D(n_1883),
.E(n_1881),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1921),
.A2(n_1887),
.B(n_1904),
.C(n_1898),
.Y(n_1955)
);

AOI211xp5_ASAP7_75t_L g1956 ( 
.A1(n_1914),
.A2(n_1897),
.B(n_1700),
.C(n_1884),
.Y(n_1956)
);

OR3x1_ASAP7_75t_L g1957 ( 
.A(n_1944),
.B(n_1930),
.C(n_1881),
.Y(n_1957)
);

AOI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1943),
.A2(n_1926),
.B(n_1927),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1943),
.B(n_1949),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1947),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1938),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1947),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1951),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1951),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1948),
.Y(n_1965)
);

AOI21xp33_ASAP7_75t_L g1966 ( 
.A1(n_1950),
.A2(n_1952),
.B(n_1953),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1936),
.Y(n_1967)
);

A2O1A1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1945),
.A2(n_1916),
.B(n_1946),
.C(n_1956),
.Y(n_1968)
);

OAI211xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1968),
.A2(n_1940),
.B(n_1955),
.C(n_1954),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1961),
.B(n_1938),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1957),
.A2(n_1930),
.B1(n_1953),
.B2(n_1935),
.Y(n_1971)
);

NOR4xp25_ASAP7_75t_L g1972 ( 
.A(n_1966),
.B(n_1942),
.C(n_1941),
.D(n_1939),
.Y(n_1972)
);

AOI322xp5_ASAP7_75t_L g1973 ( 
.A1(n_1958),
.A2(n_1919),
.A3(n_1922),
.B1(n_1937),
.B2(n_1843),
.C1(n_1832),
.C2(n_1858),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1958),
.A2(n_1919),
.B1(n_1922),
.B2(n_1937),
.C(n_1858),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1961),
.B(n_1960),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1959),
.A2(n_1881),
.B(n_1888),
.Y(n_1976)
);

NAND4xp25_ASAP7_75t_L g1977 ( 
.A(n_1963),
.B(n_1889),
.C(n_1888),
.D(n_1867),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1964),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1962),
.Y(n_1979)
);

AND3x1_ASAP7_75t_L g1980 ( 
.A(n_1972),
.B(n_1965),
.C(n_1967),
.Y(n_1980)
);

OAI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1974),
.A2(n_1969),
.B1(n_1973),
.B2(n_1979),
.C(n_1975),
.Y(n_1981)
);

NAND4xp25_ASAP7_75t_SL g1982 ( 
.A(n_1970),
.B(n_1889),
.C(n_1906),
.D(n_1680),
.Y(n_1982)
);

AOI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1971),
.A2(n_1906),
.B1(n_1864),
.B2(n_1860),
.C(n_1859),
.Y(n_1983)
);

AOI22x1_ASAP7_75t_L g1984 ( 
.A1(n_1979),
.A2(n_1793),
.B1(n_1860),
.B2(n_1855),
.Y(n_1984)
);

AOI221xp5_ASAP7_75t_L g1985 ( 
.A1(n_1978),
.A2(n_1864),
.B1(n_1855),
.B2(n_1850),
.C(n_1761),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1977),
.A2(n_1761),
.B1(n_1854),
.B2(n_1710),
.C(n_1806),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1980),
.A2(n_1976),
.B1(n_1645),
.B2(n_1804),
.Y(n_1987)
);

AO22x1_ASAP7_75t_L g1988 ( 
.A1(n_1981),
.A2(n_1793),
.B1(n_1669),
.B2(n_1812),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1983),
.A2(n_1793),
.B1(n_1812),
.B2(n_1750),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1986),
.Y(n_1990)
);

OAI211xp5_ASAP7_75t_L g1991 ( 
.A1(n_1984),
.A2(n_1793),
.B(n_1686),
.C(n_1731),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1985),
.A2(n_1823),
.B1(n_1822),
.B2(n_1821),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1982),
.A2(n_1807),
.B(n_1811),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1990),
.B(n_1746),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1988),
.B(n_1701),
.Y(n_1995)
);

NAND4xp75_ASAP7_75t_L g1996 ( 
.A(n_1987),
.B(n_1811),
.C(n_1751),
.D(n_1785),
.Y(n_1996)
);

NAND2x1p5_ASAP7_75t_L g1997 ( 
.A(n_1991),
.B(n_1701),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1993),
.A2(n_1710),
.B1(n_1806),
.B2(n_1804),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1989),
.B(n_1746),
.Y(n_1999)
);

OAI321xp33_ASAP7_75t_L g2000 ( 
.A1(n_1997),
.A2(n_1992),
.A3(n_1741),
.B1(n_1804),
.B2(n_1816),
.C(n_1806),
.Y(n_2000)
);

OAI321xp33_ASAP7_75t_L g2001 ( 
.A1(n_1994),
.A2(n_1741),
.A3(n_1804),
.B1(n_1806),
.B2(n_1816),
.C(n_1777),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_L g2002 ( 
.A(n_1995),
.B(n_1999),
.C(n_1998),
.Y(n_2002)
);

AOI211x1_ASAP7_75t_L g2003 ( 
.A1(n_1996),
.A2(n_1823),
.B(n_1822),
.C(n_1821),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_SL g2004 ( 
.A1(n_2002),
.A2(n_1731),
.B1(n_1715),
.B2(n_1705),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_2004),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2005),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_2005),
.B(n_2003),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_2007),
.B(n_2000),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_2007),
.Y(n_2009)
);

OAI21xp33_ASAP7_75t_L g2010 ( 
.A1(n_2009),
.A2(n_2006),
.B(n_2001),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_2008),
.A2(n_1816),
.B1(n_1818),
.B2(n_1775),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2010),
.Y(n_2012)
);

OR2x6_ASAP7_75t_L g2013 ( 
.A(n_2012),
.B(n_1705),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2013),
.Y(n_2014)
);

OAI221xp5_ASAP7_75t_R g2015 ( 
.A1(n_2014),
.A2(n_2011),
.B1(n_1757),
.B2(n_1675),
.C(n_1715),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_2015),
.A2(n_1755),
.B1(n_1816),
.B2(n_1749),
.Y(n_2016)
);


endmodule