module real_jpeg_6756_n_31 (n_17, n_8, n_0, n_21, n_2, n_29, n_10, n_175, n_9, n_178, n_12, n_24, n_170, n_176, n_6, n_28, n_171, n_169, n_177, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_30, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_29;
input n_10;
input n_175;
input n_9;
input n_178;
input n_12;
input n_24;
input n_170;
input n_176;
input n_6;
input n_28;
input n_171;
input n_169;
input n_177;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_30;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_0),
.Y(n_95)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_3),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_155),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_6),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_8),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_113),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_9),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_10),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_13),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_13),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_14),
.B(n_98),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_69),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_17),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_18),
.B(n_44),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_18),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_19),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_21),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_23),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_54),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_24),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_25),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_26),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_27),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_27),
.B(n_66),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_29),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_162),
.Y(n_31)
);

AO21x1_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_42),
.B(n_161),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_34),
.B(n_41),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_36),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_36),
.B(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_38),
.B(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_39),
.B(n_139),
.Y(n_138)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_40),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_41),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B(n_160),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_150),
.B(n_157),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_130),
.B(n_144),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_71),
.B(n_118),
.C(n_127),
.Y(n_51)
);

NOR4xp25_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.C(n_65),
.D(n_68),
.Y(n_52)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_91),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_112),
.B(n_117),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_105),
.B(n_111),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_82),
.B1(n_102),
.B2(n_103),
.C(n_104),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_99),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B(n_101),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_97),
.B(n_100),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_110),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.C(n_125),
.D(n_126),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.C(n_140),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_140),
.B(n_145),
.C(n_148),
.D(n_149),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_169),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_170),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_171),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_172),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_173),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_174),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_175),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_176),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_177),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_178),
.Y(n_114)
);


endmodule