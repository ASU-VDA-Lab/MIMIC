module fake_jpeg_17539_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_10),
.B1(n_16),
.B2(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_15),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_22),
.B(n_14),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_36),
.C(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_29),
.B1(n_2),
.B2(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_39),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.C(n_42),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.C(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_50),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_42),
.B(n_32),
.C(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_4),
.Y(n_59)
);


endmodule