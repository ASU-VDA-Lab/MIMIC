module real_jpeg_20609_n_17 (n_8, n_0, n_2, n_348, n_10, n_9, n_12, n_6, n_347, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_348;
input n_10;
input n_9;
input n_12;
input n_6;
input n_347;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_0),
.A2(n_52),
.B1(n_53),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_0),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_0),
.A2(n_70),
.B1(n_71),
.B2(n_106),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_106),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_106),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_1),
.A2(n_70),
.B1(n_71),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_1),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_162),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_162),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_162),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_35),
.B1(n_52),
.B2(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_3),
.A2(n_35),
.B1(n_70),
.B2(n_71),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_23),
.B1(n_70),
.B2(n_71),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_4),
.A2(n_23),
.B1(n_52),
.B2(n_53),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_70),
.B1(n_71),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_111),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_111),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_111),
.Y(n_251)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_7),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_134),
.B(n_160),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_9),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_70),
.B1(n_71),
.B2(n_94),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_94),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_63),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_53),
.B(n_66),
.C(n_91),
.D(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_12),
.B(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_12),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_12),
.A2(n_112),
.B(n_114),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_32),
.B(n_48),
.C(n_150),
.D(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_12),
.B(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_36),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_31),
.B(n_33),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_131),
.Y(n_209)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_21),
.B(n_42),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_22),
.A2(n_26),
.B1(n_36),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_24),
.A2(n_28),
.B(n_131),
.C(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_26),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_26),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_27),
.A2(n_30),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_27),
.A2(n_30),
.B1(n_220),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_27),
.A2(n_211),
.B(n_251),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_27),
.A2(n_30),
.B1(n_60),
.B2(n_295),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_30),
.A2(n_221),
.B(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_36),
.B(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_80),
.B(n_345),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_75),
.C(n_77),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_43),
.A2(n_44),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_45),
.A2(n_46),
.B1(n_64),
.B2(n_320),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_47),
.A2(n_56),
.B1(n_171),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_206),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_51),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_48),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_48),
.A2(n_51),
.B1(n_248),
.B2(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_48),
.A2(n_51),
.B1(n_267),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_50),
.Y(n_158)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_52),
.B(n_54),
.Y(n_157)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_53),
.A2(n_150),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_56),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_56),
.A2(n_172),
.B(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_58),
.A2(n_59),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_64),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_73),
.B1(n_105),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_65),
.A2(n_148),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_65),
.A2(n_73),
.B1(n_203),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_65),
.A2(n_73),
.B1(n_233),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_65),
.A2(n_73),
.B1(n_242),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_66),
.A2(n_69),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_70),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_71),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_73),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_73),
.A2(n_107),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_74),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_75),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_338),
.B(n_344),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_311),
.A3(n_331),
.B1(n_336),
.B2(n_337),
.C(n_347),
.Y(n_81)
);

AOI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_259),
.A3(n_299),
.B1(n_305),
.B2(n_310),
.C(n_348),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_214),
.C(n_255),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_186),
.B(n_213),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_165),
.B(n_185),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_142),
.B(n_164),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_117),
.B(n_141),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_89),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_104),
.C(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_114),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_125),
.B1(n_161),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_112),
.A2(n_113),
.B1(n_176),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_112),
.A2(n_196),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_112),
.A2(n_125),
.B1(n_231),
.B2(n_240),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_112),
.A2(n_125),
.B(n_240),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_121),
.B(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_113),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_128),
.B(n_140),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_131),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_135),
.B(n_139),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_132),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_155),
.B2(n_163),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_154),
.C(n_163),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_167),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_181),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_182),
.C(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_180),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_177),
.C(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_200),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_199),
.C(n_200),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_195),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_215),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_235),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_235),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.C(n_234),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_234),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_232),
.Y(n_244)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_253),
.B2(n_254),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_238),
.B(n_243),
.C(n_254),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_241),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_249),
.C(n_252),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_277),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_260),
.B(n_277),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_270),
.C(n_276),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_261),
.A2(n_262),
.B1(n_270),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_275),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_272),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_271),
.A2(n_290),
.B(n_294),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_273),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_297),
.B2(n_298),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_288),
.B2(n_289),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_289),
.C(n_298),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_285),
.B(n_287),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_285),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_286),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_287),
.A2(n_313),
.B1(n_322),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_324),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.C(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_314),
.A2(n_315),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_320),
.C(n_321),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_326),
.C(n_330),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_318),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_343),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_340),
.Y(n_342)
);


endmodule