module fake_jpeg_13979_n_519 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_26),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_50),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_54),
.Y(n_148)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_63),
.B(n_89),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_15),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_19),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_87),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_92),
.Y(n_154)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_14),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_97),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_102),
.A2(n_111),
.B1(n_144),
.B2(n_121),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_30),
.B(n_21),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_141),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_83),
.B1(n_51),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_114),
.A2(n_133),
.B1(n_17),
.B2(n_48),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_39),
.C(n_46),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_45),
.C(n_22),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_34),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_142),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_62),
.A2(n_21),
.B1(n_41),
.B2(n_30),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_77),
.B(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_38),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_36),
.B1(n_29),
.B2(n_48),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_34),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_156),
.Y(n_166)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_50),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_R g162 ( 
.A(n_134),
.B(n_60),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_69),
.B1(n_68),
.B2(n_66),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_164),
.A2(n_179),
.B1(n_186),
.B2(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_176),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_114),
.A2(n_74),
.B1(n_73),
.B2(n_41),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_168),
.A2(n_180),
.B1(n_196),
.B2(n_22),
.Y(n_242)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_39),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_175),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_101),
.B(n_36),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_38),
.B1(n_46),
.B2(n_18),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_18),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_185),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_48),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_36),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_110),
.A2(n_17),
.B1(n_45),
.B2(n_32),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_95),
.B1(n_93),
.B2(n_36),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_195),
.A3(n_121),
.B1(n_124),
.B2(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_17),
.B1(n_45),
.B2(n_27),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_33),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_201),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_136),
.B(n_25),
.C(n_23),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_149),
.A2(n_25),
.B1(n_23),
.B2(n_44),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_102),
.A2(n_59),
.B(n_56),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_128),
.B(n_44),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_44),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_206),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_212),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_109),
.B(n_205),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_150),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_243),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_161),
.B(n_108),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_195),
.B1(n_204),
.B2(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_150),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_123),
.A3(n_104),
.B1(n_115),
.B2(n_108),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_168),
.Y(n_249)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_184),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_246),
.B(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_251),
.B1(n_258),
.B2(n_263),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_229),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_235),
.B1(n_238),
.B2(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_254),
.B1(n_244),
.B2(n_229),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_161),
.B1(n_200),
.B2(n_201),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_158),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_253),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_158),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_158),
.B1(n_180),
.B2(n_196),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_203),
.B1(n_121),
.B2(n_172),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_255),
.A2(n_261),
.B1(n_193),
.B2(n_192),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_183),
.CI(n_182),
.CON(n_256),
.SN(n_256)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_217),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_159),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_257),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_111),
.B1(n_177),
.B2(n_122),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_211),
.A2(n_112),
.B1(n_124),
.B2(n_106),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_264),
.B(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_212),
.A2(n_122),
.B1(n_104),
.B2(n_115),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_197),
.B(n_170),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_218),
.A2(n_159),
.B(n_160),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_222),
.A2(n_243),
.B1(n_226),
.B2(n_216),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_270),
.B1(n_213),
.B2(n_230),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_187),
.C(n_198),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_279),
.C(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_151),
.B1(n_118),
.B2(n_100),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_169),
.B(n_22),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_275),
.B(n_277),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_112),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_216),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_237),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_228),
.B(n_171),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_190),
.C(n_181),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_252),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_301),
.C(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_289),
.B1(n_298),
.B2(n_305),
.Y(n_323)
);

NAND2x1_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_219),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_312),
.B(n_275),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_279),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_293),
.B(n_247),
.CI(n_256),
.CON(n_319),
.SN(n_319)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_306),
.Y(n_339)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_249),
.A2(n_217),
.B1(n_241),
.B2(n_165),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_304),
.B1(n_309),
.B2(n_275),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_265),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_300),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_163),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_248),
.A2(n_210),
.B1(n_240),
.B2(n_213),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_254),
.A2(n_118),
.B1(n_119),
.B2(n_148),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_209),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_209),
.Y(n_308)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_260),
.A2(n_234),
.B(n_208),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_258),
.B1(n_271),
.B2(n_260),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_317),
.A2(n_318),
.B(n_336),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_298),
.A2(n_262),
.B1(n_250),
.B2(n_251),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_330),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_281),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_338),
.B1(n_302),
.B2(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_268),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_343),
.Y(n_372)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_264),
.B(n_257),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_345),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_281),
.A2(n_256),
.B1(n_279),
.B2(n_268),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_288),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_341),
.B(n_282),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_291),
.B(n_266),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_344),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_257),
.C(n_270),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_286),
.A2(n_257),
.B1(n_263),
.B2(n_272),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_346),
.A2(n_347),
.B1(n_280),
.B2(n_210),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_286),
.A2(n_272),
.B1(n_274),
.B2(n_240),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_234),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_293),
.B1(n_299),
.B2(n_304),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_362),
.B1(n_365),
.B2(n_370),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_336),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_327),
.B(n_308),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_376),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_317),
.A2(n_282),
.B(n_302),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_377),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_305),
.B1(n_290),
.B2(n_312),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_323),
.A2(n_311),
.B1(n_280),
.B2(n_313),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_373),
.B1(n_324),
.B2(n_340),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_323),
.A2(n_301),
.B1(n_210),
.B2(n_174),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_338),
.A2(n_230),
.B1(n_234),
.B2(n_148),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_369),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_339),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_237),
.B1(n_188),
.B2(n_208),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_220),
.B1(n_214),
.B2(n_231),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_220),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_192),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_326),
.C(n_334),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_384),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_387),
.A2(n_408),
.B1(n_410),
.B2(n_397),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_380),
.B(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_376),
.B(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_325),
.Y(n_393)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_352),
.A2(n_357),
.B(n_366),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_316),
.C(n_345),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_404),
.C(n_405),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_339),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_319),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_322),
.Y(n_401)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_359),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_403),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_355),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_335),
.C(n_331),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_328),
.C(n_315),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_329),
.C(n_333),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_409),
.C(n_373),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_354),
.B(n_358),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_361),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_382),
.A2(n_357),
.B1(n_368),
.B2(n_378),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_415),
.B1(n_392),
.B2(n_409),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_382),
.A2(n_368),
.B1(n_375),
.B2(n_354),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_429),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_381),
.C(n_375),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_423),
.C(n_427),
.Y(n_439)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_367),
.C(n_363),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_424),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_367),
.B(n_363),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_426),
.A2(n_402),
.B(n_27),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_358),
.C(n_329),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_371),
.B(n_214),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_R g430 ( 
.A1(n_406),
.A2(n_389),
.B1(n_387),
.B2(n_400),
.Y(n_430)
);

OAI21xp33_ASAP7_75t_SL g443 ( 
.A1(n_430),
.A2(n_383),
.B(n_399),
.Y(n_443)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_193),
.B1(n_13),
.B2(n_12),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_432),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_231),
.B(n_191),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_405),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_445),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_407),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_441),
.B(n_452),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_442),
.A2(n_429),
.B1(n_428),
.B2(n_436),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_413),
.B1(n_422),
.B2(n_423),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_403),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_448),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_414),
.A2(n_146),
.B1(n_24),
.B2(n_12),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_453),
.B1(n_455),
.B2(n_431),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_24),
.C(n_146),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_451),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_193),
.C(n_1),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_419),
.B(n_193),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_433),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_435),
.B(n_10),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_412),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_415),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_434),
.Y(n_461)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_450),
.C(n_413),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_464),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_472),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_10),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_427),
.C(n_418),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_469),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_438),
.A2(n_421),
.B1(n_424),
.B2(n_416),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_467),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_468),
.A2(n_451),
.B1(n_455),
.B2(n_454),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_425),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_425),
.C(n_426),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_471),
.C(n_473),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_0),
.C(n_1),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_440),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_0),
.C(n_1),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_9),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_3),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_467),
.A2(n_447),
.B(n_448),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_475),
.A2(n_459),
.B(n_473),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_466),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_479),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_446),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_478),
.A2(n_6),
.B(n_7),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_453),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_480),
.B(n_484),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_483),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_2),
.Y(n_484)
);

AOI21x1_ASAP7_75t_SL g485 ( 
.A1(n_457),
.A2(n_3),
.B(n_4),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_485),
.A2(n_5),
.B(n_6),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_4),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_490),
.B(n_493),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_498),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_488),
.B(n_460),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_460),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_482),
.B(n_475),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_471),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_495),
.B(n_497),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_6),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_486),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_499),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_508),
.B(n_509),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_481),
.B(n_478),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_494),
.A2(n_476),
.B(n_479),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_496),
.C(n_491),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_513),
.C(n_502),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_490),
.C(n_485),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_6),
.C(n_8),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_510),
.C(n_506),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_516),
.A2(n_514),
.B(n_6),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_8),
.C(n_321),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_8),
.Y(n_519)
);


endmodule