module real_jpeg_16982_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_419),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_0),
.B(n_420),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_23),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

AND2x4_ASAP7_75t_SL g145 ( 
.A(n_1),
.B(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_2),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_3),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_3),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_4),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_4),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_4),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_4),
.B(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_5),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_6),
.B(n_38),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_6),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_7),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_8),
.B(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_9),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_11),
.Y(n_420)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g274 ( 
.A(n_12),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g268 ( 
.A(n_13),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_100),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_60),
.B(n_99),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_60),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_48),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.C(n_39),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_19),
.A2(n_20),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_21),
.A2(n_32),
.B1(n_41),
.B2(n_92),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_41),
.B1(n_47),
.B2(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_22),
.A2(n_47),
.B1(n_127),
.B2(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_22),
.B(n_112),
.C(n_227),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_22),
.A2(n_91),
.B(n_96),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_22),
.A2(n_47),
.B1(n_227),
.B2(n_231),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_25),
.A2(n_26),
.B1(n_236),
.B2(n_238),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_29),
.C(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_29),
.A2(n_33),
.B1(n_53),
.B2(n_57),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_29),
.B(n_112),
.C(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_29),
.B(n_286),
.C(n_287),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_29),
.B(n_266),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_29),
.A2(n_33),
.B1(n_287),
.B2(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_29),
.A2(n_33),
.B1(n_66),
.B2(n_237),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_29),
.B(n_66),
.C(n_345),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_33),
.B(n_266),
.C(n_290),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_47),
.Y(n_40)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_41),
.A2(n_142),
.B(n_171),
.C(n_177),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_41),
.B(n_142),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_41),
.A2(n_92),
.B1(n_142),
.B2(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_41),
.B(n_93),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_41),
.B(n_66),
.C(n_94),
.Y(n_257)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_98),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_46),
.B(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_46),
.A2(n_145),
.B(n_172),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_47),
.B(n_122),
.C(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_53),
.A2(n_57),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_53),
.B(n_147),
.C(n_198),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_53),
.A2(n_57),
.B1(n_144),
.B2(n_149),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_53),
.A2(n_57),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_53),
.B(n_132),
.C(n_145),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_57),
.B(n_112),
.C(n_334),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_84),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_61),
.B(n_64),
.Y(n_410)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.C(n_79),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_69),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_66),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_66),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_66),
.A2(n_237),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_67),
.A2(n_93),
.B1(n_94),
.B2(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_67),
.A2(n_94),
.B(n_123),
.C(n_177),
.Y(n_222)
);

AO22x1_ASAP7_75t_L g317 ( 
.A1(n_67),
.A2(n_207),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_67),
.B(n_153),
.C(n_318),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_207),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_79),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_75),
.A2(n_240),
.B(n_246),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_75),
.B(n_240),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_75),
.A2(n_89),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_75),
.B(n_93),
.C(n_133),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_128),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_76),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_78),
.Y(n_201)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_84),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_97),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_85),
.A2(n_86),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_90),
.B(n_97),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_96),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_93),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_184),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_93),
.A2(n_94),
.B1(n_132),
.B2(n_133),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_373),
.B(n_411),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_280),
.A3(n_360),
.B1(n_366),
.B2(n_371),
.C(n_372),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_250),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_216),
.B(n_249),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_192),
.B(n_215),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_168),
.B(n_191),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_150),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_150),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_129),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_120),
.B2(n_121),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_121),
.C(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_112),
.A2(n_119),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_117),
.A2(n_212),
.B1(n_226),
.B2(n_232),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_119),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_123),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_122),
.A2(n_123),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_127),
.A2(n_153),
.B1(n_198),
.B2(n_202),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_127),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_183),
.B(n_185),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_131),
.A2(n_142),
.B(n_149),
.Y(n_203)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_132),
.A2(n_133),
.B1(n_160),
.B2(n_161),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_145),
.B(n_147),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_145),
.Y(n_147)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_156),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_145),
.B(n_172),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_145),
.A2(n_166),
.B1(n_172),
.B2(n_175),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_164),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_153),
.B(n_202),
.C(n_257),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_164),
.B1(n_165),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_156),
.B(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_160),
.A2(n_161),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_161),
.B(n_267),
.C(n_271),
.Y(n_286)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_181),
.B(n_190),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_178),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_175),
.B1(n_227),
.B2(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_212),
.C(n_227),
.Y(n_277)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_187),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B(n_189),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_194),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_204),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_203),
.C(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_210),
.C(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_248),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_220),
.C(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_225),
.C(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_224),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_247),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_239),
.C(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_251),
.B(n_252),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_253),
.B(n_264),
.C(n_279),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_356)
);

XNOR2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_279),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_277),
.C(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_348),
.Y(n_280)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_323),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_282),
.B(n_323),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_303),
.C(n_311),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_311),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_296),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_289),
.B1(n_294),
.B2(n_295),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_295),
.C(n_296),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_301),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

XOR2x2_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_314),
.C(n_316),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_341),
.C(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_341),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_327),
.B(n_331),
.C(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_340),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_344),
.C(n_347),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

AOI31xp67_ASAP7_75t_SL g366 ( 
.A1(n_348),
.A2(n_361),
.A3(n_367),
.B(n_370),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_351),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_356),
.C(n_357),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_352),
.A2(n_353),
.B1(n_357),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_365),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_395),
.C(n_406),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_378),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_381),
.C(n_388),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_386),
.C(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_390),
.B(n_393),
.C(n_394),
.Y(n_404)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_396),
.A2(n_414),
.B(n_415),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_405),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_405),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_404),
.C(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_406),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NAND2x1_ASAP7_75t_SL g418 ( 
.A(n_407),
.B(n_409),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_416),
.B(n_417),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

CKINVDCx11_ASAP7_75t_R g417 ( 
.A(n_418),
.Y(n_417)
);


endmodule