module fake_netlist_5_1557_n_473 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_473);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_473;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_124;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_127;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_155;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_373;
wire n_147;
wire n_307;
wire n_439;
wire n_150;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_430;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_213;
wire n_129;
wire n_342;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_461;
wire n_333;
wire n_309;
wire n_462;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_463;
wire n_239;
wire n_466;
wire n_420;
wire n_310;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_441;
wire n_450;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_269;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_121;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_22),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_23),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_25),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_2),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_38),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_60),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g148 ( 
.A(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_35),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_30),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_24),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_56),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_49),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_36),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_71),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_17),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_77),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_41),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_66),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_82),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_93),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_78),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_45),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_21),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_18),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_74),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_6),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_42),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_15),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_0),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_10),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_2),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_139),
.B(n_3),
.C(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_135),
.B(n_3),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_149),
.B(n_157),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_165),
.B(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_143),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_224),
.B(n_150),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_215),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_161),
.Y(n_244)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_144),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_148),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_189),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_186),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_166),
.B1(n_146),
.B2(n_170),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_5),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_203),
.A2(n_169),
.B1(n_198),
.B2(n_154),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_231),
.B(n_154),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_120),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_229),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_241),
.B(n_267),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_205),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_199),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_180),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_254),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_200),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_238),
.A2(n_216),
.B1(n_180),
.B2(n_193),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_234),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_201),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_205),
.Y(n_309)
);

NAND2x2_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_253),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_245),
.A2(n_206),
.B1(n_201),
.B2(n_147),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

OR2x6_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_206),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_256),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_212),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

NAND2x1p5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_193),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_245),
.B1(n_258),
.B2(n_192),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_281),
.A2(n_173),
.B1(n_132),
.B2(n_142),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_186),
.B1(n_237),
.B2(n_152),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_176),
.B1(n_145),
.B2(n_155),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_196),
.B1(n_156),
.B2(n_158),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_256),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_121),
.B(n_162),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_240),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_316),
.A2(n_178),
.B1(n_171),
.B2(n_163),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_298),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_240),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_283),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_283),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_164),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_309),
.A2(n_183),
.B(n_167),
.C(n_168),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_294),
.A2(n_194),
.B1(n_179),
.B2(n_182),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_266),
.B(n_230),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_212),
.Y(n_358)
);

AO31x2_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_319),
.A3(n_185),
.B(n_188),
.Y(n_359)
);

AOI21xp33_ASAP7_75t_L g360 ( 
.A1(n_319),
.A2(n_159),
.B(n_172),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_284),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_344),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_296),
.B1(n_291),
.B2(n_310),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_333),
.A2(n_330),
.B1(n_323),
.B2(n_336),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_286),
.B1(n_296),
.B2(n_317),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_313),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_330),
.A2(n_291),
.B1(n_315),
.B2(n_312),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_302),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_286),
.B1(n_312),
.B2(n_302),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

OR2x6_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_288),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_286),
.B1(n_177),
.B2(n_174),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_341),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_295),
.B1(n_289),
.B2(n_292),
.Y(n_376)
);

CKINVDCx11_ASAP7_75t_R g377 ( 
.A(n_340),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_335),
.A2(n_349),
.B1(n_325),
.B2(n_332),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_292),
.B1(n_285),
.B2(n_293),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_293),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_325),
.A2(n_293),
.B1(n_227),
.B2(n_230),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_338),
.B(n_346),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_293),
.Y(n_386)
);

AOI222xp33_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_351),
.B1(n_327),
.B2(n_334),
.C1(n_322),
.C2(n_357),
.Y(n_387)
);

AOI222xp33_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_227),
.B1(n_7),
.B2(n_9),
.C1(n_6),
.C2(n_228),
.Y(n_388)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_364),
.A2(n_348),
.B1(n_354),
.B2(n_350),
.Y(n_390)
);

AOI221xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_360),
.B1(n_353),
.B2(n_354),
.C(n_230),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_360),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_384),
.B1(n_378),
.B2(n_383),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_359),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_266),
.B(n_320),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_362),
.A2(n_361),
.B1(n_389),
.B2(n_371),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_389),
.A2(n_228),
.B1(n_222),
.B2(n_9),
.Y(n_401)
);

AO31x2_ASAP7_75t_L g402 ( 
.A1(n_385),
.A2(n_228),
.A3(n_222),
.B(n_13),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_368),
.A2(n_320),
.B1(n_12),
.B2(n_16),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_320),
.B1(n_20),
.B2(n_26),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_381),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_390),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_376),
.B1(n_382),
.B2(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_407),
.A2(n_365),
.B1(n_377),
.B2(n_373),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_404),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_370),
.B1(n_375),
.B2(n_32),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_403),
.A2(n_390),
.B1(n_401),
.B2(n_405),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_399),
.Y(n_425)
);

OAI31xp33_ASAP7_75t_L g426 ( 
.A1(n_422),
.A2(n_417),
.A3(n_414),
.B(n_412),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

OAI33xp33_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_391),
.A3(n_402),
.B1(n_39),
.B2(n_40),
.B3(n_43),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_398),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_R g435 ( 
.A(n_418),
.B(n_37),
.Y(n_435)
);

OAI31xp33_ASAP7_75t_L g436 ( 
.A1(n_417),
.A2(n_46),
.A3(n_47),
.B(n_50),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_53),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_423),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_411),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_61),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_426),
.B(n_421),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_431),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_425),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_63),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_435),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_436),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_444),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_440),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_436),
.Y(n_455)
);

AOI21x1_ASAP7_75t_SL g456 ( 
.A1(n_451),
.A2(n_439),
.B(n_446),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_450),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_458),
.B(n_452),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_441),
.B1(n_442),
.B2(n_455),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_460),
.A2(n_443),
.B1(n_456),
.B2(n_430),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_81),
.C(n_83),
.Y(n_463)
);

OAI211xp5_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_85),
.B(n_86),
.C(n_88),
.Y(n_464)
);

AOI221xp5_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.C(n_92),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_94),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_465),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

OAI22x1_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_107),
.B1(n_108),
.B2(n_113),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_468),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_117),
.B(n_116),
.Y(n_473)
);


endmodule