module real_aes_16360_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_0), .A2(n_200), .B1(n_1147), .B2(n_1149), .Y(n_1182) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1), .Y(n_1032) );
XNOR2xp5_ASAP7_75t_L g1065 ( .A(n_2), .B(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g394 ( .A(n_3), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_4), .A2(n_244), .B1(n_723), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_4), .A2(n_177), .B1(n_666), .B2(n_837), .Y(n_836) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_5), .A2(n_408), .B(n_585), .C(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g754 ( .A(n_5), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_6), .A2(n_49), .B1(n_1147), .B2(n_1149), .Y(n_1172) );
INVx1_ASAP7_75t_L g633 ( .A(n_7), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_8), .A2(n_230), .B1(n_723), .B2(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_8), .A2(n_215), .B1(n_660), .B2(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g326 ( .A(n_9), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_9), .B(n_288), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_10), .A2(n_205), .B1(n_317), .B2(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_10), .A2(n_205), .B1(n_370), .B2(n_497), .Y(n_571) );
INVx1_ASAP7_75t_L g759 ( .A(n_11), .Y(n_759) );
INVx1_ASAP7_75t_L g692 ( .A(n_12), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_13), .A2(n_180), .B1(n_317), .B2(n_319), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_13), .A2(n_180), .B1(n_370), .B2(n_373), .Y(n_1055) );
INVx2_ASAP7_75t_L g1134 ( .A(n_14), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_14), .B(n_103), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_14), .B(n_1135), .Y(n_1154) );
OAI22xp33_ASAP7_75t_SL g1027 ( .A1(n_15), .A2(n_17), .B1(n_303), .B2(n_310), .Y(n_1027) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_15), .A2(n_17), .B1(n_576), .B2(n_1060), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_127), .B1(n_496), .B2(n_497), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_16), .A2(n_127), .B1(n_317), .B2(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_18), .A2(n_26), .B1(n_1152), .B2(n_1153), .Y(n_1164) );
INVx1_ASAP7_75t_L g1043 ( .A(n_19), .Y(n_1043) );
INVx1_ASAP7_75t_L g630 ( .A(n_20), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_21), .A2(n_157), .B1(n_319), .B2(n_593), .Y(n_967) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_21), .A2(n_255), .B1(n_372), .B2(n_694), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_22), .A2(n_119), .B1(n_1152), .B2(n_1153), .Y(n_1181) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_23), .Y(n_948) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_24), .A2(n_137), .B1(n_559), .B2(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_SL g598 ( .A1(n_24), .A2(n_137), .B1(n_372), .B2(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g416 ( .A(n_25), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_27), .A2(n_199), .B1(n_311), .B2(n_596), .Y(n_931) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_27), .A2(n_98), .B1(n_372), .B2(n_694), .Y(n_934) );
INVx1_ASAP7_75t_L g415 ( .A(n_28), .Y(n_415) );
INVx1_ASAP7_75t_L g847 ( .A(n_29), .Y(n_847) );
INVx1_ASAP7_75t_L g930 ( .A(n_30), .Y(n_930) );
OAI211xp5_ASAP7_75t_L g935 ( .A1(n_30), .A2(n_555), .B(n_601), .C(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g1080 ( .A(n_31), .Y(n_1080) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_32), .A2(n_97), .B1(n_1147), .B2(n_1158), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_33), .A2(n_100), .B1(n_1147), .B2(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1359 ( .A(n_34), .Y(n_1359) );
INVx1_ASAP7_75t_L g464 ( .A(n_35), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g953 ( .A(n_36), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_37), .Y(n_945) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_38), .A2(n_121), .B1(n_593), .B2(n_594), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_38), .A2(n_50), .B1(n_344), .B2(n_694), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_39), .A2(n_173), .B1(n_344), .B2(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_39), .A2(n_40), .B1(n_593), .B2(n_594), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_40), .A2(n_262), .B1(n_334), .B2(n_372), .Y(n_683) );
INVx1_ASAP7_75t_L g1072 ( .A(n_41), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1106 ( .A1(n_42), .A2(n_160), .B1(n_319), .B2(n_596), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_42), .A2(n_118), .B1(n_372), .B2(n_507), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_43), .A2(n_143), .B1(n_853), .B2(n_854), .Y(n_852) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_43), .Y(n_865) );
INVx1_ASAP7_75t_L g797 ( .A(n_44), .Y(n_797) );
INVx1_ASAP7_75t_L g591 ( .A(n_45), .Y(n_591) );
INVx1_ASAP7_75t_L g1103 ( .A(n_46), .Y(n_1103) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_46), .A2(n_601), .B(n_1110), .C(n_1111), .Y(n_1109) );
INVx1_ASAP7_75t_L g341 ( .A(n_47), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_47), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_48), .A2(n_125), .B1(n_1147), .B2(n_1158), .Y(n_1169) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_50), .A2(n_204), .B1(n_559), .B2(n_596), .Y(n_747) );
INVx1_ASAP7_75t_L g541 ( .A(n_51), .Y(n_541) );
XOR2x2_ASAP7_75t_L g843 ( .A(n_52), .B(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_52), .A2(n_217), .B1(n_1152), .B2(n_1153), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_53), .A2(n_76), .B1(n_723), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_53), .A2(n_238), .B1(n_608), .B2(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g534 ( .A(n_54), .Y(n_534) );
INVx1_ASAP7_75t_L g1084 ( .A(n_55), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_56), .A2(n_585), .B(n_927), .C(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g937 ( .A(n_56), .Y(n_937) );
INVx1_ASAP7_75t_L g1122 ( .A(n_57), .Y(n_1122) );
INVx1_ASAP7_75t_L g1044 ( .A(n_58), .Y(n_1044) );
INVx2_ASAP7_75t_L g337 ( .A(n_59), .Y(n_337) );
XNOR2x2_ASAP7_75t_L g524 ( .A(n_60), .B(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_61), .A2(n_236), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_61), .A2(n_174), .B1(n_726), .B2(n_728), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_62), .A2(n_220), .B1(n_303), .B2(n_568), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_62), .A2(n_220), .B1(n_507), .B2(n_576), .Y(n_575) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_63), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_63), .A2(n_143), .B1(n_564), .B2(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g1387 ( .A(n_64), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1398 ( .A1(n_64), .A2(n_164), .B1(n_319), .B2(n_596), .Y(n_1398) );
INVx1_ASAP7_75t_L g690 ( .A(n_65), .Y(n_690) );
INVx1_ASAP7_75t_L g746 ( .A(n_66), .Y(n_746) );
INVx1_ASAP7_75t_L g686 ( .A(n_67), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_68), .A2(n_252), .B1(n_334), .B2(n_344), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_68), .A2(n_252), .B1(n_593), .B2(n_594), .Y(n_1015) );
INVx1_ASAP7_75t_L g1356 ( .A(n_69), .Y(n_1356) );
OAI22xp33_ASAP7_75t_SL g1002 ( .A1(n_70), .A2(n_261), .B1(n_372), .B2(n_694), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_70), .A2(n_261), .B1(n_559), .B2(n_596), .Y(n_1010) );
INVx1_ASAP7_75t_L g535 ( .A(n_71), .Y(n_535) );
INVx1_ASAP7_75t_L g764 ( .A(n_72), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_73), .A2(n_98), .B1(n_304), .B2(n_319), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_73), .A2(n_199), .B1(n_334), .B2(n_344), .Y(n_938) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_74), .A2(n_355), .B(n_499), .C(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g517 ( .A(n_74), .Y(n_517) );
INVx1_ASAP7_75t_L g620 ( .A(n_75), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_76), .A2(n_86), .B1(n_608), .B2(n_839), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_77), .Y(n_911) );
INVx1_ASAP7_75t_L g402 ( .A(n_78), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_79), .A2(n_260), .B1(n_440), .B2(n_666), .C(n_670), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_79), .A2(n_132), .B1(n_731), .B2(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g988 ( .A(n_80), .Y(n_988) );
INVx1_ASAP7_75t_L g482 ( .A(n_81), .Y(n_482) );
INVx1_ASAP7_75t_L g590 ( .A(n_82), .Y(n_590) );
INVx1_ASAP7_75t_L g805 ( .A(n_83), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_83), .A2(n_237), .B1(n_618), .B2(n_811), .C(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g985 ( .A(n_84), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_85), .A2(n_156), .B1(n_593), .B2(n_594), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_85), .A2(n_156), .B1(n_334), .B2(n_344), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_86), .A2(n_238), .B1(n_726), .B2(n_876), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_87), .A2(n_106), .B1(n_1147), .B2(n_1149), .Y(n_1146) );
XOR2x2_ASAP7_75t_L g579 ( .A(n_88), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_89), .A2(n_120), .B1(n_1152), .B2(n_1153), .Y(n_1204) );
INVx1_ASAP7_75t_L g1360 ( .A(n_90), .Y(n_1360) );
INVx1_ASAP7_75t_L g530 ( .A(n_91), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g560 ( .A1(n_92), .A2(n_277), .B(n_561), .C(n_566), .Y(n_560) );
INVx1_ASAP7_75t_L g574 ( .A(n_92), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_93), .Y(n_1102) );
INVx1_ASAP7_75t_L g461 ( .A(n_94), .Y(n_461) );
INVx1_ASAP7_75t_L g898 ( .A(n_95), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_96), .A2(n_169), .B1(n_593), .B2(n_594), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_96), .A2(n_169), .B1(n_334), .B2(n_344), .Y(n_609) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_99), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_99), .B(n_1122), .Y(n_1132) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_101), .A2(n_215), .B1(n_820), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_101), .A2(n_230), .B1(n_829), .B2(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g1025 ( .A(n_102), .Y(n_1025) );
INVx1_ASAP7_75t_L g1135 ( .A(n_103), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_103), .B(n_1134), .Y(n_1148) );
INVx1_ASAP7_75t_L g1079 ( .A(n_104), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_105), .A2(n_167), .B1(n_1152), .B2(n_1153), .Y(n_1168) );
XOR2xp5_ASAP7_75t_L g1405 ( .A(n_107), .B(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g856 ( .A(n_108), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_109), .Y(n_950) );
INVx2_ASAP7_75t_L g382 ( .A(n_110), .Y(n_382) );
INVx1_ASAP7_75t_L g449 ( .A(n_110), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_111), .Y(n_904) );
INVx1_ASAP7_75t_L g768 ( .A(n_112), .Y(n_768) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_113), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_114), .A2(n_248), .B1(n_723), .B2(n_878), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_114), .A2(n_187), .B1(n_885), .B2(n_886), .Y(n_889) );
INVx1_ASAP7_75t_L g617 ( .A(n_115), .Y(n_617) );
INVx1_ASAP7_75t_L g994 ( .A(n_116), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_117), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_118), .A2(n_122), .B1(n_303), .B2(n_1105), .Y(n_1104) );
XNOR2xp5_ASAP7_75t_L g1017 ( .A(n_120), .B(n_1018), .Y(n_1017) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_121), .A2(n_204), .B1(n_334), .B2(n_372), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_122), .A2(n_160), .B1(n_373), .B2(n_1114), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_123), .A2(n_241), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g772 ( .A(n_124), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_126), .A2(n_129), .B1(n_1147), .B2(n_1149), .Y(n_1203) );
INVx1_ASAP7_75t_L g632 ( .A(n_128), .Y(n_632) );
INVx1_ASAP7_75t_L g1362 ( .A(n_130), .Y(n_1362) );
INVx1_ASAP7_75t_L g475 ( .A(n_131), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_132), .A2(n_213), .B1(n_440), .B2(n_666), .C(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g992 ( .A(n_133), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_134), .A2(n_136), .B1(n_1152), .B2(n_1153), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_135), .Y(n_964) );
INVx1_ASAP7_75t_L g769 ( .A(n_138), .Y(n_769) );
AOI31xp33_ASAP7_75t_L g657 ( .A1(n_139), .A2(n_658), .A3(n_682), .B(n_697), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g715 ( .A(n_139), .B(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_139), .Y(n_737) );
INVx1_ASAP7_75t_L g1007 ( .A(n_140), .Y(n_1007) );
OAI211xp5_ASAP7_75t_L g1011 ( .A1(n_140), .A2(n_584), .B(n_585), .C(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1038 ( .A(n_141), .Y(n_1038) );
INVx1_ASAP7_75t_L g1385 ( .A(n_142), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_142), .A2(n_249), .B1(n_303), .B2(n_568), .Y(n_1394) );
BUFx3_ASAP7_75t_L g339 ( .A(n_144), .Y(n_339) );
INVx1_ASAP7_75t_L g1381 ( .A(n_145), .Y(n_1381) );
OA211x2_ASAP7_75t_L g1395 ( .A1(n_145), .A2(n_284), .B(n_408), .C(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g986 ( .A(n_146), .Y(n_986) );
INVx1_ASAP7_75t_L g989 ( .A(n_147), .Y(n_989) );
INVx1_ASAP7_75t_L g762 ( .A(n_148), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_149), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_150), .A2(n_152), .B1(n_1152), .B2(n_1153), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_151), .Y(n_954) );
AOI222xp33_ASAP7_75t_L g1341 ( .A1(n_152), .A2(n_1342), .B1(n_1401), .B2(n_1404), .C1(n_1407), .C2(n_1409), .Y(n_1341) );
OAI22xp5_ASAP7_75t_SL g1344 ( .A1(n_152), .A2(n_1345), .B1(n_1392), .B2(n_1400), .Y(n_1344) );
NAND4xp25_ASAP7_75t_L g1345 ( .A(n_152), .B(n_1346), .C(n_1364), .D(n_1375), .Y(n_1345) );
INVx1_ASAP7_75t_L g505 ( .A(n_153), .Y(n_505) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_153), .A2(n_277), .B(n_515), .C(n_516), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_154), .Y(n_1006) );
INVx1_ASAP7_75t_L g532 ( .A(n_155), .Y(n_532) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_157), .A2(n_258), .B1(n_334), .B2(n_344), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_158), .Y(n_951) );
XNOR2x1_ASAP7_75t_L g980 ( .A(n_159), .B(n_981), .Y(n_980) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_161), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_162), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_163), .A2(n_224), .B1(n_1147), .B2(n_1149), .Y(n_1165) );
INVx1_ASAP7_75t_L g1384 ( .A(n_164), .Y(n_1384) );
INVx1_ASAP7_75t_L g1041 ( .A(n_165), .Y(n_1041) );
INVx1_ASAP7_75t_L g1082 ( .A(n_166), .Y(n_1082) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_167), .B(n_740), .Y(n_739) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_168), .A2(n_195), .B1(n_317), .B2(n_319), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_168), .A2(n_195), .B1(n_370), .B2(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g679 ( .A(n_170), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_170), .A2(n_236), .B1(n_719), .B2(n_723), .Y(n_718) );
INVx1_ASAP7_75t_L g539 ( .A(n_171), .Y(n_539) );
OAI211xp5_ASAP7_75t_L g1099 ( .A1(n_172), .A2(n_284), .B(n_1100), .C(n_1101), .Y(n_1099) );
INVx1_ASAP7_75t_L g1112 ( .A(n_172), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_173), .Y(n_701) );
INVx1_ASAP7_75t_L g676 ( .A(n_174), .Y(n_676) );
INVx1_ASAP7_75t_L g1074 ( .A(n_175), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1003 ( .A1(n_176), .A2(n_601), .B(n_1004), .C(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g1014 ( .A(n_176), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_177), .A2(n_240), .B1(n_820), .B2(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g1352 ( .A(n_178), .Y(n_1352) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_179), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g1031 ( .A(n_181), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_182), .Y(n_429) );
INVx1_ASAP7_75t_L g848 ( .A(n_183), .Y(n_848) );
INVx1_ASAP7_75t_L g774 ( .A(n_184), .Y(n_774) );
OAI211xp5_ASAP7_75t_SL g276 ( .A1(n_185), .A2(n_277), .B(n_284), .C(n_291), .Y(n_276) );
INVx1_ASAP7_75t_L g365 ( .A(n_185), .Y(n_365) );
INVx1_ASAP7_75t_L g397 ( .A(n_186), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_187), .A2(n_193), .B1(n_873), .B2(n_876), .Y(n_872) );
INVx1_ASAP7_75t_L g795 ( .A(n_188), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_189), .Y(n_947) );
INVx1_ASAP7_75t_L g1355 ( .A(n_190), .Y(n_1355) );
INVx1_ASAP7_75t_L g480 ( .A(n_191), .Y(n_480) );
INVx1_ASAP7_75t_L g473 ( .A(n_192), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_193), .A2(n_248), .B1(n_885), .B2(n_886), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_194), .Y(n_908) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
INVx1_ASAP7_75t_L g1351 ( .A(n_197), .Y(n_1351) );
INVx1_ASAP7_75t_L g802 ( .A(n_198), .Y(n_802) );
INVx1_ASAP7_75t_L g965 ( .A(n_201), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g970 ( .A1(n_201), .A2(n_555), .B(n_601), .C(n_971), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_202), .Y(n_903) );
INVx1_ASAP7_75t_L g745 ( .A(n_203), .Y(n_745) );
INVx1_ASAP7_75t_L g627 ( .A(n_206), .Y(n_627) );
INVx1_ASAP7_75t_L g991 ( .A(n_207), .Y(n_991) );
INVx1_ASAP7_75t_L g565 ( .A(n_208), .Y(n_565) );
OAI211xp5_ASAP7_75t_L g572 ( .A1(n_208), .A2(n_349), .B(n_355), .C(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g766 ( .A(n_209), .Y(n_766) );
INVx1_ASAP7_75t_L g296 ( .A(n_210), .Y(n_296) );
OA22x2_ASAP7_75t_L g791 ( .A1(n_211), .A2(n_792), .B1(n_841), .B2(n_842), .Y(n_791) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_211), .Y(n_842) );
INVx1_ASAP7_75t_L g468 ( .A(n_212), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_213), .A2(n_260), .B1(n_726), .B2(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g1026 ( .A(n_214), .Y(n_1026) );
OAI211xp5_ASAP7_75t_L g1056 ( .A1(n_214), .A2(n_349), .B(n_355), .C(n_1057), .Y(n_1056) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_216), .Y(n_929) );
INVx1_ASAP7_75t_L g407 ( .A(n_218), .Y(n_407) );
INVx1_ASAP7_75t_L g623 ( .A(n_219), .Y(n_623) );
BUFx3_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
INVx1_ASAP7_75t_L g309 ( .A(n_221), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_222), .A2(n_251), .B1(n_303), .B2(n_310), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_222), .A2(n_251), .B1(n_333), .B2(n_342), .Y(n_332) );
INVx1_ASAP7_75t_L g562 ( .A(n_223), .Y(n_562) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_225), .A2(n_247), .B1(n_507), .B2(n_508), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_225), .A2(n_247), .B1(n_303), .B2(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1380 ( .A(n_226), .Y(n_1380) );
INVx1_ASAP7_75t_L g1363 ( .A(n_227), .Y(n_1363) );
OAI211xp5_ASAP7_75t_L g962 ( .A1(n_228), .A2(n_585), .B(n_927), .C(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g972 ( .A(n_228), .Y(n_972) );
INVx1_ASAP7_75t_L g615 ( .A(n_229), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_231), .Y(n_915) );
INVx1_ASAP7_75t_L g995 ( .A(n_232), .Y(n_995) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_233), .A2(n_583), .B(n_585), .C(n_589), .Y(n_582) );
INVx1_ASAP7_75t_L g604 ( .A(n_233), .Y(n_604) );
INVx1_ASAP7_75t_L g330 ( .A(n_234), .Y(n_330) );
INVx2_ASAP7_75t_L g391 ( .A(n_234), .Y(n_391) );
INVx1_ASAP7_75t_L g448 ( .A(n_234), .Y(n_448) );
INVx1_ASAP7_75t_L g504 ( .A(n_235), .Y(n_504) );
OAI211xp5_ASAP7_75t_L g799 ( .A1(n_237), .A2(n_710), .B(n_800), .C(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g1070 ( .A(n_239), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_240), .A2(n_244), .B1(n_833), .B2(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_242), .A2(n_349), .B(n_355), .C(n_359), .Y(n_348) );
INVx1_ASAP7_75t_L g1035 ( .A(n_243), .Y(n_1035) );
INVx1_ASAP7_75t_L g542 ( .A(n_245), .Y(n_542) );
INVx1_ASAP7_75t_L g1076 ( .A(n_246), .Y(n_1076) );
INVx1_ASAP7_75t_L g1389 ( .A(n_249), .Y(n_1389) );
INVx1_ASAP7_75t_L g858 ( .A(n_250), .Y(n_858) );
INVx1_ASAP7_75t_L g1382 ( .A(n_253), .Y(n_1382) );
XNOR2xp5_ASAP7_75t_L g939 ( .A(n_254), .B(n_940), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_255), .A2(n_258), .B1(n_311), .B2(n_596), .Y(n_966) );
INVx1_ASAP7_75t_L g426 ( .A(n_256), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_257), .Y(n_918) );
OAI211xp5_ASAP7_75t_L g1021 ( .A1(n_259), .A2(n_566), .B(n_1022), .C(n_1024), .Y(n_1021) );
INVx1_ASAP7_75t_L g1058 ( .A(n_259), .Y(n_1058) );
INVx1_ASAP7_75t_L g699 ( .A(n_262), .Y(n_699) );
INVx1_ASAP7_75t_L g537 ( .A(n_263), .Y(n_537) );
INVx1_ASAP7_75t_L g460 ( .A(n_264), .Y(n_460) );
INVx1_ASAP7_75t_L g1036 ( .A(n_265), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_1116), .B(n_1128), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_975), .B1(n_976), .B2(n_1115), .Y(n_267) );
INVx1_ASAP7_75t_L g1115 ( .A(n_268), .Y(n_1115) );
XNOR2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_787), .Y(n_268) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_522), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B1(n_454), .B2(n_455), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_331), .C(n_386), .Y(n_274) );
OAI31xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_302), .A3(n_316), .B(n_323), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_279), .A2(n_1074), .B1(n_1075), .B2(n_1076), .Y(n_1073) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx4f_ASAP7_75t_L g491 ( .A(n_280), .Y(n_491) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_280), .Y(n_584) );
INVx4_ASAP7_75t_L g644 ( .A(n_280), .Y(n_644) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g410 ( .A(n_281), .Y(n_410) );
NAND2x1_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_282), .B(n_283), .Y(n_290) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
OR2x2_ASAP7_75t_L g307 ( .A(n_282), .B(n_283), .Y(n_307) );
INVx2_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_282), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g406 ( .A(n_282), .Y(n_406) );
BUFx2_ASAP7_75t_L g295 ( .A(n_283), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
OR2x2_ASAP7_75t_L g405 ( .A(n_283), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g722 ( .A(n_283), .Y(n_722) );
AND2x2_ASAP7_75t_L g724 ( .A(n_283), .B(n_315), .Y(n_724) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g515 ( .A(n_285), .Y(n_515) );
INVx1_ASAP7_75t_L g566 ( .A(n_285), .Y(n_566) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
AND2x2_ASAP7_75t_L g586 ( .A(n_286), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g594 ( .A(n_286), .B(n_313), .Y(n_594) );
AND2x2_ASAP7_75t_L g706 ( .A(n_286), .B(n_295), .Y(n_706) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVxp67_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g294 ( .A(n_288), .Y(n_294) );
AND2x4_ASAP7_75t_L g299 ( .A(n_288), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g419 ( .A(n_288), .B(n_326), .Y(n_419) );
BUFx3_ASAP7_75t_L g728 ( .A(n_289), .Y(n_728) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_289), .Y(n_822) );
BUFx3_ASAP7_75t_L g824 ( .A(n_289), .Y(n_824) );
BUFx3_ASAP7_75t_L g876 ( .A(n_289), .Y(n_876) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g588 ( .A(n_290), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_296), .B1(n_297), .B2(n_298), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_292), .A2(n_562), .B1(n_563), .B2(n_565), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_292), .A2(n_803), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_293), .A2(n_299), .B1(n_504), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_293), .A2(n_298), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_293), .A2(n_298), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g867 ( .A(n_293), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_293), .A2(n_803), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_293), .A2(n_563), .B1(n_1380), .B2(n_1382), .Y(n_1396) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OR2x2_ASAP7_75t_L g312 ( .A(n_294), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g869 ( .A(n_294), .B(n_733), .Y(n_869) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_294), .B(n_295), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_296), .A2(n_360), .B1(n_365), .B2(n_366), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_298), .A2(n_706), .B1(n_964), .B2(n_965), .Y(n_963) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g564 ( .A(n_299), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_299), .A2(n_686), .B1(n_690), .B2(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g804 ( .A(n_299), .Y(n_804) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x6_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
OR2x6_ASAP7_75t_L g317 ( .A(n_305), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g593 ( .A(n_305), .B(n_308), .Y(n_593) );
INVx1_ASAP7_75t_L g650 ( .A(n_305), .Y(n_650) );
BUFx4f_ASAP7_75t_L g1368 ( .A(n_305), .Y(n_1368) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx3_ASAP7_75t_L g396 ( .A(n_306), .Y(n_396) );
BUFx4f_ASAP7_75t_L g425 ( .A(n_306), .Y(n_425) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g320 ( .A(n_308), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g520 ( .A(n_312), .Y(n_520) );
INVx8_ASAP7_75t_L g400 ( .A(n_313), .Y(n_400) );
BUFx2_ASAP7_75t_L g1369 ( .A(n_313), .Y(n_1369) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g796 ( .A(n_317), .Y(n_796) );
OR2x6_ASAP7_75t_L g596 ( .A(n_318), .B(n_396), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_SL g513 ( .A(n_320), .Y(n_513) );
INVx4_ASAP7_75t_L g559 ( .A(n_320), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_320), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_320), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_320), .A2(n_847), .B1(n_848), .B2(n_861), .Y(n_860) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_321), .Y(n_727) );
BUFx3_ASAP7_75t_L g875 ( .A(n_321), .Y(n_875) );
OAI31xp33_ASAP7_75t_L g925 ( .A1(n_323), .A2(n_926), .A3(n_931), .B(n_932), .Y(n_925) );
OAI31xp33_ASAP7_75t_L g961 ( .A1(n_323), .A2(n_962), .A3(n_966), .B(n_967), .Y(n_961) );
OAI31xp33_ASAP7_75t_SL g1009 ( .A1(n_323), .A2(n_1010), .A3(n_1011), .B(n_1015), .Y(n_1009) );
OAI31xp33_ASAP7_75t_L g1098 ( .A1(n_323), .A2(n_1099), .A3(n_1104), .B(n_1106), .Y(n_1098) );
INVx1_ASAP7_75t_L g1399 ( .A(n_323), .Y(n_1399) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_SL g521 ( .A(n_324), .Y(n_521) );
BUFx3_ASAP7_75t_L g569 ( .A(n_324), .Y(n_569) );
INVx1_ASAP7_75t_L g711 ( .A(n_324), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g741 ( .A1(n_324), .A2(n_742), .A3(n_743), .B(n_747), .Y(n_741) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g1127 ( .A(n_325), .Y(n_1127) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_325), .B(n_1119), .Y(n_1403) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g385 ( .A(n_329), .Y(n_385) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI31xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_348), .A3(n_369), .B(n_379), .Y(n_331) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g507 ( .A(n_334), .Y(n_507) );
INVx2_ASAP7_75t_SL g857 ( .A(n_334), .Y(n_857) );
OR2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x4_ASAP7_75t_L g374 ( .A(n_335), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g695 ( .A(n_335), .B(n_375), .Y(n_695) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x6_ASAP7_75t_L g344 ( .A(n_336), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g356 ( .A(n_336), .B(n_357), .Y(n_356) );
OR2x4_ASAP7_75t_L g372 ( .A(n_336), .B(n_338), .Y(n_372) );
NAND3x1_ASAP7_75t_L g446 ( .A(n_336), .B(n_447), .C(n_449), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_336), .B(n_449), .Y(n_635) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_337), .B(n_382), .Y(n_433) );
BUFx3_ASAP7_75t_L g435 ( .A(n_338), .Y(n_435) );
BUFx3_ASAP7_75t_L g453 ( .A(n_338), .Y(n_453) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_338), .Y(n_616) );
INVx2_ASAP7_75t_L g778 ( .A(n_338), .Y(n_778) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_339), .B(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
AND2x4_ASAP7_75t_L g357 ( .A(n_339), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
INVx1_ASAP7_75t_L g664 ( .A(n_340), .Y(n_664) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g509 ( .A(n_344), .Y(n_509) );
INVx1_ASAP7_75t_L g577 ( .A(n_344), .Y(n_577) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_344), .Y(n_1114) );
BUFx3_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
INVx1_ASAP7_75t_L g471 ( .A(n_345), .Y(n_471) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g478 ( .A(n_346), .Y(n_478) );
INVx1_ASAP7_75t_L g353 ( .A(n_347), .Y(n_353) );
INVx2_ASAP7_75t_L g358 ( .A(n_347), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_349), .A2(n_397), .B1(n_416), .B2(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g481 ( .A(n_350), .Y(n_481) );
INVx1_ASAP7_75t_L g1033 ( .A(n_350), .Y(n_1033) );
INVx1_ASAP7_75t_L g1090 ( .A(n_350), .Y(n_1090) );
INVx1_ASAP7_75t_L g1110 ( .A(n_350), .Y(n_1110) );
INVx4_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_351), .Y(n_618) );
INVx3_ASAP7_75t_L g906 ( .A(n_351), .Y(n_906) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
BUFx2_ASAP7_75t_L g501 ( .A(n_352), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
BUFx2_ASAP7_75t_L g368 ( .A(n_353), .Y(n_368) );
BUFx2_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
AND2x4_ASAP7_75t_L g668 ( .A(n_354), .B(n_669), .Y(n_668) );
CKINVDCx8_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
CKINVDCx8_ASAP7_75t_R g601 ( .A(n_356), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_356), .B(n_809), .C(n_810), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g849 ( .A1(n_356), .A2(n_850), .B(n_851), .C(n_852), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_356), .B(n_1378), .Y(n_1377) );
BUFx3_ASAP7_75t_L g608 ( .A(n_357), .Y(n_608) );
BUFx2_ASAP7_75t_L g660 ( .A(n_357), .Y(n_660) );
INVx2_ASAP7_75t_L g688 ( .A(n_357), .Y(n_688) );
BUFx2_ASAP7_75t_L g752 ( .A(n_357), .Y(n_752) );
BUFx2_ASAP7_75t_L g851 ( .A(n_357), .Y(n_851) );
INVx1_ASAP7_75t_L g669 ( .A(n_358), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_360), .A2(n_366), .B1(n_1025), .B2(n_1058), .Y(n_1057) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g503 ( .A(n_361), .Y(n_503) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
AND2x4_ASAP7_75t_L g367 ( .A(n_362), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g603 ( .A(n_362), .B(n_364), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_362), .B(n_368), .Y(n_605) );
AND2x4_ASAP7_75t_L g691 ( .A(n_362), .B(n_364), .Y(n_691) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND3x4_ASAP7_75t_L g671 ( .A(n_363), .B(n_382), .C(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_366), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_366), .A2(n_503), .B1(n_562), .B2(n_574), .Y(n_573) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g811 ( .A(n_367), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_367), .A2(n_603), .B1(n_1102), .B2(n_1112), .Y(n_1111) );
AOI222xp33_ASAP7_75t_L g1379 ( .A1(n_367), .A2(n_660), .B1(n_691), .B2(n_1380), .C1(n_1381), .C2(n_1382), .Y(n_1379) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_372), .Y(n_496) );
INVx2_ASAP7_75t_SL g814 ( .A(n_372), .Y(n_814) );
INVx1_ASAP7_75t_L g1388 ( .A(n_372), .Y(n_1388) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g497 ( .A(n_374), .Y(n_497) );
INVx1_ASAP7_75t_L g599 ( .A(n_374), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_374), .A2(n_795), .B1(n_797), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_374), .A2(n_814), .B1(n_847), .B2(n_848), .Y(n_846) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
INVx1_ASAP7_75t_L g474 ( .A(n_375), .Y(n_474) );
INVx2_ASAP7_75t_L g834 ( .A(n_375), .Y(n_834) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_375), .Y(n_885) );
INVx2_ASAP7_75t_L g1094 ( .A(n_375), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_376), .Y(n_467) );
BUFx8_ASAP7_75t_L g622 ( .A(n_376), .Y(n_622) );
INVx2_ASAP7_75t_L g914 ( .A(n_376), .Y(n_914) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x4_ASAP7_75t_L g663 ( .A(n_378), .B(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_L g578 ( .A(n_379), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_379), .A2(n_521), .B1(n_845), .B2(n_859), .C(n_870), .Y(n_844) );
OAI31xp33_ASAP7_75t_L g1054 ( .A1(n_379), .A2(n_1055), .A3(n_1056), .B(n_1059), .Y(n_1054) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_380), .B(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g510 ( .A(n_380), .B(n_383), .Y(n_510) );
AND2x2_ASAP7_75t_L g610 ( .A(n_380), .B(n_383), .Y(n_610) );
AND2x2_ASAP7_75t_L g696 ( .A(n_380), .B(n_383), .Y(n_696) );
AND2x4_ASAP7_75t_L g1391 ( .A(n_380), .B(n_383), .Y(n_1391) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
OR2x2_ASAP7_75t_L g432 ( .A(n_385), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_SL g647 ( .A(n_385), .B(n_419), .Y(n_647) );
NOR2xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_430), .Y(n_386) );
OAI33xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .A3(n_401), .B1(n_411), .B2(n_417), .B3(n_422), .Y(n_387) );
INVx2_ASAP7_75t_SL g717 ( .A(n_388), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_388), .A2(n_1069), .A3(n_1073), .B1(n_1077), .B2(n_1081), .B3(n_1085), .Y(n_1068) );
INVx4_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g485 ( .A(n_389), .Y(n_485) );
INVx2_ASAP7_75t_L g528 ( .A(n_389), .Y(n_528) );
INVx2_ASAP7_75t_L g639 ( .A(n_389), .Y(n_639) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g634 ( .A(n_390), .B(n_635), .Y(n_634) );
OR2x6_ASAP7_75t_L g681 ( .A(n_390), .B(n_635), .Y(n_681) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g672 ( .A(n_391), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_397), .B2(n_398), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_394), .A2(n_415), .B1(n_435), .B2(n_436), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_395), .A2(n_398), .B1(n_468), .B2(n_475), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_395), .A2(n_398), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_395), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g529 ( .A1(n_398), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_529) );
INVx6_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
INVx1_ASAP7_75t_L g488 ( .A(n_400), .Y(n_488) );
INVx4_ASAP7_75t_L g651 ( .A(n_400), .Y(n_651) );
INVx2_ASAP7_75t_L g761 ( .A(n_400), .Y(n_761) );
INVx2_ASAP7_75t_SL g773 ( .A(n_400), .Y(n_773) );
INVx2_ASAP7_75t_L g1083 ( .A(n_400), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_407), .B2(n_408), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_402), .A2(n_426), .B1(n_439), .B2(n_441), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_403), .A2(n_410), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g1052 ( .A(n_403), .Y(n_1052) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g765 ( .A(n_404), .Y(n_765) );
BUFx2_ASAP7_75t_L g1373 ( .A(n_404), .Y(n_1373) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g414 ( .A(n_405), .Y(n_414) );
INVx1_ASAP7_75t_L g642 ( .A(n_405), .Y(n_642) );
BUFx2_ASAP7_75t_L g923 ( .A(n_405), .Y(n_923) );
AND2x2_ASAP7_75t_L g721 ( .A(n_406), .B(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_429), .B1(n_441), .B2(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_408), .A2(n_412), .B1(n_1035), .B2(n_1038), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_408), .A2(n_1032), .B1(n_1044), .B2(n_1051), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_408), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
INVx5_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_410), .A2(n_412), .B1(n_415), .B2(n_416), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_410), .A2(n_412), .B1(n_461), .B2(n_482), .Y(n_492) );
BUFx2_ASAP7_75t_SL g538 ( .A(n_410), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_410), .A2(n_617), .B1(n_633), .B2(n_641), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_410), .A2(n_904), .B1(n_918), .B2(n_923), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_410), .A2(n_765), .B1(n_947), .B2(n_948), .Y(n_946) );
BUFx3_ASAP7_75t_L g1023 ( .A(n_410), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_412), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx4_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
INVx2_ASAP7_75t_L g1075 ( .A(n_413), .Y(n_1075) );
INVx4_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI33xp33_ASAP7_75t_L g483 ( .A1(n_417), .A2(n_484), .A3(n_486), .B1(n_489), .B2(n_492), .B3(n_493), .Y(n_483) );
OAI33xp33_ASAP7_75t_L g527 ( .A1(n_417), .A2(n_528), .A3(n_529), .B1(n_533), .B2(n_536), .B3(n_540), .Y(n_527) );
OAI33xp33_ASAP7_75t_L g1045 ( .A1(n_417), .A2(n_485), .A3(n_1046), .B1(n_1049), .B2(n_1050), .B3(n_1053), .Y(n_1045) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g880 ( .A(n_418), .B(n_881), .C(n_882), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_418), .Y(n_1085) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_423), .A2(n_427), .B1(n_1036), .B2(n_1041), .Y(n_1053) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g487 ( .A(n_424), .Y(n_487) );
INVx3_ASAP7_75t_L g1071 ( .A(n_424), .Y(n_1071) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g531 ( .A(n_425), .Y(n_531) );
INVx4_ASAP7_75t_L g638 ( .A(n_425), .Y(n_638) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_428), .A2(n_638), .B1(n_988), .B2(n_991), .Y(n_997) );
OAI33xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .A3(n_438), .B1(n_442), .B2(n_444), .B3(n_450), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g458 ( .A1(n_431), .A2(n_444), .A3(n_459), .B1(n_463), .B2(n_472), .B3(n_479), .Y(n_458) );
OAI33xp33_ASAP7_75t_L g1086 ( .A1(n_431), .A2(n_1087), .A3(n_1091), .B1(n_1093), .B2(n_1095), .B3(n_1096), .Y(n_1086) );
BUFx8_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_432), .Y(n_544) );
BUFx4f_ASAP7_75t_L g613 ( .A(n_432), .Y(n_613) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_432), .Y(n_1348) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_435), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_435), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_435), .A2(n_1004), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_435), .A2(n_618), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_437), .Y(n_462) );
INVx2_ASAP7_75t_L g549 ( .A(n_437), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_437), .A2(n_616), .B1(n_632), .B2(n_633), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_437), .A2(n_759), .B1(n_768), .B2(n_777), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_437), .A2(n_777), .B1(n_917), .B2(n_918), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_437), .A2(n_777), .B1(n_945), .B2(n_951), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_437), .A2(n_616), .B1(n_991), .B2(n_992), .Y(n_990) );
BUFx6f_ASAP7_75t_L g1004 ( .A(n_437), .Y(n_1004) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_441), .A2(n_535), .B1(n_542), .B2(n_552), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_441), .A2(n_443), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_441), .A2(n_1038), .B1(n_1039), .B2(n_1041), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_441), .A2(n_1074), .B1(n_1082), .B2(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_443), .A2(n_766), .B1(n_774), .B2(n_783), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_443), .A2(n_781), .B1(n_908), .B2(n_909), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_443), .A2(n_781), .B1(n_947), .B2(n_953), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g553 ( .A(n_445), .Y(n_553) );
INVx2_ASAP7_75t_L g1095 ( .A(n_445), .Y(n_1095) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g891 ( .A(n_446), .Y(n_891) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_453), .Y(n_547) );
INVx1_ASAP7_75t_L g1089 ( .A(n_453), .Y(n_1089) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_494), .C(n_511), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_483), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_460), .A2(n_480), .B1(n_487), .B2(n_488), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_464), .A2(n_473), .B1(n_490), .B2(n_491), .Y(n_489) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_466), .A2(n_476), .B1(n_534), .B2(n_541), .Y(n_550) );
INVx8_ASAP7_75t_L g1040 ( .A(n_466), .Y(n_1040) );
INVx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g552 ( .A(n_467), .Y(n_552) );
INVx3_ASAP7_75t_L g780 ( .A(n_467), .Y(n_780) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g624 ( .A(n_471), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_472) );
INVx1_ASAP7_75t_L g837 ( .A(n_474), .Y(n_837) );
OAI22xp33_ASAP7_75t_SL g1093 ( .A1(n_476), .A2(n_1076), .B1(n_1084), .B2(n_1094), .Y(n_1093) );
CKINVDCx8_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g781 ( .A(n_477), .Y(n_781) );
INVx3_ASAP7_75t_L g783 ( .A(n_477), .Y(n_783) );
INVx3_ASAP7_75t_L g959 ( .A(n_477), .Y(n_959) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g629 ( .A(n_478), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_481), .A2(n_616), .B1(n_762), .B2(n_769), .Y(n_784) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI33xp33_ASAP7_75t_L g757 ( .A1(n_485), .A2(n_758), .A3(n_763), .B1(n_767), .B2(n_770), .B3(n_771), .Y(n_757) );
OAI33xp33_ASAP7_75t_L g942 ( .A1(n_485), .A2(n_770), .A3(n_943), .B1(n_946), .B2(n_949), .B3(n_952), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_488), .A2(n_615), .B1(n_632), .B2(n_638), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_488), .A2(n_1031), .B1(n_1043), .B2(n_1047), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_491), .A2(n_765), .B1(n_768), .B2(n_769), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_491), .A2(n_923), .B1(n_985), .B2(n_994), .Y(n_998) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .A3(n_506), .B(n_510), .Y(n_494) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_509), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g1107 ( .A1(n_510), .A2(n_1108), .A3(n_1109), .B(n_1113), .Y(n_1107) );
OAI31xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_514), .A3(n_518), .B(n_521), .Y(n_511) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_520), .A2(n_856), .B1(n_858), .B2(n_869), .Y(n_868) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_520), .Y(n_1105) );
OAI31xp33_ASAP7_75t_SL g581 ( .A1(n_521), .A2(n_582), .A3(n_592), .B(n_595), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_654), .B1(n_785), .B2(n_786), .Y(n_522) );
INVx1_ASAP7_75t_L g785 ( .A(n_523), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_579), .B1(n_652), .B2(n_653), .Y(n_523) );
INVx1_ASAP7_75t_L g653 ( .A(n_524), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_557), .C(n_570), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_543), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_530), .A2(n_537), .B1(n_546), .B2(n_548), .Y(n_545) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_531), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_532), .A2(n_539), .B1(n_546), .B2(n_555), .Y(n_554) );
OAI33xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .A3(n_550), .B1(n_551), .B2(n_553), .B3(n_554), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_546), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_552), .A2(n_948), .B1(n_954), .B2(n_959), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_552), .A2(n_624), .B1(n_994), .B2(n_995), .Y(n_993) );
OAI33xp33_ASAP7_75t_L g1029 ( .A1(n_553), .A2(n_613), .A3(n_1030), .B1(n_1034), .B2(n_1037), .B3(n_1042), .Y(n_1029) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI31xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .A3(n_567), .B(n_569), .Y(n_557) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI31xp33_ASAP7_75t_L g1019 ( .A1(n_569), .A2(n_1020), .A3(n_1021), .B(n_1027), .Y(n_1019) );
OAI31xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .A3(n_575), .B(n_578), .Y(n_570) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_577), .A2(n_695), .B1(n_1384), .B2(n_1385), .Y(n_1383) );
INVx2_ASAP7_75t_SL g652 ( .A(n_579), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_597), .C(n_611), .Y(n_580) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_584), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_584), .A2(n_765), .B1(n_950), .B2(n_951), .Y(n_949) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g710 ( .A(n_586), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g862 ( .A1(n_586), .A2(n_863), .B(n_865), .C(n_866), .Y(n_862) );
INVx1_ASAP7_75t_L g709 ( .A(n_587), .Y(n_709) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g864 ( .A(n_588), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_590), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_591), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g700 ( .A(n_596), .Y(n_700) );
INVx1_ASAP7_75t_L g861 ( .A(n_596), .Y(n_861) );
OAI31xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .A3(n_609), .B(n_610), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .C(n_606), .Y(n_600) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_601), .B(n_685), .C(n_689), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g750 ( .A(n_601), .B(n_751), .C(n_753), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_605), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_605), .A2(n_691), .B1(n_745), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g854 ( .A(n_605), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_605), .A2(n_691), .B1(n_929), .B2(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_605), .A2(n_691), .B1(n_964), .B2(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_605), .A2(n_691), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g675 ( .A(n_608), .Y(n_675) );
OAI31xp33_ASAP7_75t_SL g933 ( .A1(n_610), .A2(n_934), .A3(n_935), .B(n_938), .Y(n_933) );
OAI31xp33_ASAP7_75t_SL g968 ( .A1(n_610), .A2(n_969), .A3(n_970), .B(n_973), .Y(n_968) );
OAI31xp33_ASAP7_75t_L g1001 ( .A1(n_610), .A2(n_1002), .A3(n_1003), .B(n_1008), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_636), .Y(n_611) );
OAI33xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .A3(n_619), .B1(n_625), .B2(n_631), .B3(n_634), .Y(n_612) );
OAI33xp33_ASAP7_75t_L g775 ( .A1(n_613), .A2(n_634), .A3(n_776), .B1(n_779), .B2(n_782), .B3(n_784), .Y(n_775) );
OAI33xp33_ASAP7_75t_L g901 ( .A1(n_613), .A2(n_634), .A3(n_902), .B1(n_907), .B2(n_910), .B3(n_916), .Y(n_901) );
OAI33xp33_ASAP7_75t_L g955 ( .A1(n_613), .A2(n_634), .A3(n_956), .B1(n_957), .B2(n_958), .B3(n_960), .Y(n_955) );
OAI33xp33_ASAP7_75t_L g983 ( .A1(n_613), .A2(n_634), .A3(n_984), .B1(n_987), .B2(n_990), .B3(n_993), .Y(n_983) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_616), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_902) );
OAI22xp5_ASAP7_75t_SL g987 ( .A1(n_616), .A2(n_905), .B1(n_988), .B2(n_989), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_618), .A2(n_777), .B1(n_944), .B2(n_950), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_623), .B2(n_624), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_620), .A2(n_627), .B1(n_641), .B2(n_643), .Y(n_640) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g626 ( .A(n_622), .Y(n_626) );
INVx3_ASAP7_75t_L g1358 ( .A(n_622), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_623), .A2(n_630), .B1(n_649), .B2(n_651), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_624), .A2(n_911), .B1(n_912), .B2(n_915), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_628), .B2(n_630), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_628), .A2(n_1354), .B1(n_1355), .B2(n_1356), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_628), .A2(n_1358), .B1(n_1359), .B2(n_1360), .Y(n_1357) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI33xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .A3(n_640), .B1(n_645), .B2(n_646), .B3(n_648), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_638), .A2(n_759), .B1(n_760), .B2(n_762), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_638), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_638), .A2(n_760), .B1(n_903), .B2(n_917), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_638), .A2(n_651), .B1(n_909), .B2(n_915), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_638), .A2(n_773), .B1(n_944), .B2(n_945), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_638), .A2(n_760), .B1(n_953), .B2(n_954), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_638), .A2(n_651), .B1(n_986), .B2(n_995), .Y(n_1000) );
OAI33xp33_ASAP7_75t_L g919 ( .A1(n_639), .A2(n_770), .A3(n_920), .B1(n_921), .B2(n_922), .B3(n_924), .Y(n_919) );
OAI33xp33_ASAP7_75t_L g996 ( .A1(n_639), .A2(n_646), .A3(n_997), .B1(n_998), .B2(n_999), .B3(n_1000), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_641), .A2(n_643), .B1(n_989), .B2(n_992), .Y(n_999) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g1078 ( .A(n_642), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_643), .A2(n_765), .B1(n_908), .B2(n_911), .Y(n_921) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g800 ( .A(n_644), .Y(n_800) );
INVx1_ASAP7_75t_L g927 ( .A(n_644), .Y(n_927) );
INVx2_ASAP7_75t_L g1100 ( .A(n_644), .Y(n_1100) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI33xp33_ASAP7_75t_L g716 ( .A1(n_647), .A2(n_717), .A3(n_718), .B1(n_725), .B2(n_729), .B3(n_730), .Y(n_716) );
INVx2_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
AOI33xp33_ASAP7_75t_L g816 ( .A1(n_647), .A2(n_717), .A3(n_817), .B1(n_819), .B2(n_823), .B3(n_825), .Y(n_816) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g786 ( .A(n_654), .Y(n_786) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
XNOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_739), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_712), .Y(n_656) );
INVx1_ASAP7_75t_L g714 ( .A(n_658), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_665), .B(n_673), .Y(n_658) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx8_ASAP7_75t_L g839 ( .A(n_662), .Y(n_839) );
INVx8_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx3_ASAP7_75t_L g678 ( .A(n_663), .Y(n_678) );
BUFx3_ASAP7_75t_L g830 ( .A(n_663), .Y(n_830) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_R g835 ( .A(n_667), .Y(n_835) );
INVx5_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx12f_ASAP7_75t_L g886 ( .A(n_668), .Y(n_886) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI33xp33_ASAP7_75t_L g827 ( .A1(n_671), .A2(n_828), .A3(n_832), .B1(n_836), .B2(n_838), .B3(n_840), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_671), .B(n_884), .C(n_887), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_674) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g840 ( .A(n_681), .Y(n_840) );
OAI33xp33_ASAP7_75t_L g1347 ( .A1(n_681), .A2(n_1348), .A3(n_1349), .B1(n_1353), .B2(n_1357), .B3(n_1361), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_682), .B(n_697), .Y(n_713) );
OAI31xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .A3(n_693), .B(n_696), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g831 ( .A(n_688), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_691), .B(n_802), .Y(n_812) );
INVx1_ASAP7_75t_L g853 ( .A(n_691), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_692), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI31xp33_ASAP7_75t_SL g748 ( .A1(n_696), .A2(n_749), .A3(n_750), .B(n_755), .Y(n_748) );
INVx1_ASAP7_75t_L g815 ( .A(n_696), .Y(n_815) );
AO21x1_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B(n_711), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .C(n_710), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_706), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_706), .A2(n_803), .B1(n_929), .B2(n_930), .Y(n_928) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AO21x1_ASAP7_75t_L g793 ( .A1(n_711), .A2(n_794), .B(n_798), .Y(n_793) );
OAI31xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .A3(n_715), .B(n_736), .Y(n_712) );
INVx1_ASAP7_75t_L g738 ( .A(n_716), .Y(n_738) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_717), .Y(n_879) );
INVx1_ASAP7_75t_L g1366 ( .A(n_717), .Y(n_1366) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g878 ( .A(n_720), .Y(n_878) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_721), .Y(n_733) );
BUFx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g735 ( .A(n_724), .Y(n_735) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g821 ( .A(n_727), .Y(n_821) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_SL g826 ( .A(n_732), .Y(n_826) );
INVx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_733), .Y(n_818) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND3xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_748), .C(n_756), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_746), .B(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_775), .Y(n_756) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_764), .A2(n_772), .B1(n_780), .B2(n_781), .Y(n_779) );
OAI33xp33_ASAP7_75t_L g1365 ( .A1(n_770), .A2(n_1366), .A3(n_1367), .B1(n_1370), .B2(n_1371), .B3(n_1374), .Y(n_1365) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_773), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_773), .A2(n_1356), .B1(n_1360), .B2(n_1368), .Y(n_1374) );
INVx2_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx3_ASAP7_75t_L g1350 ( .A(n_778), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_780), .A2(n_783), .B1(n_985), .B2(n_986), .Y(n_984) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B1(n_895), .B2(n_974), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
XNOR2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_843), .Y(n_790) );
INVx1_ASAP7_75t_L g841 ( .A(n_792), .Y(n_841) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_793), .B(n_807), .C(n_816), .D(n_827), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_796), .B(n_1127), .Y(n_1126) );
AND2x4_ASAP7_75t_SL g1402 ( .A(n_796), .B(n_1403), .Y(n_1402) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_806), .Y(n_798) );
OAI22xp5_ASAP7_75t_SL g1370 ( .A1(n_800), .A2(n_923), .B1(n_1355), .B2(n_1359), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_800), .A2(n_1352), .B1(n_1363), .B2(n_1372), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_803), .A2(n_1006), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AO21x1_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_813), .B(n_815), .Y(n_807) );
INVx2_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
BUFx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g894 ( .A(n_830), .Y(n_894) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .C(n_855), .Y(n_845) );
INVx2_ASAP7_75t_L g1060 ( .A(n_857), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1386 ( .A1(n_857), .A2(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1386) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .C(n_868), .Y(n_859) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_880), .C(n_883), .D(n_888), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_877), .C(n_879), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .C(n_892), .Y(n_888) );
BUFx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
BUFx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g974 ( .A(n_896), .Y(n_974) );
XNOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_939), .Y(n_896) );
XNOR2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
AND3x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_925), .C(n_933), .Y(n_899) );
NOR2xp33_ASAP7_75t_SL g900 ( .A(n_901), .B(n_919), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_905), .A2(n_1350), .B1(n_1351), .B2(n_1352), .Y(n_1349) );
INVx3_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g1097 ( .A(n_906), .Y(n_1097) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g1092 ( .A(n_913), .Y(n_1092) );
INVx3_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
BUFx2_ASAP7_75t_L g1354 ( .A(n_914), .Y(n_1354) );
AND3x1_ASAP7_75t_L g940 ( .A(n_941), .B(n_961), .C(n_968), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_955), .Y(n_941) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_1062), .B2(n_1063), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B1(n_1016), .B2(n_1061), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AND3x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_1001), .C(n_1009), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_983), .B(n_996), .Y(n_982) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1016), .Y(n_1061) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
AND3x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1028), .C(n_1054), .Y(n_1018) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
NOR2xp33_ASAP7_75t_SL g1028 ( .A(n_1029), .B(n_1045), .Y(n_1028) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1098), .C(n_1107), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1086), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_1070), .A2(n_1079), .B1(n_1088), .B2(n_1090), .Y(n_1087) );
OAI22xp33_ASAP7_75t_L g1096 ( .A1(n_1072), .A2(n_1080), .B1(n_1088), .B2(n_1097), .Y(n_1096) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
BUFx4f_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx3_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1125), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NOR2xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1123), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1408 ( .A(n_1121), .B(n_1124), .Y(n_1408) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1121), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1413 ( .A(n_1124), .B(n_1410), .Y(n_1413) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1136), .B(n_1341), .Y(n_1128) );
CKINVDCx20_ASAP7_75t_R g1129 ( .A(n_1130), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
AND2x6_ASAP7_75t_L g1147 ( .A(n_1132), .B(n_1148), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1132), .B(n_1150), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1132), .B(n_1133), .Y(n_1152) );
AND2x6_ASAP7_75t_L g1153 ( .A(n_1132), .B(n_1154), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1132), .B(n_1150), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1132), .B(n_1150), .Y(n_1218) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1133), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
AND4x1_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1259), .C(n_1289), .D(n_1318), .Y(n_1136) );
AOI211xp5_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1201), .B(n_1205), .C(n_1244), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
A2O1A1Ixp33_ASAP7_75t_L g1272 ( .A1(n_1139), .A2(n_1230), .B(n_1234), .C(n_1273), .Y(n_1272) );
NOR2xp33_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1189), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1183), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1160), .B1(n_1173), .B2(n_1176), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1142), .B(n_1184), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1142), .B(n_1162), .Y(n_1283) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1155), .Y(n_1143) );
OAI32xp33_ASAP7_75t_L g1212 ( .A1(n_1144), .A2(n_1213), .A3(n_1215), .B1(n_1220), .B2(n_1222), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1144), .B(n_1162), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1144), .B(n_1298), .Y(n_1297) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1144), .Y(n_1316) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1145), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1145), .B(n_1162), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1145), .B(n_1156), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1145), .B(n_1155), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1151), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1155), .B(n_1201), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1155), .B(n_1216), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1155), .B(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1155), .B(n_1202), .Y(n_1280) );
OAI32xp33_ASAP7_75t_L g1294 ( .A1(n_1155), .A2(n_1156), .A3(n_1227), .B1(n_1295), .B2(n_1297), .Y(n_1294) );
HB1xp67_ASAP7_75t_SL g1319 ( .A(n_1155), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1156), .B(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1156), .B(n_1239), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1156), .B(n_1202), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1156), .B(n_1163), .Y(n_1328) );
AND2x4_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1159), .Y(n_1156) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1161), .B(n_1198), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1166), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1162), .B(n_1223), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1162), .B(n_1198), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1162), .B(n_1228), .Y(n_1301) );
CKINVDCx14_ASAP7_75t_R g1308 ( .A(n_1162), .Y(n_1308) );
INVx3_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_1163), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1163), .B(n_1180), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1163), .B(n_1166), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1163), .B(n_1285), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1163), .B(n_1195), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1305 ( .A(n_1163), .B(n_1186), .Y(n_1305) );
AND2x4_ASAP7_75t_SL g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1166), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1166), .B(n_1198), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1166), .B(n_1188), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1166), .B(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1170), .Y(n_1166) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1167), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1167), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1167), .B(n_1198), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_1167), .B(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1167), .B(n_1180), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1167), .B(n_1180), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1170), .Y(n_1187) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1170), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1170), .B(n_1198), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1170), .B(n_1179), .Y(n_1250) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1170), .Y(n_1282) );
NAND2x1_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1173), .B(n_1239), .Y(n_1258) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1174), .B(n_1177), .Y(n_1200) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1174), .Y(n_1303) );
OAI21xp33_ASAP7_75t_L g1190 ( .A1(n_1175), .A2(n_1191), .B(n_1194), .Y(n_1190) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1175), .Y(n_1208) );
OAI21xp5_ASAP7_75t_L g1302 ( .A1(n_1176), .A2(n_1191), .B(n_1303), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1177), .B(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1177), .B(n_1195), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1177), .B(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1177), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1177), .B(n_1315), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1177), .B(n_1306), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1179), .B(n_1193), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1180), .B(n_1193), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1180), .B(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1180), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1180), .B(n_1211), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1180), .B(n_1293), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1180), .B(n_1250), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1184), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1188), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1185), .B(n_1198), .Y(n_1223) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1186), .B(n_1198), .Y(n_1291) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1188), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1188), .B(n_1195), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1196), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1245 ( .A1(n_1191), .A2(n_1194), .B1(n_1209), .B2(n_1246), .C(n_1247), .Y(n_1245) );
NOR2xp33_ASAP7_75t_SL g1327 ( .A(n_1192), .B(n_1223), .Y(n_1327) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_1195), .A2(n_1197), .B(n_1199), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1195), .B(n_1268), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1277 ( .A1(n_1195), .A2(n_1226), .B1(n_1250), .B2(n_1278), .C(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1195), .Y(n_1340) );
A2O1A1Ixp33_ASAP7_75t_L g1252 ( .A1(n_1197), .A2(n_1253), .B(n_1254), .C(n_1255), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1198), .B(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1198), .B(n_1282), .Y(n_1336) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_1200), .A2(n_1339), .B(n_1340), .Y(n_1338) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_1201), .A2(n_1237), .B1(n_1292), .B2(n_1332), .C(n_1335), .Y(n_1331) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1202), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1202), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
NAND4xp25_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1224), .C(n_1232), .D(n_1235), .Y(n_1205) );
O2A1O1Ixp33_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1209), .B(n_1210), .C(n_1212), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1208), .B(n_1239), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1208), .B(n_1275), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1208), .B(n_1296), .Y(n_1323) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1209), .Y(n_1265) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1214), .Y(n_1315) );
INVxp67_ASAP7_75t_SL g1317 ( .A(n_1215), .Y(n_1317) );
INVx3_ASAP7_75t_L g1231 ( .A(n_1216), .Y(n_1231) );
NAND3xp33_ASAP7_75t_SL g1274 ( .A(n_1216), .B(n_1234), .C(n_1275), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1216), .B(n_1239), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1219), .Y(n_1216) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1221), .Y(n_1278) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
OAI211xp5_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1227), .B(n_1228), .C(n_1230), .Y(n_1224) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
A2O1A1Ixp33_ASAP7_75t_L g1266 ( .A1(n_1229), .A2(n_1230), .B(n_1267), .C(n_1270), .Y(n_1266) );
A2O1A1Ixp33_ASAP7_75t_L g1290 ( .A1(n_1229), .A2(n_1291), .B(n_1292), .C(n_1294), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1330 ( .A(n_1229), .B(n_1310), .Y(n_1330) );
AOI21xp33_ASAP7_75t_L g1304 ( .A1(n_1230), .A2(n_1305), .B(n_1306), .Y(n_1304) );
CKINVDCx14_ASAP7_75t_R g1230 ( .A(n_1231), .Y(n_1230) );
AOI31xp33_ASAP7_75t_L g1244 ( .A1(n_1231), .A2(n_1245), .A3(n_1252), .B(n_1256), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1231), .B(n_1238), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1312 ( .A1(n_1231), .A2(n_1313), .B(n_1316), .Y(n_1312) );
A2O1A1Ixp33_ASAP7_75t_L g1335 ( .A1(n_1231), .A2(n_1336), .B(n_1337), .C(n_1338), .Y(n_1335) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1241), .Y(n_1235) );
A2O1A1Ixp33_ASAP7_75t_L g1259 ( .A1(n_1236), .A2(n_1260), .B(n_1262), .C(n_1272), .Y(n_1259) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1240), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1248 ( .A(n_1239), .B(n_1249), .C(n_1251), .Y(n_1248) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1239), .Y(n_1275) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1240), .Y(n_1306) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1262 ( .A1(n_1242), .A2(n_1263), .B1(n_1264), .B2(n_1265), .C(n_1266), .Y(n_1262) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1243), .B(n_1269), .Y(n_1326) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1250), .B(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1254), .Y(n_1339) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1255), .Y(n_1264) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1261), .B(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
CKINVDCx14_ASAP7_75t_R g1270 ( .A(n_1271), .Y(n_1270) );
A2O1A1O1Ixp25_ASAP7_75t_L g1318 ( .A1(n_1271), .A2(n_1319), .B(n_1320), .C(n_1321), .D(n_1331), .Y(n_1318) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1276), .B1(n_1277), .B2(n_1280), .C(n_1281), .Y(n_1273) );
AOI21xp5_ASAP7_75t_L g1289 ( .A1(n_1275), .A2(n_1290), .B(n_1299), .Y(n_1289) );
O2A1O1Ixp33_ASAP7_75t_L g1281 ( .A1(n_1282), .A2(n_1283), .B(n_1284), .C(n_1286), .Y(n_1281) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1283), .Y(n_1337) );
NOR2xp33_ASAP7_75t_SL g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1297), .Y(n_1311) );
AOI331xp33_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1302), .A3(n_1304), .B1(n_1307), .B2(n_1311), .B3(n_1312), .C1(n_1317), .Y(n_1299) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1307), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
NOR2xp33_ASAP7_75t_SL g1324 ( .A(n_1316), .B(n_1325), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_1322), .A2(n_1324), .B1(n_1327), .B2(n_1328), .C(n_1329), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVxp67_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVxp67_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
HB1xp67_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVxp67_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
NOR4xp25_ASAP7_75t_L g1400 ( .A(n_1347), .B(n_1365), .C(n_1376), .D(n_1392), .Y(n_1400) );
OAI22xp33_ASAP7_75t_L g1367 ( .A1(n_1351), .A2(n_1362), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
INVxp67_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx4_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVxp67_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
AOI31xp33_ASAP7_75t_L g1376 ( .A1(n_1377), .A2(n_1383), .A3(n_1386), .B(n_1390), .Y(n_1376) );
INVxp67_ASAP7_75t_SL g1378 ( .A(n_1379), .Y(n_1378) );
CKINVDCx14_ASAP7_75t_R g1390 ( .A(n_1391), .Y(n_1390) );
AOI31xp67_ASAP7_75t_SL g1392 ( .A1(n_1393), .A2(n_1395), .A3(n_1397), .B(n_1399), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVxp67_ASAP7_75t_SL g1397 ( .A(n_1398), .Y(n_1397) );
INVxp33_ASAP7_75t_L g1406 ( .A(n_1400), .Y(n_1406) );
BUFx3_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVxp67_ASAP7_75t_SL g1404 ( .A(n_1405), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
OAI21xp5_ASAP7_75t_L g1409 ( .A1(n_1410), .A2(n_1411), .B(n_1412), .Y(n_1409) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
endmodule