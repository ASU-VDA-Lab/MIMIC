module real_jpeg_32503_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_0),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_32),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_32),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_2),
.A2(n_32),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_71),
.B1(n_75),
.B2(n_80),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_80),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_5),
.A2(n_80),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_5),
.A2(n_80),
.B1(n_348),
.B2(n_350),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_6),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_15),
.B(n_18),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_53),
.B1(n_150),
.B2(n_154),
.Y(n_149)
);

AOI22x1_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_53),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_8),
.A2(n_53),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_8),
.B(n_417),
.Y(n_416)
);

OAI32xp33_ASAP7_75t_L g438 ( 
.A1(n_8),
.A2(n_439),
.A3(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_8),
.B(n_192),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_11),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_11),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_11),
.A2(n_267),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_L g399 ( 
.A1(n_11),
.A2(n_267),
.B1(n_400),
.B2(n_403),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_11),
.A2(n_267),
.B1(n_460),
.B2(n_462),
.Y(n_459)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_302),
.B(n_535),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_300),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_277),
.B(n_293),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_237),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_SL g304 ( 
.A(n_23),
.B(n_294),
.C(n_296),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_183),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_24),
.B(n_183),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_158),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_67),
.B1(n_156),
.B2(n_157),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_68),
.C(n_120),
.Y(n_67)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_26),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_26),
.A2(n_156),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_26),
.B(n_158),
.C(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_49),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_27),
.A2(n_174),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_27),
.B(n_263),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_28),
.B(n_57),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_34),
.Y(n_176)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_38),
.B(n_50),
.Y(n_262)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OA21x2_ASAP7_75t_SL g173 ( 
.A1(n_39),
.A2(n_174),
.B(n_181),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_SL g356 ( 
.A(n_39),
.B(n_53),
.Y(n_356)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2x1p5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_40),
.A2(n_50),
.B(n_57),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_40),
.B(n_264),
.Y(n_315)
);

AO22x2_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_45),
.Y(n_340)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_47),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_49),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_54),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_55),
.Y(n_54)
);

AOI32xp33_ASAP7_75t_L g410 ( 
.A1(n_53),
.A2(n_411),
.A3(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_53),
.B(n_440),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_R g479 ( 
.A(n_53),
.B(n_137),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_53),
.B(n_213),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_54),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_57),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_57),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_64),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_66),
.Y(n_332)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_69),
.B(n_121),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_81),
.B(n_109),
.Y(n_69)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g162 ( 
.A(n_82),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_82),
.B(n_320),
.Y(n_355)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_83),
.B(n_166),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_83),
.A2(n_166),
.B(n_287),
.Y(n_286)
);

AO21x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_99),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_85),
.Y(n_414)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_90),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_102),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_102),
.Y(n_402)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_106),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_109),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_110),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_112),
.Y(n_287)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_116),
.Y(n_329)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_121),
.B1(n_160),
.B2(n_172),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_120),
.A2(n_121),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_121),
.B(n_160),
.C(n_173),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_121),
.B(n_314),
.C(n_318),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_148),
.B(n_149),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_122),
.B(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_122),
.B(n_149),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_122),
.B(n_399),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_128),
.B1(n_131),
.B2(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_144),
.B2(n_147),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_140),
.Y(n_453)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

NAND2x1p5_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_148),
.B(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_148),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_195),
.Y(n_194)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_153),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_153),
.Y(n_413)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_157),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_173),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2x1p5_ASAP7_75t_L g318 ( 
.A(n_162),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_164),
.B(n_355),
.Y(n_376)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_170),
.Y(n_324)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_181),
.B(n_262),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_L g384 ( 
.A(n_182),
.B(n_315),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_205),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_189),
.A2(n_190),
.B(n_193),
.Y(n_272)
);

NAND2x1_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_192),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_194),
.B(n_431),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_196),
.B(n_243),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_196),
.B(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_208),
.B(n_235),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_206),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_223),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_207),
.A2(n_208),
.B1(n_236),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_207),
.A2(n_208),
.B1(n_410),
.B2(n_421),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_207),
.A2(n_208),
.B1(n_223),
.B2(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_208),
.B(n_410),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B(n_218),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_211),
.A2(n_347),
.B(n_361),
.Y(n_369)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_212),
.B(n_219),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_212),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_214),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_216),
.Y(n_349)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_216),
.Y(n_462)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_217),
.Y(n_461)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_217),
.Y(n_487)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_246),
.Y(n_245)
);

BUFx4f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_223),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_233),
.B(n_234),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_234),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_234),
.B(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_235),
.B(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_236),
.A2(n_298),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_238),
.B(n_240),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_271),
.C(n_273),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_241),
.B(n_531),
.Y(n_530)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_257),
.C(n_260),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_242),
.B(n_521),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_SL g387 ( 
.A(n_244),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

AND2x4_ASAP7_75t_SL g457 ( 
.A(n_245),
.B(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_250),
.A2(n_343),
.B(n_347),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_250),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_251),
.B(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_258),
.B(n_261),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_259),
.Y(n_407)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2x1_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_272),
.B(n_274),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_294),
.B(n_296),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_291),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_291),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_288),
.C(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g515 ( 
.A(n_285),
.B(n_384),
.C(n_385),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_286),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_299),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_298),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_506),
.B(n_532),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_392),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_377),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_364),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_312),
.B(n_365),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_325),
.C(n_352),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_313),
.B(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_319),
.B(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2x2_ASAP7_75t_L g502 ( 
.A(n_325),
.B(n_353),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_342),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_326),
.B(n_342),
.Y(n_373)
);

OAI31xp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.A3(n_333),
.B(n_334),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_338),
.B(n_341),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.C(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_426),
.Y(n_428)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_359),
.Y(n_483)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_361),
.B(n_458),
.Y(n_480)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_372),
.C(n_391),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_370),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_371),
.B(n_398),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_375),
.C(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_390),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g507 ( 
.A1(n_378),
.A2(n_390),
.B(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_378),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_379),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_386),
.B1(n_387),
.B2(n_389),
.Y(n_381)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_382),
.Y(n_512)
);

XOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_386),
.B(n_511),
.C(n_513),
.Y(n_510)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_390),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_500),
.B(n_504),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_433),
.B(n_499),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_422),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_395),
.B(n_422),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_406),
.C(n_408),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g497 ( 
.A(n_397),
.B(n_406),
.Y(n_497)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_409),
.B(n_497),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_423),
.B(n_430),
.C(n_432),
.Y(n_503)
);

OAI22x1_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_424),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_492),
.B(n_498),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_468),
.B(n_491),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_456),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_456),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_454),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_437),
.A2(n_438),
.B1(n_454),
.B2(n_455),
.Y(n_470)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_463),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_457),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_464),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_465),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_465),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_494),
.C(n_495),
.Y(n_493)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_477),
.B(n_490),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_471),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_483),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21x1_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_481),
.B(n_489),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_480),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_488),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_496),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_503),
.Y(n_505)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_509),
.C(n_524),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_514),
.B1(n_522),
.B2(n_523),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_514),
.Y(n_534)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_518),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_520),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_524),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_530),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_530),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.C(n_528),
.Y(n_525)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule