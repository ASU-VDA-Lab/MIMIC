module fake_jpeg_16094_n_18 (n_3, n_2, n_1, n_0, n_4, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_2),
.Y(n_5)
);

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_5),
.A2(n_4),
.B1(n_0),
.B2(n_3),
.Y(n_11)
);

NOR3xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_12),
.C(n_13),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_4),
.B(n_6),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_6),
.C(n_7),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_12),
.C(n_15),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_15),
.B(n_12),
.Y(n_18)
);


endmodule