module real_aes_1037_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_784, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_784;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_0), .B(n_132), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_1), .A2(n_141), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_2), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_3), .B(n_132), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_4), .B(n_148), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_5), .B(n_148), .Y(n_211) );
INVx1_ASAP7_75t_L g139 ( .A(n_6), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_7), .B(n_148), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_8), .Y(n_778) );
NAND2xp33_ASAP7_75t_L g149 ( .A(n_9), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g467 ( .A(n_10), .B(n_158), .Y(n_467) );
AND2x2_ASAP7_75t_L g527 ( .A(n_11), .B(n_127), .Y(n_527) );
INVx2_ASAP7_75t_L g129 ( .A(n_12), .Y(n_129) );
AOI221x1_ASAP7_75t_L g227 ( .A1(n_13), .A2(n_25), .B1(n_132), .B2(n_141), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_14), .B(n_148), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_15), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_16), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_17), .B(n_132), .Y(n_131) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_18), .A2(n_127), .B(n_130), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_19), .B(n_166), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_20), .B(n_148), .Y(n_175) );
AO21x1_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_132), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_22), .B(n_132), .Y(n_532) );
INVx1_ASAP7_75t_L g113 ( .A(n_23), .Y(n_113) );
NOR2xp33_ASAP7_75t_SL g775 ( .A(n_23), .B(n_114), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_24), .A2(n_87), .B1(n_132), .B2(n_472), .Y(n_471) );
NAND2x1_ASAP7_75t_L g197 ( .A(n_26), .B(n_148), .Y(n_197) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_27), .B(n_150), .Y(n_185) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_28), .A2(n_84), .B(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g153 ( .A(n_28), .B(n_84), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_29), .B(n_150), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_30), .B(n_148), .Y(n_147) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_31), .A2(n_158), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_32), .B(n_150), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_33), .A2(n_141), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_34), .B(n_148), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_35), .A2(n_141), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g138 ( .A(n_36), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g142 ( .A(n_36), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g480 ( .A(n_36), .Y(n_480) );
OR2x6_ASAP7_75t_L g111 ( .A(n_37), .B(n_112), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_37), .B(n_777), .C(n_779), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_38), .B(n_132), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_39), .B(n_132), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_40), .B(n_148), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_41), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_42), .B(n_150), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_43), .B(n_132), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_44), .A2(n_141), .B(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_45), .A2(n_141), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_46), .B(n_150), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_47), .B(n_150), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_48), .B(n_132), .Y(n_498) );
INVx1_ASAP7_75t_L g135 ( .A(n_49), .Y(n_135) );
INVx1_ASAP7_75t_L g145 ( .A(n_49), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_50), .B(n_148), .Y(n_465) );
AND2x2_ASAP7_75t_L g487 ( .A(n_51), .B(n_166), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_52), .B(n_150), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_53), .B(n_148), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_54), .B(n_150), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_55), .A2(n_141), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_56), .B(n_132), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_57), .B(n_132), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_58), .A2(n_141), .B(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_59), .Y(n_753) );
AO21x1_ASAP7_75t_L g208 ( .A1(n_60), .A2(n_141), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g538 ( .A(n_61), .B(n_167), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_62), .B(n_132), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_64), .B(n_150), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_65), .B(n_132), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_66), .B(n_150), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_67), .A2(n_91), .B1(n_141), .B2(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g221 ( .A(n_68), .B(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_69), .B(n_148), .Y(n_535) );
INVx1_ASAP7_75t_L g137 ( .A(n_70), .Y(n_137) );
INVx1_ASAP7_75t_L g143 ( .A(n_70), .Y(n_143) );
AND2x2_ASAP7_75t_L g189 ( .A(n_71), .B(n_158), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_72), .B(n_150), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_73), .A2(n_141), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_74), .A2(n_141), .B(n_455), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_75), .A2(n_141), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g510 ( .A(n_76), .B(n_167), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_77), .A2(n_445), .B1(n_446), .B2(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_77), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_78), .B(n_166), .Y(n_469) );
INVx1_ASAP7_75t_L g114 ( .A(n_79), .Y(n_114) );
AND2x2_ASAP7_75t_L g157 ( .A(n_80), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_81), .B(n_132), .Y(n_177) );
AND2x2_ASAP7_75t_L g458 ( .A(n_82), .B(n_127), .Y(n_458) );
AND2x2_ASAP7_75t_L g207 ( .A(n_83), .B(n_152), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_85), .B(n_150), .Y(n_176) );
AND2x2_ASAP7_75t_L g201 ( .A(n_86), .B(n_158), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_88), .B(n_148), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_89), .A2(n_141), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_90), .B(n_150), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_92), .A2(n_141), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_93), .B(n_148), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_94), .B(n_148), .Y(n_164) );
BUFx2_ASAP7_75t_L g537 ( .A(n_95), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_96), .Y(n_759) );
BUFx2_ASAP7_75t_L g104 ( .A(n_97), .Y(n_104) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_97), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_98), .A2(n_141), .B(n_146), .Y(n_140) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_772), .B(n_780), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_116), .B(n_763), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_106), .A2(n_768), .B(n_770), .Y(n_767) );
NOR2xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_115), .Y(n_106) );
INVx1_ASAP7_75t_SL g771 ( .A(n_107), .Y(n_771) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OR2x6_ASAP7_75t_SL g444 ( .A(n_109), .B(n_110), .Y(n_444) );
AND2x6_ASAP7_75t_SL g752 ( .A(n_109), .B(n_111), .Y(n_752) );
OR2x2_ASAP7_75t_L g762 ( .A(n_109), .B(n_111), .Y(n_762) );
CKINVDCx16_ASAP7_75t_R g779 ( .A(n_109), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_753), .B(n_754), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_442), .B1(n_445), .B2(n_749), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_120), .A2(n_446), .B1(n_756), .B2(n_757), .Y(n_755) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_363), .Y(n_120) );
NOR3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_275), .C(n_315), .Y(n_121) );
OAI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_190), .B1(n_239), .B2(n_254), .C(n_257), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_154), .Y(n_124) );
INVx2_ASAP7_75t_L g272 ( .A(n_125), .Y(n_272) );
AND2x2_ASAP7_75t_L g302 ( .A(n_125), .B(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g240 ( .A(n_126), .B(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g247 ( .A(n_126), .B(n_180), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_126), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_126), .B(n_156), .Y(n_262) );
INVx1_ASAP7_75t_L g278 ( .A(n_126), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_126), .B(n_324), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_127), .A2(n_532), .B(n_533), .Y(n_531) );
BUFx4f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
AND2x4_ASAP7_75t_L g152 ( .A(n_129), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_129), .B(n_153), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_140), .B(n_152), .Y(n_130) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_138), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
AND2x6_ASAP7_75t_L g150 ( .A(n_134), .B(n_143), .Y(n_150) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g148 ( .A(n_136), .B(n_145), .Y(n_148) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx5_ASAP7_75t_L g151 ( .A(n_138), .Y(n_151) );
AND2x2_ASAP7_75t_L g144 ( .A(n_139), .B(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_139), .Y(n_475) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx3_ASAP7_75t_L g476 ( .A(n_142), .Y(n_476) );
INVx2_ASAP7_75t_L g482 ( .A(n_143), .Y(n_482) );
AND2x4_ASAP7_75t_L g478 ( .A(n_144), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g474 ( .A(n_145), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_151), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_150), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_151), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_151), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_151), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_151), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_151), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_151), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_151), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_151), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_151), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_151), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_151), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_151), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_151), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_151), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_SL g171 ( .A(n_152), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_152), .B(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_152), .A2(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_168), .Y(n_154) );
INVx4_ASAP7_75t_L g243 ( .A(n_155), .Y(n_243) );
AND2x2_ASAP7_75t_L g274 ( .A(n_155), .B(n_181), .Y(n_274) );
AND2x2_ASAP7_75t_L g350 ( .A(n_155), .B(n_324), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_155), .B(n_180), .Y(n_392) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_156), .B(n_180), .Y(n_279) );
AND2x2_ASAP7_75t_L g303 ( .A(n_156), .B(n_181), .Y(n_303) );
BUFx2_ASAP7_75t_L g319 ( .A(n_156), .Y(n_319) );
NOR2x1_ASAP7_75t_SL g422 ( .A(n_156), .B(n_324), .Y(n_422) );
OR2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_160), .Y(n_156) );
INVx3_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_159), .A2(n_461), .B(n_467), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_166), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_166), .Y(n_188) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_166), .A2(n_227), .B(n_231), .Y(n_226) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_166), .A2(n_227), .B(n_231), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_166), .A2(n_453), .B(n_454), .Y(n_452) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_166), .A2(n_471), .B(n_477), .Y(n_470) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g299 ( .A(n_168), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_168), .A2(n_366), .B1(n_368), .B2(n_370), .C(n_375), .Y(n_365) );
AND2x2_ASAP7_75t_L g385 ( .A(n_168), .B(n_278), .Y(n_385) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_180), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g241 ( .A(n_170), .Y(n_241) );
INVx1_ASAP7_75t_L g294 ( .A(n_170), .Y(n_294) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_178), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_171), .B(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_171), .A2(n_172), .B(n_178), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_180), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g263 ( .A(n_180), .B(n_251), .Y(n_263) );
INVx2_ASAP7_75t_L g305 ( .A(n_180), .Y(n_305) );
AND2x2_ASAP7_75t_L g438 ( .A(n_180), .B(n_253), .Y(n_438) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_181), .Y(n_295) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_188), .B(n_189), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
AOI21x1_ASAP7_75t_L g520 ( .A1(n_188), .A2(n_521), .B(n_527), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_222), .C(n_237), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
INVx2_ASAP7_75t_L g352 ( .A(n_192), .Y(n_352) );
AND2x2_ASAP7_75t_L g397 ( .A(n_192), .B(n_274), .Y(n_397) );
BUFx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g342 ( .A(n_193), .Y(n_342) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_193), .B(n_269), .Y(n_357) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_200), .B(n_201), .Y(n_193) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_194), .A2(n_200), .B(n_201), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_199), .Y(n_194) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_200), .A2(n_215), .B(n_221), .Y(n_214) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_200), .A2(n_215), .B(n_221), .Y(n_234) );
AO21x1_ASAP7_75t_SL g503 ( .A1(n_200), .A2(n_504), .B(n_510), .Y(n_503) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_200), .A2(n_504), .B(n_510), .Y(n_561) );
INVx2_ASAP7_75t_L g311 ( .A(n_202), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_202), .B(n_341), .Y(n_367) );
AND2x4_ASAP7_75t_L g400 ( .A(n_202), .B(n_347), .Y(n_400) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_214), .Y(n_202) );
AND2x2_ASAP7_75t_L g238 ( .A(n_203), .B(n_233), .Y(n_238) );
OR2x2_ASAP7_75t_L g268 ( .A(n_203), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_203), .B(n_289), .Y(n_337) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g256 ( .A(n_205), .Y(n_256) );
OAI21x1_ASAP7_75t_SL g205 ( .A1(n_206), .A2(n_208), .B(n_212), .Y(n_205) );
INVx1_ASAP7_75t_L g213 ( .A(n_207), .Y(n_213) );
INVx2_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_216), .B(n_220), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_222), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_232), .Y(n_223) );
AND2x2_ASAP7_75t_L g237 ( .A(n_224), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g310 ( .A(n_224), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g395 ( .A(n_224), .Y(n_395) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g255 ( .A(n_225), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g374 ( .A(n_225), .B(n_234), .Y(n_374) );
AND2x2_ASAP7_75t_L g378 ( .A(n_225), .B(n_244), .Y(n_378) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g347 ( .A(n_226), .Y(n_347) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_226), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_232), .B(n_255), .Y(n_331) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_233), .B(n_256), .Y(n_441) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g245 ( .A(n_234), .B(n_236), .Y(n_245) );
AND2x2_ASAP7_75t_L g327 ( .A(n_234), .B(n_289), .Y(n_327) );
AND2x2_ASAP7_75t_L g346 ( .A(n_234), .B(n_235), .Y(n_346) );
BUFx2_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_235), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g244 ( .A(n_236), .Y(n_244) );
INVxp67_ASAP7_75t_L g287 ( .A(n_236), .Y(n_287) );
INVx1_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
AND2x2_ASAP7_75t_L g296 ( .A(n_238), .B(n_267), .Y(n_296) );
NAND2xp33_ASAP7_75t_L g377 ( .A(n_238), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g414 ( .A(n_238), .B(n_415), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_242), .B1(n_245), .B2(n_246), .C(n_248), .Y(n_239) );
AND2x2_ASAP7_75t_L g343 ( .A(n_240), .B(n_243), .Y(n_343) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_240), .B(n_303), .Y(n_362) );
AND2x2_ASAP7_75t_L g380 ( .A(n_240), .B(n_305), .Y(n_380) );
AND2x2_ASAP7_75t_L g435 ( .A(n_240), .B(n_274), .Y(n_435) );
INVx1_ASAP7_75t_L g251 ( .A(n_241), .Y(n_251) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_242), .Y(n_387) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_243), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_243), .B(n_294), .Y(n_369) );
AND2x2_ASAP7_75t_L g336 ( .A(n_244), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g372 ( .A(n_244), .Y(n_372) );
AND2x2_ASAP7_75t_L g281 ( .A(n_245), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_245), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g423 ( .A(n_245), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_245), .B(n_347), .Y(n_433) );
AND2x4_ASAP7_75t_L g349 ( .A(n_246), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g420 ( .A(n_247), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
OR2x2_ASAP7_75t_L g291 ( .A(n_252), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g298 ( .A(n_253), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g329 ( .A(n_253), .B(n_303), .Y(n_329) );
AND2x2_ASAP7_75t_L g403 ( .A(n_253), .B(n_324), .Y(n_403) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g351 ( .A(n_255), .B(n_352), .Y(n_351) );
OAI32xp33_ASAP7_75t_L g416 ( .A1(n_255), .A2(n_417), .A3(n_419), .B1(n_420), .B2(n_423), .Y(n_416) );
AND2x4_ASAP7_75t_L g288 ( .A(n_256), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g386 ( .A(n_256), .B(n_289), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B1(n_264), .B2(n_270), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g375 ( .A1(n_259), .A2(n_273), .B(n_376), .C(n_377), .Y(n_375) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g359 ( .A(n_260), .B(n_287), .Y(n_359) );
INVx1_ASAP7_75t_SL g430 ( .A(n_261), .Y(n_430) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x4_ASAP7_75t_L g333 ( .A(n_263), .B(n_272), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_263), .A2(n_412), .B1(n_413), .B2(n_414), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_268), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_271), .A2(n_301), .B1(n_354), .B2(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_272), .A2(n_390), .B(n_398), .C(n_411), .Y(n_389) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g309 ( .A(n_274), .B(n_278), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_280), .B(n_283), .C(n_312), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g426 ( .A(n_278), .B(n_422), .Y(n_426) );
OAI32xp33_ASAP7_75t_L g383 ( .A1(n_279), .A2(n_384), .A3(n_386), .B1(n_387), .B2(n_388), .Y(n_383) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_282), .B(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_290), .B1(n_296), .B2(n_297), .C(n_300), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g440 ( .A(n_287), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_288), .B(n_352), .Y(n_354) );
A2O1A1O1Ixp25_ASAP7_75t_L g425 ( .A1(n_288), .A2(n_357), .B(n_373), .C(n_419), .D(n_426), .Y(n_425) );
AOI31xp33_ASAP7_75t_L g427 ( .A1(n_288), .A2(n_309), .A3(n_419), .B(n_426), .Y(n_427) );
AND2x2_ASAP7_75t_L g341 ( .A(n_289), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_291), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx2_ASAP7_75t_L g418 ( .A(n_293), .Y(n_418) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g413 ( .A(n_294), .B(n_305), .Y(n_413) );
INVx1_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
AND2x2_ASAP7_75t_L g313 ( .A(n_297), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AOI31xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .A3(n_308), .B(n_310), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_303), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g436 ( .A(n_303), .B(n_382), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g381 ( .A(n_305), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g407 ( .A(n_305), .Y(n_407) );
INVxp67_ASAP7_75t_L g376 ( .A(n_306), .Y(n_376) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g314 ( .A(n_310), .Y(n_314) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_332), .C(n_348), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_325), .B1(n_329), .B2(n_330), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g402 ( .A(n_319), .Y(n_402) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_323), .Y(n_382) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_323), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_323), .B(n_392), .Y(n_409) );
NAND2xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B1(n_343), .B2(n_344), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_335), .B(n_338), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_346), .B1(n_380), .B2(n_381), .C(n_383), .Y(n_379) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g419 ( .A(n_346), .Y(n_419) );
AND2x2_ASAP7_75t_L g356 ( .A(n_347), .B(n_357), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_SL g404 ( .A1(n_347), .A2(n_405), .B(n_409), .C(n_410), .Y(n_404) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_353), .C(n_358), .Y(n_348) );
AND2x2_ASAP7_75t_L g399 ( .A(n_352), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
AOI21xp33_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_360), .B(n_361), .Y(n_358) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_389), .C(n_424), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_379), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
INVxp67_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g396 ( .A(n_386), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_396), .B2(n_397), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_404), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g437 ( .A(n_422), .B(n_438), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B1(n_428), .B2(n_431), .C(n_434), .Y(n_424) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI31xp33_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .A3(n_437), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx4f_ASAP7_75t_SL g756 ( .A(n_442), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx11_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_SL g446 ( .A(n_447), .B(n_645), .Y(n_446) );
NOR3xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_554), .C(n_586), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_483), .B1(n_511), .B2(n_528), .C(n_539), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_459), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g517 ( .A(n_451), .B(n_460), .Y(n_517) );
INVx4_ASAP7_75t_L g545 ( .A(n_451), .Y(n_545) );
AND2x4_ASAP7_75t_SL g585 ( .A(n_451), .B(n_519), .Y(n_585) );
BUFx2_ASAP7_75t_L g595 ( .A(n_451), .Y(n_595) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_451), .B(n_600), .Y(n_661) );
AND2x2_ASAP7_75t_L g670 ( .A(n_451), .B(n_598), .Y(n_670) );
OR2x2_ASAP7_75t_L g678 ( .A(n_451), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g704 ( .A(n_451), .B(n_543), .Y(n_704) );
AND2x4_ASAP7_75t_L g723 ( .A(n_451), .B(n_724), .Y(n_723) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_458), .Y(n_451) );
INVx2_ASAP7_75t_SL g636 ( .A(n_459), .Y(n_636) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_468), .Y(n_459) );
AND2x2_ASAP7_75t_L g543 ( .A(n_460), .B(n_520), .Y(n_543) );
INVx2_ASAP7_75t_L g570 ( .A(n_460), .Y(n_570) );
INVx2_ASAP7_75t_L g600 ( .A(n_460), .Y(n_600) );
AND2x2_ASAP7_75t_L g614 ( .A(n_460), .B(n_519), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
AND2x2_ASAP7_75t_L g544 ( .A(n_468), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g567 ( .A(n_468), .Y(n_567) );
BUFx3_ASAP7_75t_L g581 ( .A(n_468), .Y(n_581) );
AND2x2_ASAP7_75t_L g610 ( .A(n_468), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
AND2x4_ASAP7_75t_L g515 ( .A(n_469), .B(n_470), .Y(n_515) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR2x1p5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g616 ( .A(n_483), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_494), .Y(n_483) );
OR2x2_ASAP7_75t_L g727 ( .A(n_484), .B(n_528), .Y(n_727) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g583 ( .A(n_485), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_485), .B(n_494), .Y(n_644) );
OR2x2_ASAP7_75t_L g742 ( .A(n_485), .B(n_664), .Y(n_742) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_529), .Y(n_553) );
OR2x2_ASAP7_75t_SL g563 ( .A(n_486), .B(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_486), .Y(n_625) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_486), .B(n_530), .Y(n_631) );
AND2x2_ASAP7_75t_L g656 ( .A(n_486), .B(n_496), .Y(n_656) );
OR2x2_ASAP7_75t_L g677 ( .A(n_486), .B(n_560), .Y(n_677) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g572 ( .A(n_494), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_494), .A2(n_666), .B(n_669), .C(n_671), .Y(n_665) );
AND2x2_ASAP7_75t_L g738 ( .A(n_494), .B(n_514), .Y(n_738) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx1_ASAP7_75t_L g605 ( .A(n_495), .Y(n_605) );
AND2x2_ASAP7_75t_L g675 ( .A(n_495), .B(n_530), .Y(n_675) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g549 ( .A(n_496), .Y(n_549) );
OR2x2_ASAP7_75t_L g564 ( .A(n_496), .B(n_530), .Y(n_564) );
INVx1_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
AND2x2_ASAP7_75t_L g592 ( .A(n_496), .B(n_503), .Y(n_592) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_496), .Y(n_698) );
NOR2x1_ASAP7_75t_SL g529 ( .A(n_503), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
OR2x2_ASAP7_75t_L g662 ( .A(n_513), .B(n_597), .Y(n_662) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_514), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g744 ( .A(n_514), .B(n_641), .Y(n_744) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g589 ( .A(n_515), .B(n_570), .Y(n_589) );
AND2x2_ASAP7_75t_L g685 ( .A(n_515), .B(n_598), .Y(n_685) );
INVx1_ASAP7_75t_L g602 ( .A(n_516), .Y(n_602) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g652 ( .A(n_517), .Y(n_652) );
INVx2_ASAP7_75t_L g619 ( .A(n_518), .Y(n_619) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g569 ( .A(n_519), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g599 ( .A(n_519), .Y(n_599) );
INVx1_ASAP7_75t_L g724 ( .A(n_519), .Y(n_724) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_520), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
OR2x2_ASAP7_75t_L g695 ( .A(n_528), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g550 ( .A(n_530), .Y(n_550) );
OR2x2_ASAP7_75t_L g573 ( .A(n_530), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g584 ( .A(n_530), .B(n_560), .Y(n_584) );
AND2x2_ASAP7_75t_L g658 ( .A(n_530), .B(n_574), .Y(n_658) );
BUFx2_ASAP7_75t_L g741 ( .A(n_530), .Y(n_741) );
OR2x6_ASAP7_75t_L g530 ( .A(n_531), .B(n_538), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_546), .B(n_551), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x2_ASAP7_75t_L g693 ( .A(n_542), .B(n_615), .Y(n_693) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g552 ( .A(n_543), .B(n_545), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_544), .B(n_614), .Y(n_715) );
INVx1_ASAP7_75t_L g745 ( .A(n_544), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_545), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_545), .B(n_681), .Y(n_718) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_548), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_548), .B(n_576), .Y(n_729) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_549), .B(n_631), .Y(n_687) );
AND2x2_ASAP7_75t_L g705 ( .A(n_549), .B(n_658), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_550), .B(n_592), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_550), .A2(n_596), .B(n_638), .C(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_552), .A2(n_625), .B1(n_733), .B2(n_739), .C(n_743), .Y(n_732) );
INVx1_ASAP7_75t_SL g720 ( .A(n_553), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_565), .B1(n_571), .B2(n_575), .C(n_784), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g630 ( .A(n_559), .Y(n_630) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g604 ( .A(n_560), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g635 ( .A(n_560), .B(n_580), .Y(n_635) );
INVx2_ASAP7_75t_L g668 ( .A(n_560), .Y(n_668) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI32xp33_ASAP7_75t_L g719 ( .A1(n_563), .A2(n_610), .A3(n_641), .B1(n_720), .B2(n_721), .Y(n_719) );
OR2x2_ASAP7_75t_L g690 ( .A(n_564), .B(n_677), .Y(n_690) );
INVx1_ASAP7_75t_L g700 ( .A(n_565), .Y(n_700) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx2_ASAP7_75t_L g615 ( .A(n_566), .Y(n_615) );
AND2x2_ASAP7_75t_L g686 ( .A(n_566), .B(n_661), .Y(n_686) );
OR2x2_ASAP7_75t_L g717 ( .A(n_566), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_567), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g611 ( .A(n_570), .Y(n_611) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_SL g576 ( .A(n_573), .Y(n_576) );
OR2x2_ASAP7_75t_L g663 ( .A(n_573), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_574), .B(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_574), .B(n_698), .Y(n_697) );
BUFx2_ASAP7_75t_L g710 ( .A(n_574), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_582), .C(n_585), .Y(n_575) );
AND2x2_ASAP7_75t_L g725 ( .A(n_577), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g651 ( .A(n_581), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_581), .B(n_585), .Y(n_672) );
AND2x2_ASAP7_75t_L g703 ( .A(n_581), .B(n_704), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_583), .A2(n_714), .B(n_716), .C(n_719), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_584), .A2(n_588), .B1(n_590), .B2(n_593), .C1(n_601), .C2(n_603), .Y(n_587) );
AND2x2_ASAP7_75t_L g655 ( .A(n_584), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g588 ( .A(n_585), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g609 ( .A(n_585), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g586 ( .A(n_587), .B(n_606), .C(n_627), .D(n_637), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_589), .B(n_595), .Y(n_649) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g657 ( .A(n_592), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g664 ( .A(n_592), .Y(n_664) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_594), .A2(n_628), .B(n_632), .C(n_636), .Y(n_627) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_595), .B(n_610), .Y(n_731) );
OR2x2_ASAP7_75t_L g735 ( .A(n_595), .B(n_621), .Y(n_735) );
INVx1_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_SL g642 ( .A(n_599), .Y(n_642) );
INVx1_ASAP7_75t_L g622 ( .A(n_600), .Y(n_622) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_602), .B(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g626 ( .A(n_604), .Y(n_626) );
AOI322xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .A3(n_610), .B1(n_612), .B2(n_616), .C1(n_617), .C2(n_623), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_SL g688 ( .A1(n_609), .A2(n_689), .B(n_690), .C(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g711 ( .A(n_610), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g669 ( .A(n_615), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_621), .Y(n_691) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx3_ASAP7_75t_L g634 ( .A(n_631), .Y(n_634) );
OR2x2_ASAP7_75t_L g702 ( .A(n_631), .B(n_664), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_631), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_SL g734 ( .A(n_635), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_636), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND3xp33_ASAP7_75t_SL g739 ( .A(n_644), .B(n_740), .C(n_742), .Y(n_739) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_683), .C(n_712), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_665), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B(n_653), .C(n_659), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g692 ( .A1(n_648), .A2(n_670), .A3(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx2_ASAP7_75t_L g707 ( .A(n_655), .Y(n_707) );
INVx1_ASAP7_75t_L g682 ( .A(n_657), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g709 ( .A(n_667), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g748 ( .A(n_668), .Y(n_748) );
OAI22xp33_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_673), .B1(n_678), .B2(n_682), .Y(n_671) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_677), .Y(n_689) );
OR2x2_ASAP7_75t_L g740 ( .A(n_677), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_692), .C(n_699), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B(n_687), .C(n_688), .Y(n_684) );
INVx2_ASAP7_75t_L g721 ( .A(n_685), .Y(n_721) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_709), .B2(n_711), .Y(n_706) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_722), .C(n_732), .Y(n_712) );
INVxp33_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_725), .B1(n_728), .B2(n_730), .Y(n_722) );
INVx2_ASAP7_75t_L g736 ( .A(n_723), .Y(n_736) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp33_ASAP7_75t_SL g743 ( .A1(n_742), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx6p67_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx4_ASAP7_75t_SL g757 ( .A(n_750), .Y(n_757) );
INVx3_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_755), .B(n_758), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g782 ( .A(n_773), .Y(n_782) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x4_ASAP7_75t_SL g774 ( .A(n_775), .B(n_776), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
endmodule