module fake_jpeg_26974_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_58),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_47),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_77),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_54),
.Y(n_96)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_51),
.B1(n_45),
.B2(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_70),
.B1(n_88),
.B2(n_83),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_60),
.B1(n_55),
.B2(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_92),
.B1(n_50),
.B2(n_49),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_59),
.B(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_52),
.B1(n_43),
.B2(n_25),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_102),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_53),
.B1(n_81),
.B2(n_56),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_106),
.B1(n_97),
.B2(n_83),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_89),
.B(n_95),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_111),
.B(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_113),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_91),
.B(n_84),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_23),
.B(n_39),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_22),
.B1(n_38),
.B2(n_37),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_19),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_31),
.C(n_10),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_121),
.Y(n_130)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_106),
.B1(n_3),
.B2(n_5),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_122),
.B(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_0),
.B(n_5),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_126),
.B1(n_9),
.B2(n_12),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_107),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_8),
.B(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_8),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_125),
.B1(n_15),
.B2(n_16),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_118),
.C(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_128),
.B1(n_130),
.B2(n_129),
.Y(n_136)
);

OAI221xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_130),
.B1(n_127),
.B2(n_27),
.C(n_32),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_137),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_13),
.B(n_21),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_33),
.Y(n_143)
);


endmodule