module fake_ariane_3110_n_1209 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1209);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1209;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_1118;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_1187;
wire n_985;
wire n_421;
wire n_245;
wire n_1167;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_443;
wire n_586;
wire n_286;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_515;
wire n_379;
wire n_445;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_1067;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_1018;
wire n_597;
wire n_269;
wire n_816;
wire n_784;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1201;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_271;
wire n_1153;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_478;
wire n_222;
wire n_703;
wire n_1207;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_957;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_705;
wire n_658;
wire n_630;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_262;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_741;
wire n_371;
wire n_845;
wire n_1135;
wire n_199;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_217;
wire n_673;
wire n_1114;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_249;
wire n_1108;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_851;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_785;
wire n_669;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_608;
wire n_959;
wire n_494;
wire n_892;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_33),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_177),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_54),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_89),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_55),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_147),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_41),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_36),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_141),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_72),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_105),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_100),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_13),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_131),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_96),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_107),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_51),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_90),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_29),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_124),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_171),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_93),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_94),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_67),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_13),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_82),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_73),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_88),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_120),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_87),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_130),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_81),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_159),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_156),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_15),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_74),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_180),
.Y(n_274)
);

BUFx2_ASAP7_75t_SL g275 ( 
.A(n_117),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_163),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_115),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_28),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_37),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_139),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_132),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_16),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_168),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_1),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_40),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_153),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_64),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_95),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_2),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_270),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_184),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_194),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_202),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_199),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_211),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_272),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_188),
.B(n_0),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_279),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_219),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_229),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_232),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_191),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_239),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_207),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_240),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_251),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_187),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_301),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_259),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_280),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_212),
.B(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_221),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_223),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_182),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_182),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_215),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_2),
.Y(n_349)
);

INVx4_ASAP7_75t_R g350 ( 
.A(n_216),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_215),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_254),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_216),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_246),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_3),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_295),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_181),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_185),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_254),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g363 ( 
.A(n_230),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_186),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_252),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_192),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_196),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_253),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_264),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_256),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_197),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_198),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_263),
.B(n_3),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_266),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_296),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_224),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_200),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_284),
.B(n_4),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_224),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_285),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_284),
.B(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_293),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_205),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_206),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_360),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_361),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_305),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_365),
.B(n_190),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_190),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_298),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_298),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_363),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_242),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_238),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_242),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_383),
.B(n_193),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_193),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_310),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_309),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_312),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_323),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_225),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_303),
.B(n_275),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_363),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_311),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_313),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_380),
.B(n_208),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_314),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_315),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_316),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_382),
.B(n_193),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_307),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_320),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_324),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_318),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_373),
.B(n_209),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_375),
.B(n_210),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_383),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_350),
.B(n_193),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_391),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_321),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_328),
.B(n_195),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_338),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_325),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_327),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_330),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_332),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_344),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_308),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_302),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_195),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_319),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_412),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_456),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_336),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_308),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_326),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_444),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_410),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_335),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_401),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_462),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_411),
.B(n_384),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_339),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_384),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_343),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_410),
.B(n_348),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_446),
.B(n_358),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_335),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

CKINVDCx6p67_ASAP7_75t_R g507 ( 
.A(n_452),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_437),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_451),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_435),
.B(n_374),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_461),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_431),
.B(n_344),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_449),
.A2(n_189),
.B1(n_377),
.B2(n_370),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_435),
.B(n_347),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_411),
.B(n_5),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_347),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_458),
.B(n_213),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_429),
.B(n_418),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

NOR2x1p5_ASAP7_75t_L g528 ( 
.A(n_398),
.B(n_351),
.Y(n_528)
);

INVx4_ASAP7_75t_SL g529 ( 
.A(n_451),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_458),
.B(n_214),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_515),
.A2(n_448),
.B1(n_379),
.B2(n_370),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_521),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_472),
.B(n_450),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_513),
.B(n_480),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_493),
.B(n_450),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_476),
.B(n_458),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_493),
.B(n_450),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_475),
.B(n_455),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_481),
.B(n_424),
.Y(n_546)
);

AO22x2_ASAP7_75t_L g547 ( 
.A1(n_487),
.A2(n_492),
.B1(n_514),
.B2(n_448),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_490),
.B(n_443),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_483),
.B(n_458),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_487),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_497),
.B(n_455),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_487),
.A2(n_353),
.B1(n_379),
.B2(n_377),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_501),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_502),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_452),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_L g562 ( 
.A1(n_463),
.A2(n_500),
.B(n_499),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_511),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_504),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_504),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_505),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_469),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_505),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_526),
.B(n_452),
.Y(n_569)
);

OAI221xp5_ASAP7_75t_L g570 ( 
.A1(n_469),
.A2(n_417),
.B1(n_409),
.B2(n_453),
.C(n_439),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_526),
.B(n_478),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_465),
.B(n_455),
.Y(n_572)
);

OAI221xp5_ASAP7_75t_L g573 ( 
.A1(n_512),
.A2(n_417),
.B1(n_409),
.B2(n_453),
.C(n_439),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_511),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_525),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_518),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_478),
.B(n_459),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_459),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

AO22x2_ASAP7_75t_L g583 ( 
.A1(n_492),
.A2(n_351),
.B1(n_362),
.B2(n_353),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

OAI221xp5_ASAP7_75t_L g585 ( 
.A1(n_512),
.A2(n_453),
.B1(n_439),
.B2(n_436),
.C(n_433),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_471),
.Y(n_586)
);

AO22x2_ASAP7_75t_L g587 ( 
.A1(n_492),
.A2(n_362),
.B1(n_306),
.B2(n_317),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_473),
.Y(n_589)
);

BUFx8_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_473),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_465),
.B(n_455),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_532),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_465),
.B(n_459),
.Y(n_596)
);

AO22x2_ASAP7_75t_L g597 ( 
.A1(n_519),
.A2(n_522),
.B1(n_520),
.B2(n_317),
.Y(n_597)
);

AO22x2_ASAP7_75t_L g598 ( 
.A1(n_519),
.A2(n_304),
.B1(n_306),
.B2(n_322),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_532),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_522),
.A2(n_304),
.B1(n_322),
.B2(n_404),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_520),
.A2(n_405),
.B1(n_404),
.B2(n_418),
.Y(n_602)
);

OAI221xp5_ASAP7_75t_L g603 ( 
.A1(n_491),
.A2(n_396),
.B1(n_400),
.B2(n_408),
.C(n_414),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_507),
.B(n_402),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_507),
.B(n_402),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_520),
.B(n_428),
.C(n_427),
.Y(n_609)
);

AO22x2_ASAP7_75t_L g610 ( 
.A1(n_528),
.A2(n_405),
.B1(n_404),
.B2(n_418),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_474),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_467),
.B(n_418),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_529),
.B(n_405),
.Y(n_613)
);

OAI221xp5_ASAP7_75t_L g614 ( 
.A1(n_524),
.A2(n_393),
.B1(n_400),
.B2(n_414),
.C(n_415),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_467),
.B(n_412),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_485),
.A2(n_429),
.B1(n_454),
.B2(n_422),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_479),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_486),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

NAND2x1_ASAP7_75t_L g621 ( 
.A(n_468),
.B(n_440),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_498),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_498),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_530),
.A2(n_429),
.B1(n_454),
.B2(n_428),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_508),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_506),
.B(n_427),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_506),
.A2(n_429),
.B1(n_454),
.B2(n_403),
.Y(n_627)
);

AO22x2_ASAP7_75t_L g628 ( 
.A1(n_506),
.A2(n_454),
.B1(n_421),
.B2(n_393),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_580),
.B(n_470),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_580),
.B(n_470),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_529),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_581),
.B(n_470),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_581),
.B(n_412),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_560),
.B(n_412),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_560),
.B(n_412),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_544),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_569),
.B(n_412),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_569),
.B(n_468),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_536),
.B(n_445),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_572),
.B(n_447),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_571),
.B(n_468),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_567),
.B(n_509),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_562),
.B(n_545),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_541),
.B(n_509),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_SL g645 ( 
.A(n_593),
.B(n_434),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_543),
.B(n_509),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_SL g647 ( 
.A(n_596),
.B(n_434),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_552),
.B(n_467),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_535),
.B(n_466),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_613),
.B(n_466),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_613),
.B(n_466),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_607),
.B(n_466),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_608),
.B(n_626),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_542),
.B(n_440),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_609),
.B(n_477),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_549),
.B(n_546),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_557),
.B(n_477),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_551),
.B(n_534),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_534),
.B(n_488),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_561),
.B(n_488),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_602),
.B(n_467),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_606),
.B(n_503),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_590),
.B(n_503),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_590),
.B(n_510),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_621),
.B(n_440),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g666 ( 
.A(n_550),
.B(n_440),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_SL g667 ( 
.A(n_556),
.B(n_394),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_612),
.B(n_510),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_537),
.B(n_527),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_537),
.B(n_527),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_558),
.B(n_396),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_588),
.B(n_531),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_588),
.B(n_531),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_SL g674 ( 
.A(n_559),
.B(n_564),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_589),
.B(n_437),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_597),
.B(n_415),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_589),
.B(n_437),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_591),
.B(n_437),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_554),
.B(n_419),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_565),
.B(n_419),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_591),
.B(n_508),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_594),
.B(n_421),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_SL g683 ( 
.A(n_566),
.B(n_568),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_594),
.B(n_425),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_625),
.B(n_529),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_620),
.B(n_425),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_620),
.B(n_508),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_597),
.B(n_432),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_622),
.B(n_516),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_622),
.B(n_516),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_576),
.B(n_577),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_623),
.B(n_516),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_623),
.B(n_529),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_625),
.B(n_579),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_584),
.B(n_416),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_595),
.B(n_416),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_599),
.B(n_416),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_582),
.B(n_420),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_SL g699 ( 
.A(n_548),
.B(n_420),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_586),
.B(n_420),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_611),
.B(n_438),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_617),
.B(n_438),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_618),
.B(n_432),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_619),
.B(n_441),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_600),
.B(n_441),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_615),
.B(n_441),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_538),
.B(n_401),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_602),
.B(n_467),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_539),
.B(n_217),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_540),
.B(n_218),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_467),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_604),
.B(n_220),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_605),
.B(n_222),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_563),
.B(n_227),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_574),
.B(n_231),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_601),
.B(n_6),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_575),
.B(n_235),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_578),
.B(n_553),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_555),
.B(n_236),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_627),
.B(n_244),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_573),
.B(n_423),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_627),
.B(n_628),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_628),
.B(n_250),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_639),
.A2(n_585),
.B(n_614),
.C(n_603),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_682),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_643),
.A2(n_273),
.B(n_258),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_636),
.B(n_616),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_676),
.B(n_600),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_691),
.A2(n_624),
.B(n_610),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_649),
.A2(n_616),
.B(n_110),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_698),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_666),
.A2(n_271),
.B(n_257),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_700),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_653),
.B(n_547),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_688),
.B(n_705),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_681),
.A2(n_108),
.B(n_160),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_656),
.B(n_547),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_631),
.B(n_195),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_684),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_644),
.A2(n_260),
.B(n_261),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_704),
.A2(n_274),
.B(n_262),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_716),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_631),
.B(n_195),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_681),
.A2(n_102),
.B(n_142),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_SL g745 ( 
.A1(n_716),
.A2(n_533),
.B(n_598),
.Y(n_745)
);

AOI221x1_ASAP7_75t_L g746 ( 
.A1(n_720),
.A2(n_683),
.B1(n_674),
.B2(n_708),
.C(n_661),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_685),
.B(n_204),
.Y(n_747)
);

AOI221x1_ASAP7_75t_L g748 ( 
.A1(n_667),
.A2(n_533),
.B1(n_598),
.B2(n_583),
.C(n_554),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_652),
.B(n_583),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_686),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_646),
.A2(n_265),
.B(n_267),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_658),
.B(n_268),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_716),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_633),
.B(n_587),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_695),
.Y(n_755)
);

OAI21x1_ASAP7_75t_SL g756 ( 
.A1(n_648),
.A2(n_6),
.B(n_7),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

AO32x2_ASAP7_75t_L g758 ( 
.A1(n_722),
.A2(n_587),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_758)
);

AOI31xp67_ASAP7_75t_L g759 ( 
.A1(n_675),
.A2(n_677),
.A3(n_678),
.B(n_706),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_634),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_645),
.A2(n_297),
.B(n_292),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_696),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_647),
.A2(n_289),
.B(n_286),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_640),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_671),
.A2(n_281),
.B(n_276),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_697),
.A2(n_269),
.B(n_8),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_641),
.B(n_7),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_680),
.A2(n_249),
.B(n_234),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_635),
.B(n_637),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_721),
.A2(n_249),
.B(n_234),
.C(n_226),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_654),
.A2(n_249),
.B(n_234),
.C(n_226),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_679),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_694),
.A2(n_79),
.B(n_179),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_650),
.Y(n_774)
);

AO31x2_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_249),
.A3(n_226),
.B(n_204),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_629),
.B(n_10),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_642),
.A2(n_226),
.B(n_204),
.Y(n_777)
);

OA21x2_ASAP7_75t_L g778 ( 
.A1(n_703),
.A2(n_75),
.B(n_169),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_630),
.B(n_11),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_687),
.A2(n_11),
.B(n_12),
.C(n_15),
.Y(n_780)
);

AOI221x1_ASAP7_75t_L g781 ( 
.A1(n_699),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_781)
);

AO21x2_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_80),
.B(n_167),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_632),
.B(n_17),
.Y(n_783)
);

AO31x2_ASAP7_75t_L g784 ( 
.A1(n_718),
.A2(n_83),
.A3(n_165),
.B(n_161),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_665),
.A2(n_70),
.B(n_158),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_689),
.A2(n_63),
.B(n_157),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_SL g787 ( 
.A1(n_772),
.A2(n_663),
.B1(n_664),
.B2(n_659),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_767),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_764),
.B(n_657),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_730),
.A2(n_693),
.B(n_692),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_757),
.B(n_651),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_729),
.B(n_655),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_753),
.B(n_660),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_754),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_777),
.A2(n_690),
.B(n_673),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_713),
.B1(n_712),
.B2(n_710),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_785),
.A2(n_669),
.B(n_670),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_757),
.B(n_758),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_773),
.A2(n_672),
.B(n_702),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_736),
.A2(n_701),
.B(n_668),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_744),
.A2(n_746),
.B(n_768),
.Y(n_802)
);

CKINVDCx6p67_ASAP7_75t_R g803 ( 
.A(n_742),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_767),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_726),
.A2(n_709),
.B1(n_717),
.B2(n_715),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_757),
.B(n_707),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_SL g807 ( 
.A(n_766),
.B(n_714),
.C(n_719),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_776),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_757),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_728),
.A2(n_662),
.B1(n_638),
.B2(n_22),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_726),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_778),
.A2(n_78),
.B(n_152),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_778),
.A2(n_62),
.B(n_150),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_725),
.B(n_61),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_747),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_733),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_779),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_756),
.A2(n_60),
.B(n_149),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_742),
.B(n_745),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_747),
.Y(n_820)
);

OA21x2_ASAP7_75t_L g821 ( 
.A1(n_770),
.A2(n_58),
.B(n_144),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_739),
.B(n_750),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_738),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_727),
.B(n_20),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_737),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_781),
.B(n_21),
.C(n_23),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_752),
.B(n_84),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_745),
.B(n_23),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_749),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_760),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_734),
.B(n_24),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_755),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_760),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_786),
.A2(n_86),
.B(n_136),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_762),
.B(n_85),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_759),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_766),
.A2(n_25),
.B(n_26),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_738),
.A2(n_57),
.B(n_134),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_769),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_740),
.B(n_25),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_735),
.B(n_774),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_840),
.A2(n_783),
.B(n_780),
.C(n_740),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_836),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_832),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_790),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_832),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_839),
.B(n_748),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_830),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_797),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_816),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_840),
.A2(n_751),
.B(n_761),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_816),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_833),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_841),
.B(n_775),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_788),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_790),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_841),
.B(n_775),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_804),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_825),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_799),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_828),
.A2(n_782),
.B1(n_758),
.B2(n_751),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_802),
.A2(n_771),
.B(n_775),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_822),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_799),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_822),
.B(n_758),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_792),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_792),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_812),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_809),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_801),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_801),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_800),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_837),
.A2(n_782),
.B(n_763),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_800),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_817),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_814),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_809),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_812),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_818),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_838),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_838),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_795),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_824),
.B(n_743),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_809),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_795),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_815),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_824),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_835),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_815),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_830),
.B(n_831),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_869),
.B(n_814),
.Y(n_898)
);

CKINVDCx11_ASAP7_75t_R g899 ( 
.A(n_865),
.Y(n_899)
);

XNOR2xp5_ASAP7_75t_L g900 ( 
.A(n_849),
.B(n_787),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_894),
.B(n_794),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_R g902 ( 
.A(n_869),
.B(n_807),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_856),
.B(n_859),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_856),
.B(n_829),
.Y(n_904)
);

BUFx10_ASAP7_75t_L g905 ( 
.A(n_879),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_860),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_863),
.B(n_789),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_865),
.B(n_881),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_881),
.B(n_809),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_897),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_R g911 ( 
.A(n_867),
.B(n_835),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_R g912 ( 
.A(n_867),
.B(n_835),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_860),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_871),
.B(n_895),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_871),
.B(n_823),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_854),
.B(n_861),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_895),
.B(n_890),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_871),
.B(n_823),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_893),
.B(n_823),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_873),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_873),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_880),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_883),
.B(n_803),
.Y(n_923)
);

XNOR2xp5_ASAP7_75t_L g924 ( 
.A(n_861),
.B(n_811),
.Y(n_924)
);

BUFx10_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_859),
.B(n_789),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_862),
.B(n_819),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_R g929 ( 
.A(n_848),
.B(n_821),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_893),
.B(n_820),
.Y(n_930)
);

CKINVDCx11_ASAP7_75t_R g931 ( 
.A(n_845),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_R g932 ( 
.A(n_893),
.B(n_821),
.Y(n_932)
);

XNOR2xp5_ASAP7_75t_L g933 ( 
.A(n_866),
.B(n_827),
.Y(n_933)
);

XNOR2xp5_ASAP7_75t_L g934 ( 
.A(n_866),
.B(n_796),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_845),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_868),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_914),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_SL g938 ( 
.A(n_910),
.B(n_852),
.C(n_842),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_926),
.B(n_868),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_844),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_SL g941 ( 
.A1(n_898),
.A2(n_877),
.B1(n_826),
.B2(n_805),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_903),
.B(n_870),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_903),
.B(n_855),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_920),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_905),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_935),
.B(n_855),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_906),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_914),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_908),
.B(n_844),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_898),
.B(n_870),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_913),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_927),
.Y(n_952)
);

OAI221xp5_ASAP7_75t_L g953 ( 
.A1(n_902),
.A2(n_810),
.B1(n_882),
.B2(n_885),
.C(n_793),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_905),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_898),
.B(n_909),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_907),
.B(n_843),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_927),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_904),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_904),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_909),
.B(n_843),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_917),
.B(n_858),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_934),
.B(n_858),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_901),
.B(n_874),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_921),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_931),
.B(n_874),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_919),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_929),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_921),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_924),
.B(n_875),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_928),
.A2(n_852),
.B1(n_877),
.B2(n_853),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_919),
.B(n_915),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_921),
.B(n_875),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_915),
.B(n_847),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_918),
.B(n_876),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_967),
.B(n_918),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_947),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_959),
.B(n_847),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_952),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_L g979 ( 
.A1(n_967),
.A2(n_911),
.B1(n_912),
.B2(n_932),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_952),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_944),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_959),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_941),
.A2(n_900),
.B1(n_933),
.B2(n_885),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_957),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_958),
.B(n_930),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_947),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_938),
.A2(n_899),
.B1(n_877),
.B2(n_806),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_951),
.Y(n_988)
);

NAND2x1_ASAP7_75t_L g989 ( 
.A(n_937),
.B(n_948),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_937),
.B(n_846),
.Y(n_990)
);

AO21x2_ASAP7_75t_L g991 ( 
.A1(n_938),
.A2(n_882),
.B(n_886),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_951),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_956),
.Y(n_993)
);

AOI31xp33_ASAP7_75t_L g994 ( 
.A1(n_941),
.A2(n_886),
.A3(n_887),
.B(n_923),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_957),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_948),
.B(n_846),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_955),
.B(n_846),
.Y(n_997)
);

BUFx12f_ASAP7_75t_L g998 ( 
.A(n_954),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_958),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_978),
.B(n_958),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_975),
.B(n_982),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_975),
.B(n_965),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_984),
.B(n_969),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_984),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_945),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_995),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_978),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_975),
.B(n_965),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_995),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_975),
.B(n_955),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_989),
.B(n_969),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_989),
.B(n_974),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_981),
.B(n_955),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_980),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_976),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_980),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_999),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_999),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_993),
.B(n_963),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1003),
.B(n_940),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_R g1022 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1008),
.B(n_940),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_1004),
.B(n_945),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1000),
.B(n_1015),
.Y(n_1025)
);

AO221x2_ASAP7_75t_L g1026 ( 
.A1(n_1004),
.A2(n_983),
.B1(n_1015),
.B2(n_1017),
.C(n_979),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_1004),
.Y(n_1027)
);

AO221x2_ASAP7_75t_L g1028 ( 
.A1(n_1017),
.A2(n_994),
.B1(n_962),
.B2(n_981),
.C(n_954),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1000),
.B(n_977),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_1006),
.B(n_954),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_R g1031 ( 
.A(n_1012),
.B(n_962),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1028),
.B(n_1002),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_1027),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_1030),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1026),
.A2(n_994),
.B1(n_987),
.B2(n_1011),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_1031),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1028),
.B(n_1002),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1025),
.B(n_1011),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1033),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1033),
.B(n_1029),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1034),
.B(n_1023),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_1036),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1042),
.B(n_1038),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1041),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1039),
.B(n_1038),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1039),
.B(n_1032),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1040),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1040),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1042),
.B(n_1038),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_1038),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_1042),
.B(n_1035),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1045),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_1048),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1048),
.Y(n_1056)
);

INVxp33_ASAP7_75t_SL g1057 ( 
.A(n_1044),
.Y(n_1057)
);

INVxp33_ASAP7_75t_SL g1058 ( 
.A(n_1051),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_1052),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1043),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_1047),
.Y(n_1061)
);

INVx6_ASAP7_75t_L g1062 ( 
.A(n_1046),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1049),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1050),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1045),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1045),
.B(n_1032),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_1048),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1045),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1059),
.B(n_1037),
.Y(n_1070)
);

AOI211xp5_ASAP7_75t_L g1071 ( 
.A1(n_1065),
.A2(n_1037),
.B(n_1024),
.C(n_953),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1058),
.A2(n_1009),
.B1(n_1011),
.B2(n_1014),
.Y(n_1072)
);

NAND5xp2_ASAP7_75t_L g1073 ( 
.A(n_1058),
.B(n_1009),
.C(n_1022),
.D(n_1001),
.E(n_987),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1057),
.B(n_1010),
.Y(n_1074)
);

NAND4xp25_ASAP7_75t_L g1075 ( 
.A(n_1068),
.B(n_1001),
.C(n_1013),
.D(n_1014),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1061),
.B(n_953),
.C(n_1010),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1059),
.B(n_1021),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1059),
.B(n_1011),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_SL g1079 ( 
.A1(n_1068),
.A2(n_1014),
.B(n_1013),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1059),
.B(n_1010),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1056),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_L g1082 ( 
.A(n_1056),
.B(n_1005),
.Y(n_1082)
);

AO21x1_ASAP7_75t_L g1083 ( 
.A1(n_1063),
.A2(n_1005),
.B(n_1007),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_L g1084 ( 
.A(n_1063),
.B(n_1007),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1055),
.A2(n_991),
.B(n_1019),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1062),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1067),
.A2(n_991),
.B(n_1019),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1081),
.Y(n_1088)
);

AOI221xp5_ASAP7_75t_L g1089 ( 
.A1(n_1076),
.A2(n_1069),
.B1(n_1066),
.B2(n_1054),
.C(n_1060),
.Y(n_1089)
);

AOI222xp33_ASAP7_75t_L g1090 ( 
.A1(n_1070),
.A2(n_1086),
.B1(n_1064),
.B2(n_1080),
.C1(n_1074),
.C2(n_1077),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1082),
.B(n_1062),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_1084),
.B(n_1062),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1071),
.A2(n_991),
.B1(n_970),
.B2(n_1018),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_1018),
.B1(n_765),
.B2(n_1016),
.C(n_936),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1078),
.B(n_990),
.Y(n_1095)
);

AOI211xp5_ASAP7_75t_L g1096 ( 
.A1(n_1083),
.A2(n_963),
.B(n_996),
.C(n_990),
.Y(n_1096)
);

OAI211xp5_ASAP7_75t_SL g1097 ( 
.A1(n_1087),
.A2(n_1079),
.B(n_1085),
.C(n_1072),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1075),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1086),
.B(n_1020),
.C(n_936),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1086),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1081),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1076),
.A2(n_1016),
.B1(n_964),
.B2(n_968),
.Y(n_1102)
);

AOI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1070),
.A2(n_1016),
.B1(n_992),
.B2(n_988),
.C1(n_986),
.C2(n_976),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1081),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1088),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_981),
.Y(n_1106)
);

AND4x1_ASAP7_75t_L g1107 ( 
.A(n_1090),
.B(n_732),
.C(n_30),
.D(n_31),
.Y(n_1107)
);

NAND4xp75_ASAP7_75t_L g1108 ( 
.A(n_1092),
.B(n_821),
.C(n_803),
.D(n_964),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1093),
.A2(n_968),
.B1(n_1020),
.B2(n_997),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1101),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1089),
.B(n_939),
.C(n_741),
.Y(n_1111)
);

XNOR2xp5_ASAP7_75t_L g1112 ( 
.A(n_1098),
.B(n_26),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1100),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1091),
.B(n_31),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1102),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1095),
.Y(n_1116)
);

NAND4xp75_ASAP7_75t_L g1117 ( 
.A(n_1094),
.B(n_939),
.C(n_985),
.D(n_973),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_L g1118 ( 
.A(n_1097),
.B(n_32),
.Y(n_1118)
);

AO22x1_ASAP7_75t_L g1119 ( 
.A1(n_1103),
.A2(n_981),
.B1(n_944),
.B2(n_997),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1099),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_1096),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_SL g1122 ( 
.A(n_1091),
.B(n_981),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1093),
.A2(n_997),
.B1(n_950),
.B2(n_974),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_1104),
.B(n_32),
.Y(n_1124)
);

XNOR2xp5_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_34),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1104),
.B(n_996),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1088),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1088),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1114),
.B(n_35),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_1105),
.B(n_1110),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_1105),
.B(n_35),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1118),
.B(n_981),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_SL g1133 ( 
.A(n_1128),
.B(n_944),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_1112),
.B(n_37),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1116),
.B(n_944),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1107),
.B(n_38),
.C(n_39),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_R g1137 ( 
.A(n_1125),
.B(n_39),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1113),
.B(n_942),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1127),
.B(n_42),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1124),
.B(n_942),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1106),
.B(n_806),
.C(n_972),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_SL g1142 ( 
.A(n_1106),
.B(n_997),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_1126),
.B(n_43),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_L g1144 ( 
.A(n_1120),
.B(n_972),
.C(n_973),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1121),
.B(n_971),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1111),
.B(n_950),
.C(n_820),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1115),
.B(n_950),
.C(n_820),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1117),
.B(n_950),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1122),
.B(n_986),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1109),
.B(n_971),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_R g1151 ( 
.A(n_1108),
.B(n_44),
.Y(n_1151)
);

OAI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1132),
.A2(n_1123),
.B1(n_1119),
.B2(n_988),
.C(n_992),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_SL g1153 ( 
.A(n_1133),
.B(n_798),
.C(n_961),
.Y(n_1153)
);

OR3x1_ASAP7_75t_L g1154 ( 
.A(n_1136),
.B(n_887),
.C(n_878),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1129),
.B(n_993),
.Y(n_1155)
);

AND3x1_ASAP7_75t_L g1156 ( 
.A(n_1130),
.B(n_966),
.C(n_891),
.Y(n_1156)
);

NOR2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1138),
.B(n_1140),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1151),
.A2(n_943),
.B1(n_930),
.B2(n_961),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1135),
.A2(n_834),
.B(n_971),
.Y(n_1159)
);

NAND4xp75_ASAP7_75t_L g1160 ( 
.A(n_1145),
.B(n_891),
.C(n_949),
.D(n_864),
.Y(n_1160)
);

XOR2xp5_ASAP7_75t_L g1161 ( 
.A(n_1137),
.B(n_943),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1131),
.B(n_971),
.Y(n_1162)
);

OAI222xp33_ASAP7_75t_L g1163 ( 
.A1(n_1148),
.A2(n_955),
.B1(n_946),
.B2(n_966),
.C1(n_791),
.C2(n_876),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1134),
.B(n_1143),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1149),
.Y(n_1165)
);

OA22x2_ASAP7_75t_L g1166 ( 
.A1(n_1150),
.A2(n_966),
.B1(n_892),
.B2(n_888),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1141),
.A2(n_946),
.B1(n_846),
.B2(n_857),
.Y(n_1167)
);

XNOR2x1_ASAP7_75t_L g1168 ( 
.A(n_1139),
.B(n_813),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1144),
.A2(n_857),
.B1(n_878),
.B2(n_888),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1146),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1147),
.Y(n_1171)
);

CKINVDCx11_ASAP7_75t_R g1172 ( 
.A(n_1165),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_1142),
.C(n_820),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1161),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1162),
.A2(n_1170),
.B(n_1153),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1157),
.Y(n_1176)
);

OR5x1_ASAP7_75t_L g1177 ( 
.A(n_1154),
.B(n_920),
.C(n_925),
.D(n_50),
.E(n_52),
.Y(n_1177)
);

AOI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1171),
.A2(n_872),
.B1(n_889),
.B2(n_884),
.C(n_857),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1157),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1159),
.A2(n_834),
.B(n_892),
.Y(n_1180)
);

NAND4xp25_ASAP7_75t_L g1181 ( 
.A(n_1155),
.B(n_857),
.C(n_949),
.D(n_960),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1168),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1176),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_1179),
.A2(n_1160),
.B1(n_1167),
.B2(n_1169),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1177),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1172),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1174),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1182),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1175),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1173),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1180),
.B(n_1156),
.Y(n_1191)
);

AOI31xp33_ASAP7_75t_L g1192 ( 
.A1(n_1186),
.A2(n_1152),
.A3(n_1158),
.B(n_1178),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1188),
.A2(n_1166),
.B1(n_1181),
.B2(n_1163),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1190),
.A2(n_884),
.B1(n_872),
.B2(n_889),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1191),
.A2(n_872),
.B1(n_889),
.B2(n_864),
.Y(n_1195)
);

AOI31xp33_ASAP7_75t_L g1196 ( 
.A1(n_1189),
.A2(n_1183),
.A3(n_1187),
.B(n_1185),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1183),
.A2(n_864),
.B1(n_853),
.B2(n_850),
.Y(n_1197)
);

AOI31xp33_ASAP7_75t_L g1198 ( 
.A1(n_1184),
.A2(n_791),
.A3(n_47),
.B(n_53),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1184),
.A2(n_864),
.B1(n_850),
.B2(n_851),
.Y(n_1199)
);

NOR5xp2_ASAP7_75t_L g1200 ( 
.A(n_1196),
.B(n_45),
.C(n_56),
.D(n_101),
.E(n_103),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1193),
.A2(n_896),
.B1(n_893),
.B2(n_815),
.Y(n_1201)
);

NAND4xp25_ASAP7_75t_L g1202 ( 
.A(n_1199),
.B(n_104),
.C(n_106),
.D(n_109),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1192),
.Y(n_1203)
);

AO22x1_ASAP7_75t_L g1204 ( 
.A1(n_1198),
.A2(n_815),
.B1(n_784),
.B2(n_896),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1203),
.A2(n_1195),
.B(n_1194),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1202),
.A2(n_1197),
.B1(n_851),
.B2(n_956),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1205),
.Y(n_1207)
);

OAI221xp5_ASAP7_75t_R g1208 ( 
.A1(n_1207),
.A2(n_1201),
.B1(n_1200),
.B2(n_1206),
.C(n_1204),
.Y(n_1208)
);

AOI211xp5_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_111),
.B(n_114),
.C(n_116),
.Y(n_1209)
);


endmodule