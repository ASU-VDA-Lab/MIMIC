module real_jpeg_27428_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_0),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_0),
.B(n_182),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_3),
.A2(n_4),
.B1(n_33),
.B2(n_64),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_33),
.B1(n_68),
.B2(n_69),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_4),
.A2(n_5),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_65),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_45),
.Y(n_53)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.Y(n_173)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_9),
.A2(n_10),
.B(n_43),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_25),
.B1(n_68),
.B2(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_10),
.B(n_64),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_64),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_91),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_81),
.Y(n_177)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_129),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_128),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_110),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_16),
.B(n_110),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_87),
.B2(n_109),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_21),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_22),
.A2(n_27),
.B(n_35),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_22),
.B(n_35),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_25),
.A2(n_69),
.B(n_82),
.C(n_138),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_25),
.A2(n_39),
.B(n_43),
.C(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_25),
.B(n_37),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_25),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_26),
.B(n_197),
.Y(n_196)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx5_ASAP7_75t_SL g198 ( 
.A(n_27),
.Y(n_198)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_53),
.B(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_30),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_35),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_37),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_38),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_38),
.B(n_58),
.Y(n_163)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_43),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_46),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_47),
.B(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_59),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_54),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_54),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_56),
.B(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_57),
.B(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_58),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.C(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_70),
.Y(n_103)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_79),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_73),
.B(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_78),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_78),
.B(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_127),
.Y(n_153)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.C(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_102),
.B(n_107),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_115),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_111),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_114),
.B(n_115),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.C(n_123),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_116),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_225),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_221),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_208),
.B(n_220),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_166),
.B(n_207),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_149),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_135),
.B(n_149),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.C(n_145),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_140),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_160),
.B2(n_161),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_162),
.C(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_202),
.B(n_206),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_201),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_200),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_194),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.B1(n_214),
.B2(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_222)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);


endmodule