module fake_jpeg_23549_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_26),
.Y(n_34)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_19),
.B1(n_27),
.B2(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_27),
.B1(n_24),
.B2(n_62),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_46),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_19),
.B1(n_24),
.B2(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_64),
.B1(n_51),
.B2(n_61),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_28),
.B1(n_19),
.B2(n_24),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_48),
.B1(n_45),
.B2(n_38),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_0),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_11),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_28),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_99),
.B1(n_101),
.B2(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_61),
.B1(n_51),
.B2(n_69),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_46),
.C(n_52),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_61),
.B1(n_65),
.B2(n_27),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_109),
.B1(n_73),
.B2(n_62),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_65),
.B1(n_81),
.B2(n_59),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_55),
.B1(n_44),
.B2(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_67),
.B1(n_73),
.B2(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_116),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_129),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_125),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_83),
.Y(n_125)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_131),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_63),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_72),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_54),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_84),
.B1(n_74),
.B2(n_39),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_140),
.B1(n_105),
.B2(n_110),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_79),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_94),
.B(n_117),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_152),
.B(n_156),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_94),
.B(n_80),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_150),
.A2(n_160),
.B(n_13),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_29),
.B(n_15),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_116),
.B1(n_92),
.B2(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_163),
.B1(n_127),
.B2(n_122),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_164),
.B1(n_42),
.B2(n_60),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_29),
.B(n_21),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_97),
.C(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_132),
.C(n_130),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_80),
.B(n_9),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_97),
.B1(n_105),
.B2(n_42),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_76),
.B(n_29),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_42),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_60),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_181),
.C(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_178),
.B(n_186),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_137),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_193),
.B(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_139),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_187),
.B(n_20),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_153),
.B1(n_171),
.B2(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_156),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_71),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_152),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_75),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_162),
.B1(n_163),
.B2(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_25),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_20),
.CON(n_202),
.SN(n_202)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_207),
.B(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_193),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_178),
.B1(n_177),
.B2(n_186),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_149),
.B(n_169),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_166),
.C(n_147),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_207),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_171),
.B1(n_166),
.B2(n_147),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_221),
.B1(n_177),
.B2(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_148),
.A3(n_165),
.B1(n_17),
.B2(n_20),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_194),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_12),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_180),
.C(n_12),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_25),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_181),
.C(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_191),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

AO21x2_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_98),
.B(n_79),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_236),
.B(n_242),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_212),
.B(n_213),
.C(n_238),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_234),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_221),
.B1(n_222),
.B2(n_201),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_204),
.B1(n_221),
.B2(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_241),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_235),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_193),
.Y(n_235)
);

FAx1_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_180),
.CI(n_2),
.CON(n_236),
.SN(n_236)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_202),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_98),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_243),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_16),
.B(n_15),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_98),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_22),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_21),
.C(n_30),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_263),
.B1(n_266),
.B2(n_21),
.Y(n_278)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_259),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_221),
.B1(n_210),
.B2(n_224),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_221),
.B1(n_210),
.B2(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_214),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_236),
.B1(n_227),
.B2(n_240),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_205),
.B1(n_216),
.B2(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_234),
.C(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_274),
.C(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_245),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_257),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_239),
.B(n_31),
.C(n_16),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_278),
.B1(n_259),
.B2(n_17),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_263),
.C(n_254),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_12),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_10),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_20),
.B(n_17),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_30),
.C(n_23),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_31),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_266),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_30),
.C(n_23),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_283),
.C(n_15),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_23),
.C(n_21),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_288),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_262),
.Y(n_288)
);

FAx1_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_256),
.CI(n_260),
.CON(n_289),
.SN(n_289)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_10),
.B(n_2),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_11),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_11),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_10),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_275),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_297),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_1),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_296),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_270),
.B1(n_272),
.B2(n_23),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_15),
.C(n_16),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_16),
.C(n_2),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_1),
.B(n_2),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_318),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_319),
.B1(n_305),
.B2(n_299),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_318),
.A2(n_3),
.B(n_4),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_326),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_310),
.B1(n_309),
.B2(n_5),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_324),
.A3(n_321),
.B1(n_320),
.B2(n_322),
.C1(n_326),
.C2(n_7),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_328),
.B(n_329),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_310),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_3),
.C(n_4),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_6),
.Y(n_335)
);


endmodule