module real_jpeg_24308_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_29),
.B1(n_34),
.B2(n_62),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_1),
.A2(n_40),
.B1(n_44),
.B2(n_62),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_65),
.B1(n_71),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_2),
.A2(n_40),
.B1(n_44),
.B2(n_65),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_3),
.B(n_73),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_55),
.C(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_109),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_66),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_3),
.B(n_40),
.C(n_89),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_3),
.A2(n_39),
.B(n_203),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_7),
.A2(n_40),
.B1(n_44),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_8),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_40),
.B1(n_44),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_34),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_12),
.A2(n_40),
.B1(n_44),
.B2(n_70),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_40),
.B1(n_44),
.B2(n_94),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_40),
.B1(n_44),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_124)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_16),
.Y(n_157)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_16),
.A2(n_38),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_21),
.B(n_112),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_96),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_22),
.B(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_23),
.B(n_51),
.C(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_24),
.B(n_37),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_26),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_73)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_26),
.B(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_39),
.A2(n_41),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_39),
.A2(n_83),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_39),
.A2(n_43),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_39),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_39),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_40),
.A2(n_44),
.B1(n_89),
.B2(n_91),
.Y(n_92)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_44),
.B(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_47),
.A2(n_217),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_67),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_63),
.Y(n_51)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_52),
.A2(n_63),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_53),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_53),
.A2(n_137),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_55),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_55),
.B(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_66),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_103),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_69),
.A2(n_73),
.B1(n_78),
.B2(n_133),
.Y(n_132)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_105),
.B(n_111),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_80),
.B(n_96),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_85),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_86),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_86),
.A2(n_191),
.B(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_87),
.A2(n_125),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_93),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_92),
.A2(n_99),
.B(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_92),
.B(n_109),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_100),
.B(n_125),
.Y(n_191)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_110),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_109),
.B(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_128),
.B2(n_129),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_246),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_160),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_144),
.B(n_158),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_145),
.A2(n_146),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_149),
.B(n_150),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_240),
.B(n_245),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_192),
.B(n_239),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_181),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_163),
.B(n_181),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_174),
.C(n_178),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_164),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_167),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B(n_172),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_178),
.B1(n_179),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_233),
.B(n_238),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_213),
.B(n_232),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_207),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_207),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_231),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_244),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule