module fake_jpeg_25930_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_25),
.B1(n_33),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_25),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_33),
.B1(n_25),
.B2(n_24),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_70),
.Y(n_125)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_71),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_45),
.Y(n_127)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_95),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_67),
.B1(n_53),
.B2(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_33),
.B1(n_23),
.B2(n_24),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_85),
.B1(n_91),
.B2(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_43),
.B1(n_41),
.B2(n_47),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_47),
.B1(n_39),
.B2(n_36),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_92),
.B1(n_26),
.B2(n_35),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_23),
.B1(n_27),
.B2(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_39),
.B1(n_36),
.B2(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_99),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_36),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_26),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_45),
.C(n_46),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_45),
.C(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_32),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_19),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_131),
.C(n_127),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_74),
.B1(n_79),
.B2(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_121),
.B1(n_101),
.B2(n_83),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_92),
.B1(n_78),
.B2(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_46),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_80),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_35),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_136),
.A2(n_18),
.B1(n_52),
.B2(n_48),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_162),
.B1(n_108),
.B2(n_111),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_125),
.B1(n_113),
.B2(n_71),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_154),
.B1(n_156),
.B2(n_165),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.C(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_141),
.Y(n_197)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_129),
.B(n_122),
.C(n_127),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_151),
.B(n_142),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_103),
.C(n_118),
.Y(n_183)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_90),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_160),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_102),
.B1(n_82),
.B2(n_103),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_72),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_40),
.B(n_19),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_106),
.B(n_72),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_103),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_77),
.B1(n_103),
.B2(n_73),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_164),
.Y(n_189)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_107),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_184),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_111),
.B(n_124),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_168),
.A2(n_173),
.B(n_179),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_187),
.B1(n_163),
.B2(n_141),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_117),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_155),
.A3(n_144),
.B1(n_145),
.B2(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_112),
.A3(n_118),
.B1(n_119),
.B2(n_26),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_114),
.B1(n_119),
.B2(n_112),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_189),
.B(n_170),
.C(n_191),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_181),
.B(n_29),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_188),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_52),
.C(n_105),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_77),
.B1(n_114),
.B2(n_69),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_35),
.C(n_40),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_35),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_192),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_40),
.B(n_105),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_146),
.B(n_139),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_40),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_68),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_48),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_199),
.B1(n_0),
.B2(n_1),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_19),
.B1(n_28),
.B2(n_31),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_229),
.B1(n_206),
.B2(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_12),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_224),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_210),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_221),
.B(n_207),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_225),
.B(n_187),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_214),
.Y(n_241)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_94),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_172),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_227),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_31),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_228),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_68),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_68),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_14),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_12),
.B(n_10),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_29),
.B1(n_28),
.B2(n_14),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_0),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_169),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_194),
.B(n_168),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_250),
.B1(n_216),
.B2(n_226),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_177),
.B1(n_173),
.B2(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_183),
.C(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.C(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_186),
.C(n_198),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_255),
.B1(n_229),
.B2(n_205),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_180),
.C(n_199),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_244),
.B(n_214),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_169),
.C(n_176),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_219),
.C(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_252),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_263),
.C(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_216),
.B1(n_200),
.B2(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_213),
.C(n_215),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_213),
.C(n_211),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_275),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_225),
.C(n_207),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_205),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_207),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_273),
.B1(n_232),
.B2(n_253),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_3),
.C(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_3),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_277),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_292),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_236),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_290),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_234),
.B1(n_235),
.B2(n_247),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_286),
.B1(n_248),
.B2(n_231),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_235),
.B1(n_253),
.B2(n_255),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_237),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_237),
.C(n_233),
.Y(n_291)
);

BUFx12f_ASAP7_75t_SL g307 ( 
.A(n_291),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_3),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_254),
.B(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_301),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_275),
.B(n_254),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_248),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_304),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_231),
.B(n_263),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_282),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_306),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_261),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_3),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.C(n_4),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_4),
.B(n_5),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_292),
.C(n_294),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_283),
.B(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_280),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_300),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_280),
.B(n_294),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_303),
.B(n_296),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_5),
.B(n_6),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_5),
.B(n_6),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_328),
.B(n_310),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_311),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_297),
.B1(n_305),
.B2(n_7),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_320),
.B1(n_314),
.B2(n_9),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_6),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_333),
.B(n_326),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_332),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_323),
.C(n_316),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_325),
.C(n_8),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_9),
.B(n_7),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_7),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_8),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_8),
.B(n_328),
.Y(n_342)
);


endmodule