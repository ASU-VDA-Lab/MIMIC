module fake_aes_1980_n_43 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
NOR2xp67_ASAP7_75t_L g12 ( .A(n_8), .B(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_2), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_18), .Y(n_22) );
OR2x6_ASAP7_75t_L g23 ( .A(n_18), .B(n_0), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_15), .B(n_1), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_22), .B(n_13), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_22), .B(n_13), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_17), .B1(n_16), .B2(n_12), .Y(n_27) );
AO22x1_ASAP7_75t_L g28 ( .A1(n_24), .A2(n_16), .B1(n_14), .B2(n_5), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_23), .B1(n_21), .B2(n_20), .C(n_19), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI221xp5_ASAP7_75t_SL g31 ( .A1(n_25), .A2(n_21), .B1(n_20), .B2(n_19), .C(n_23), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_26), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_30), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
AOI21xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_29), .B(n_30), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_23), .B1(n_31), .B2(n_21), .Y(n_37) );
AND4x2_ASAP7_75t_L g38 ( .A(n_34), .B(n_4), .C(n_5), .D(n_6), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g39 ( .A(n_38), .B(n_20), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_37), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
OAI222xp33_ASAP7_75t_L g42 ( .A1(n_39), .A2(n_4), .B1(n_9), .B2(n_19), .C1(n_36), .C2(n_40), .Y(n_42) );
NAND3xp33_ASAP7_75t_L g43 ( .A(n_41), .B(n_19), .C(n_42), .Y(n_43) );
endmodule