module fake_jpeg_10131_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_55),
.B1(n_38),
.B2(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_38),
.B1(n_33),
.B2(n_39),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_77),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_73),
.B1(n_44),
.B2(n_53),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_38),
.A3(n_42),
.B1(n_26),
.B2(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_23),
.B(n_22),
.C(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_15),
.Y(n_103)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_27),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_62),
.B1(n_51),
.B2(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_92),
.B1(n_104),
.B2(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_36),
.B1(n_49),
.B2(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_103),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_71),
.B1(n_58),
.B2(n_32),
.Y(n_117)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_46),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_46),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_32),
.B1(n_49),
.B2(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_32),
.B1(n_16),
.B2(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_122),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_37),
.C(n_36),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_92),
.C(n_89),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_120),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_125),
.B1(n_99),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_104),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_18),
.B(n_22),
.C(n_23),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_129),
.B(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_58),
.B1(n_16),
.B2(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_29),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_91),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.C(n_137),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_141),
.B(n_142),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_92),
.C(n_91),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_92),
.B(n_101),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_139),
.B(n_149),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_101),
.B(n_103),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_85),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_106),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_115),
.B(n_126),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_145),
.B1(n_131),
.B2(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_120),
.B(n_108),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_36),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_36),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_113),
.C(n_108),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_31),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_36),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_110),
.B1(n_116),
.B2(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_161),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_29),
.B(n_28),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_166),
.B(n_16),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_126),
.B1(n_97),
.B2(n_76),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_165),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_28),
.B(n_16),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_149),
.B1(n_140),
.B2(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_31),
.C(n_12),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_144),
.A3(n_130),
.B1(n_136),
.B2(n_133),
.C1(n_150),
.C2(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_173),
.Y(n_193)
);

OA21x2_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_130),
.B(n_31),
.Y(n_170)
);

OA21x2_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_166),
.B(n_159),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_174),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_182),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_36),
.C(n_107),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_180),
.C(n_183),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_36),
.C(n_107),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_19),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_2),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_31),
.C(n_19),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_192),
.B(n_7),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_162),
.B1(n_164),
.B2(n_151),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_176),
.B1(n_180),
.B2(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_162),
.B1(n_160),
.B2(n_14),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_2),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_31),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_3),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_172),
.B(n_174),
.CI(n_183),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_195),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_189),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_13),
.C(n_4),
.Y(n_199)
);

OR2x6_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_186),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_3),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_192),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_194),
.B1(n_193),
.B2(n_186),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_191),
.B(n_9),
.C(n_10),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_202),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_196),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_199),
.B(n_195),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_211),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_208),
.B1(n_190),
.B2(n_10),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_208),
.B(n_8),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_8),
.B(n_9),
.C(n_216),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_224),
.B(n_218),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.Y(n_228)
);


endmodule