module fake_jpeg_30873_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

BUFx8_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_20),
.B(n_21),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_24),
.B1(n_15),
.B2(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_8),
.B1(n_14),
.B2(n_11),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_25),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_31),
.Y(n_35)
);

OAI221xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B1(n_30),
.B2(n_15),
.C(n_9),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_30),
.B(n_23),
.Y(n_36)
);

AOI21x1_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_26),
.B(n_5),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_1),
.B1(n_7),
.B2(n_36),
.Y(n_40)
);


endmodule