module fake_ariane_725_n_3783 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_363, n_720, n_354, n_41, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_733, n_500, n_665, n_59, n_336, n_731, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_738, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_711, n_453, n_734, n_74, n_491, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_718, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_3783);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_363;
input n_720;
input n_354;
input n_41;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_733;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_738;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_3783;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_3416;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_754;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_829;
wire n_1761;
wire n_1062;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2391;
wire n_2332;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_3739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_772;
wire n_1216;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_3698;
wire n_3716;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_3678;
wire n_762;
wire n_1468;
wire n_1661;
wire n_1253;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3624;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_3306;
wire n_2748;
wire n_2185;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_1376;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_1178;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_1623;
wire n_990;
wire n_3559;
wire n_1903;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3724;
wire n_1920;
wire n_2083;
wire n_815;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2898;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_3467;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3569;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_1162;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3035;
wire n_887;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3766;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1975;
wire n_1373;
wire n_742;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1714;
wire n_1044;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_3097;
wire n_3507;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_854;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_1784;
wire n_3110;
wire n_771;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_3753;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_3718;
wire n_756;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_3381;
wire n_3455;
wire n_807;
wire n_3736;
wire n_891;
wire n_3313;
wire n_1659;
wire n_885;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_3605;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_3769;
wire n_825;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3731;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_3255;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1065;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3241;
wire n_1584;
wire n_1157;
wire n_848;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_3106;
wire n_2977;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_3470;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_3521;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_761;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_758;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_2897;
wire n_816;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_2775;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2705;
wire n_2664;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3194;
wire n_3143;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_881;
wire n_1477;
wire n_1777;
wire n_1019;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_3094;
wire n_741;
wire n_1410;
wire n_2297;
wire n_939;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_1923;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_3763;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3593;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3293;
wire n_3361;
wire n_1683;
wire n_1229;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_2269;
wire n_1474;
wire n_937;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_3547;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g740 ( 
.A(n_299),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_227),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_647),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_491),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_721),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_648),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_691),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_325),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_62),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_201),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_564),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_527),
.Y(n_751)
);

CKINVDCx16_ASAP7_75t_R g752 ( 
.A(n_643),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_438),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_98),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_129),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_22),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_120),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_441),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_725),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_626),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_633),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_206),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_366),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_456),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_154),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_87),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_153),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_133),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_527),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_201),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_591),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_327),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_724),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_705),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_606),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_78),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_292),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_214),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_712),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_522),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_134),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_509),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_462),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_171),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_194),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_31),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_672),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_252),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_342),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_45),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_528),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_110),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_385),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_204),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_173),
.Y(n_795)
);

BUFx2_ASAP7_75t_SL g796 ( 
.A(n_428),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_566),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_503),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_200),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_419),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_707),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_163),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_184),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_710),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_306),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_690),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_695),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_616),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_513),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_539),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_337),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_356),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_130),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_145),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_736),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_114),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_435),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_216),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_727),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_7),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_602),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_87),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_362),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_67),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_168),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_739),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_526),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_352),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_682),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_127),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_339),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_450),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_423),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_395),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_220),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_187),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_498),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_149),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_63),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_222),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_342),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_194),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_362),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_681),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_145),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_536),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_733),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_450),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_245),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_518),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_284),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_78),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_698),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_323),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_90),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_716),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_504),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_457),
.Y(n_858)
);

CKINVDCx16_ASAP7_75t_R g859 ( 
.A(n_170),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_701),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_149),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_678),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_594),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_542),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_706),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_178),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_49),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_34),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_476),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_628),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_520),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_108),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_323),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_667),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_694),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_466),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_689),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_16),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_642),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_268),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_358),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_138),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_666),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_532),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_526),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_413),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_316),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_480),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_27),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_475),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_8),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_102),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_599),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_374),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_456),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_123),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_455),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_651),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_732),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_388),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_25),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_218),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_60),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_446),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_569),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_146),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_118),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_361),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_333),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_256),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_696),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_187),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_179),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_165),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_98),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_412),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_208),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_384),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_658),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_662),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_659),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_279),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_134),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_391),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_653),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_461),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_516),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_458),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_586),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_688),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_20),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_620),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_533),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_635),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_469),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_266),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_714),
.Y(n_937)
);

BUFx10_ASAP7_75t_L g938 ( 
.A(n_49),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_665),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_559),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_500),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_79),
.Y(n_942)
);

BUFx8_ASAP7_75t_SL g943 ( 
.A(n_541),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_346),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_311),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_107),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_304),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_216),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_660),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_205),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_624),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_649),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_95),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_141),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_118),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_108),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_93),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_452),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_249),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_622),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_40),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_738),
.Y(n_962)
);

BUFx8_ASAP7_75t_SL g963 ( 
.A(n_403),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_62),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_361),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_627),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_234),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_266),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_619),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_537),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_440),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_429),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_223),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_380),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_8),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_544),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_730),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_416),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_535),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_636),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_143),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_14),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_207),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_55),
.Y(n_984)
);

CKINVDCx16_ASAP7_75t_R g985 ( 
.A(n_287),
.Y(n_985)
);

BUFx10_ASAP7_75t_L g986 ( 
.A(n_341),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_522),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_369),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_231),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_543),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_422),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_406),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_109),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_652),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_717),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_123),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_141),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_107),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_597),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_472),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_467),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_669),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_541),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_337),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_488),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_646),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_175),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_260),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_211),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_483),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_15),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_325),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_377),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_75),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_630),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_679),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_428),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_197),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_155),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_242),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_548),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_202),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_645),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_354),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_99),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_608),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_369),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_184),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_507),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_562),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_719),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_6),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_663),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_60),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_155),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_54),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_576),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_700),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_621),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_708),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_718),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_685),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_692),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_321),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_366),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_629),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_693),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_80),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_442),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_113),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_77),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_510),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_684),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_499),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_11),
.Y(n_1055)
);

CKINVDCx14_ASAP7_75t_R g1056 ( 
.A(n_110),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_661),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_437),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_151),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_540),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_10),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_729),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_32),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_600),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_398),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_455),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_650),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_265),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_687),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_44),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_159),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_545),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_102),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_133),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_180),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_542),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_116),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_442),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_46),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_723),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_592),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_115),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_203),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_374),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_213),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_404),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_731),
.Y(n_1087)
);

BUFx8_ASAP7_75t_SL g1088 ( 
.A(n_262),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_144),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_584),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_280),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_699),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_264),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_371),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_326),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_235),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_511),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_106),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_70),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_491),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_657),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_86),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_531),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_77),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_702),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_329),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_173),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_262),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_158),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_655),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_722),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_588),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_227),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_334),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_204),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_409),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_737),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_28),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_421),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_355),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_534),
.Y(n_1121)
);

INVx5_ASAP7_75t_SL g1122 ( 
.A(n_207),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_673),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_70),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_211),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_19),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_151),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_644),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_387),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_319),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_390),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_31),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_483),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_375),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_181),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_558),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_452),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_89),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_203),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_675),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_563),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_355),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_321),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_172),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_425),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_234),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_403),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_162),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_617),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_263),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_463),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_437),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_6),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_253),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_475),
.Y(n_1155)
);

BUFx8_ASAP7_75t_SL g1156 ( 
.A(n_683),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_345),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_517),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_557),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_90),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_220),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_121),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_568),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_728),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_73),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_525),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_294),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_320),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_477),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_252),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_233),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_309),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_248),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_734),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_76),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_331),
.Y(n_1176)
);

BUFx5_ASAP7_75t_L g1177 ( 
.A(n_726),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_388),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_404),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_103),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_179),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_539),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_711),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_704),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_709),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_214),
.Y(n_1186)
);

INVxp33_ASAP7_75t_SL g1187 ( 
.A(n_116),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_37),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_632),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_464),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_572),
.Y(n_1191)
);

BUFx2_ASAP7_75t_R g1192 ( 
.A(n_331),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_164),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_357),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_664),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_505),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_671),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_413),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_668),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_554),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_596),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_613),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_198),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_551),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_674),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_654),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_530),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_677),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_247),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_535),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_680),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_478),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_235),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_191),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_55),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_670),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_314),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_20),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_538),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_715),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_676),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_735),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_251),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_132),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_354),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_336),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_114),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_267),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_52),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_505),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_14),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_638),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_529),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_292),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_130),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_466),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_458),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_47),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_242),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_254),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_293),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_132),
.Y(n_1242)
);

BUFx8_ASAP7_75t_SL g1243 ( 
.A(n_418),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_277),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_478),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_377),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_697),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_100),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_398),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_334),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_495),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_720),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_122),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_215),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_656),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_703),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_15),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_244),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_686),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_138),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_137),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_170),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_713),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_412),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_281),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_537),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_245),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_449),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_481),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_520),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_376),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_513),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_748),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_830),
.B(n_0),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_748),
.Y(n_1275)
);

INVxp33_ASAP7_75t_L g1276 ( 
.A(n_755),
.Y(n_1276)
);

BUFx2_ASAP7_75t_SL g1277 ( 
.A(n_1201),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_943),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_943),
.Y(n_1279)
);

CKINVDCx16_ASAP7_75t_R g1280 ( 
.A(n_1056),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_772),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1056),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_772),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_833),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_861),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_833),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_1066),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1109),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_842),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_842),
.Y(n_1290)
);

INVxp33_ASAP7_75t_SL g1291 ( 
.A(n_1227),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_895),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_895),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_896),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_963),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_896),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1086),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_770),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_770),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_955),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1086),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1102),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_829),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_963),
.Y(n_1304)
);

INVxp33_ASAP7_75t_SL g1305 ( 
.A(n_1094),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_770),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_770),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1258),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1102),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1134),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1134),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_770),
.Y(n_1312)
);

INVxp67_ASAP7_75t_SL g1313 ( 
.A(n_764),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_770),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_770),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1088),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_740),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1088),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_753),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_756),
.Y(n_1320)
);

INVxp33_ASAP7_75t_L g1321 ( 
.A(n_1243),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_767),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_777),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_764),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_776),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1243),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1156),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_776),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_782),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_784),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1156),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_836),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_862),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_778),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_836),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_776),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1039),
.Y(n_1337)
);

INVxp33_ASAP7_75t_SL g1338 ( 
.A(n_796),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_785),
.Y(n_1339)
);

CKINVDCx14_ASAP7_75t_R g1340 ( 
.A(n_1201),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_789),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_793),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_799),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_859),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_802),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_809),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_810),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_816),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_985),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_820),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_825),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1201),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_834),
.Y(n_1353)
);

INVxp33_ASAP7_75t_L g1354 ( 
.A(n_835),
.Y(n_1354)
);

CKINVDCx16_ASAP7_75t_R g1355 ( 
.A(n_993),
.Y(n_1355)
);

INVxp33_ASAP7_75t_L g1356 ( 
.A(n_840),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_841),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_843),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_846),
.Y(n_1359)
);

BUFx2_ASAP7_75t_SL g1360 ( 
.A(n_1263),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_851),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_862),
.Y(n_1362)
);

INVxp33_ASAP7_75t_SL g1363 ( 
.A(n_741),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_864),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_868),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_871),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_872),
.Y(n_1367)
);

INVxp33_ASAP7_75t_L g1368 ( 
.A(n_889),
.Y(n_1368)
);

INVxp33_ASAP7_75t_SL g1369 ( 
.A(n_743),
.Y(n_1369)
);

CKINVDCx16_ASAP7_75t_R g1370 ( 
.A(n_1254),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_908),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_909),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_912),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_882),
.Y(n_1374)
);

CKINVDCx14_ASAP7_75t_R g1375 ( 
.A(n_1263),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_882),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_877),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_923),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_924),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_776),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_928),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_931),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_935),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_824),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_950),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_877),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_945),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_752),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_940),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_954),
.Y(n_1390)
);

INVxp33_ASAP7_75t_SL g1391 ( 
.A(n_747),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_958),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_L g1393 ( 
.A(n_894),
.B(n_0),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_945),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_961),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_964),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_972),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_988),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1187),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_979),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_940),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_979),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_751),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_989),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_949),
.Y(n_1405)
);

CKINVDCx16_ASAP7_75t_R g1406 ( 
.A(n_1255),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1020),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1022),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1034),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_754),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_829),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1325),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1328),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1277),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1312),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1340),
.B(n_1122),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1314),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1303),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1352),
.B(n_801),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1303),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1334),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1337),
.B(n_997),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1273),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1303),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1411),
.Y(n_1425)
);

INVx5_ASAP7_75t_L g1426 ( 
.A(n_1411),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1315),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1411),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

OAI22x1_ASAP7_75t_R g1430 ( 
.A1(n_1304),
.A2(n_749),
.B1(n_837),
.B2(n_769),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1344),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1349),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_1280),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1336),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1327),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1285),
.B(n_997),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1380),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1317),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1384),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1298),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1285),
.B(n_1045),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_807),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1319),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1300),
.A2(n_769),
.B1(n_837),
.B2(n_749),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1300),
.A2(n_1308),
.B1(n_1305),
.B2(n_1291),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1275),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1299),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1331),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1320),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1306),
.A2(n_779),
.B(n_746),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1274),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1363),
.B(n_1200),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1322),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1360),
.B(n_1122),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1307),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_L g1456 ( 
.A(n_1281),
.B(n_761),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1287),
.B(n_1045),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1278),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1323),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1276),
.B(n_1122),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1283),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1308),
.A2(n_1031),
.B1(n_1037),
.B2(n_949),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1284),
.B(n_1232),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1286),
.B(n_804),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1289),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1333),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1329),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1290),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1292),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1330),
.Y(n_1470)
);

XNOR2x2_ASAP7_75t_L g1471 ( 
.A(n_1362),
.B(n_1192),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1339),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1342),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1279),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1343),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1345),
.A2(n_919),
.B(n_745),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1293),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1287),
.B(n_1051),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1294),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1296),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1346),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1388),
.A2(n_1037),
.B1(n_1072),
.B2(n_1031),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1377),
.Y(n_1483)
);

CKINVDCx6p67_ASAP7_75t_R g1484 ( 
.A(n_1406),
.Y(n_1484)
);

AND2x6_ASAP7_75t_L g1485 ( 
.A(n_1297),
.B(n_761),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1347),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

BUFx8_ASAP7_75t_L g1488 ( 
.A(n_1321),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1313),
.B(n_1051),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1403),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1350),
.Y(n_1491)
);

XNOR2x2_ASAP7_75t_L g1492 ( 
.A(n_1386),
.B(n_758),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1354),
.B(n_838),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1313),
.B(n_1091),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1351),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1301),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1353),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1302),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1295),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1357),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1309),
.B(n_821),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1332),
.B(n_1091),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1358),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1355),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1316),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1359),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1310),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1361),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1311),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1364),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1410),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1365),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1366),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1367),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1370),
.A2(n_1164),
.B1(n_1206),
.B2(n_1072),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1371),
.A2(n_919),
.B(n_745),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1409),
.A2(n_856),
.B(n_826),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1332),
.B(n_1265),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1338),
.Y(n_1519)
);

XOR2xp5_ASAP7_75t_L g1520 ( 
.A(n_1389),
.B(n_1269),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1372),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1374),
.B(n_1265),
.Y(n_1522)
);

INVxp33_ASAP7_75t_SL g1523 ( 
.A(n_1318),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1401),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1373),
.A2(n_898),
.B(n_874),
.Y(n_1525)
);

OAI22x1_ASAP7_75t_L g1526 ( 
.A1(n_1288),
.A2(n_813),
.B1(n_867),
.B2(n_839),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1378),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1374),
.B(n_905),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1379),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1381),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1382),
.Y(n_1531)
);

BUFx8_ASAP7_75t_L g1532 ( 
.A(n_1383),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1326),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1390),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1356),
.B(n_1368),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1376),
.B(n_786),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1376),
.B(n_1394),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1434),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1440),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1466),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1490),
.B(n_1399),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1468),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1469),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1536),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1477),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1479),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1480),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1434),
.Y(n_1549)
);

AND2x6_ASAP7_75t_L g1550 ( 
.A(n_1416),
.B(n_951),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1439),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1498),
.Y(n_1552)
);

AND2x2_ASAP7_75t_R g1553 ( 
.A(n_1430),
.B(n_1405),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1454),
.B(n_1394),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1507),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1504),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1438),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1439),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1493),
.B(n_1460),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1412),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1443),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1504),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1415),
.B(n_1369),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1449),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1413),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1453),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1459),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1418),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1467),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1437),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1421),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1447),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1470),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1475),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1455),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1472),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1452),
.A2(n_1391),
.B1(n_1206),
.B2(n_1252),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1481),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1414),
.B(n_1442),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1538),
.B(n_1519),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1483),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1418),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1417),
.B(n_1400),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1486),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1420),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1472),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1487),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1473),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1421),
.B(n_1288),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1420),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1495),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1473),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1424),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1424),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1491),
.Y(n_1595)
);

AND2x6_ASAP7_75t_L g1596 ( 
.A(n_1489),
.B(n_951),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1497),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1427),
.B(n_1400),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1500),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1425),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1503),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1425),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1506),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1519),
.B(n_1511),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1428),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1476),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1513),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1521),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1524),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1517),
.A2(n_1174),
.B(n_1136),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1527),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1519),
.B(n_1393),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1428),
.Y(n_1615)
);

AND2x2_ASAP7_75t_SL g1616 ( 
.A(n_1433),
.B(n_1335),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1530),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1491),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1525),
.A2(n_1174),
.B(n_1136),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1508),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1508),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1429),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1435),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1510),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1485),
.B(n_1324),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1510),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1512),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1484),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1429),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1431),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1441),
.B(n_1282),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1512),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1441),
.B(n_1164),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1514),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1432),
.B(n_1324),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1457),
.B(n_1387),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1514),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1419),
.B(n_1392),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1528),
.B(n_1395),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1529),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1444),
.Y(n_1641)
);

BUFx8_ASAP7_75t_L g1642 ( 
.A(n_1533),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1529),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1531),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1485),
.B(n_1387),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1457),
.B(n_1478),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1531),
.Y(n_1647)
);

XNOR2xp5_ASAP7_75t_L g1648 ( 
.A(n_1520),
.B(n_1462),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1478),
.B(n_1535),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1534),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1534),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1445),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1422),
.B(n_1335),
.Y(n_1653)
);

INVx4_ASAP7_75t_L g1654 ( 
.A(n_1489),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1537),
.B(n_1396),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1450),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1423),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1446),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1465),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1509),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1426),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1461),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1537),
.B(n_1397),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1496),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1476),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1458),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1426),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1463),
.B(n_1398),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1458),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1426),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1464),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1501),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1516),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1494),
.B(n_762),
.C(n_757),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1671),
.B(n_1485),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1568),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1672),
.B(n_1638),
.Y(n_1677)
);

BUFx4f_ASAP7_75t_L g1678 ( 
.A(n_1550),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1568),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1560),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1589),
.B(n_1474),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1607),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1568),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1565),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1556),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1582),
.Y(n_1686)
);

BUFx8_ASAP7_75t_SL g1687 ( 
.A(n_1541),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1639),
.B(n_1494),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1623),
.Y(n_1689)
);

INVx8_ASAP7_75t_L g1690 ( 
.A(n_1610),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1635),
.B(n_1474),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1540),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1540),
.Y(n_1694)
);

INVx4_ASAP7_75t_L g1695 ( 
.A(n_1654),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1571),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1554),
.B(n_1502),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1557),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1570),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1554),
.A2(n_1259),
.B1(n_1252),
.B2(n_1502),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1572),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1561),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1668),
.B(n_1579),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1559),
.A2(n_1259),
.B1(n_1522),
.B2(n_1518),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1580),
.B(n_1596),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1636),
.B(n_1499),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1607),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1636),
.B(n_1499),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1616),
.B(n_1562),
.Y(n_1709)
);

INVxp33_ASAP7_75t_L g1710 ( 
.A(n_1629),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1630),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1581),
.B(n_1482),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1564),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1566),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1575),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1596),
.B(n_1518),
.Y(n_1716)
);

INVx4_ASAP7_75t_L g1717 ( 
.A(n_1596),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1596),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1641),
.A2(n_1451),
.B1(n_1516),
.B2(n_1526),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1543),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1545),
.B(n_1523),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1544),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1673),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1604),
.B(n_1613),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1666),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1563),
.B(n_1451),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1546),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1652),
.B(n_1515),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1604),
.B(n_1522),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1613),
.B(n_1422),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1646),
.A2(n_936),
.B1(n_944),
.B2(n_917),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1622),
.B(n_1505),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1547),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1582),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1653),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1655),
.B(n_1456),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1548),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1633),
.B(n_1448),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1655),
.B(n_1067),
.Y(n_1739)
);

AND2x2_ASAP7_75t_SL g1740 ( 
.A(n_1577),
.B(n_1471),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1649),
.B(n_917),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1669),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1552),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1567),
.A2(n_944),
.B1(n_1003),
.B2(n_936),
.Y(n_1744)
);

NOR2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1663),
.B(n_1488),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1569),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1663),
.B(n_1532),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1555),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_L g1749 ( 
.A(n_1674),
.B(n_765),
.C(n_763),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1573),
.Y(n_1750)
);

OAI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1583),
.A2(n_1012),
.B1(n_1013),
.B2(n_1003),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1673),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1582),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1598),
.B(n_849),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1662),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1631),
.B(n_1404),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1574),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1640),
.B(n_1012),
.Y(n_1758)
);

INVx5_ASAP7_75t_L g1759 ( 
.A(n_1550),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_L g1760 ( 
.A(n_1550),
.B(n_824),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1625),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1628),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1640),
.B(n_1013),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1605),
.B(n_1407),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1578),
.B(n_1001),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1593),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1584),
.B(n_1587),
.Y(n_1767)
);

BUFx10_ASAP7_75t_L g1768 ( 
.A(n_1550),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1665),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1665),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1591),
.B(n_1597),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1599),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1601),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1558),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1657),
.B(n_1408),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1558),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1642),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1603),
.B(n_1129),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1608),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1609),
.A2(n_992),
.B1(n_1073),
.B2(n_1071),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1612),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1617),
.Y(n_1782)
);

INVx4_ASAP7_75t_L g1783 ( 
.A(n_1661),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1576),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1645),
.B(n_1664),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1642),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1656),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1539),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1593),
.Y(n_1789)
);

NAND3xp33_ASAP7_75t_L g1790 ( 
.A(n_1542),
.B(n_768),
.C(n_766),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1648),
.Y(n_1791)
);

AND2x2_ASAP7_75t_SL g1792 ( 
.A(n_1553),
.B(n_1492),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1586),
.Y(n_1793)
);

AND2x6_ASAP7_75t_L g1794 ( 
.A(n_1656),
.B(n_1658),
.Y(n_1794)
);

BUFx4f_ASAP7_75t_L g1795 ( 
.A(n_1593),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1600),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1620),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1621),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1600),
.Y(n_1799)
);

BUFx4f_ASAP7_75t_L g1800 ( 
.A(n_1600),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1624),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1588),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1626),
.B(n_1238),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1644),
.Y(n_1804)
);

NAND2xp33_ASAP7_75t_R g1805 ( 
.A(n_1611),
.B(n_1520),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1650),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1592),
.A2(n_1073),
.B1(n_1079),
.B2(n_1071),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1606),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1659),
.B(n_1272),
.Y(n_1809)
);

AND2x4_ASAP7_75t_SL g1810 ( 
.A(n_1660),
.B(n_1595),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1618),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1627),
.B(n_780),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1632),
.Y(n_1813)
);

BUFx8_ASAP7_75t_SL g1814 ( 
.A(n_1634),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1656),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1637),
.B(n_781),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1606),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_SL g1818 ( 
.A(n_1643),
.B(n_1488),
.Y(n_1818)
);

NAND2xp33_ASAP7_75t_L g1819 ( 
.A(n_1661),
.B(n_824),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1647),
.B(n_783),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1606),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1651),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1549),
.A2(n_1104),
.B1(n_1131),
.B2(n_1079),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1611),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1614),
.B(n_1104),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1585),
.B(n_1253),
.Y(n_1826)
);

INVxp67_ASAP7_75t_SL g1827 ( 
.A(n_1585),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1670),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1590),
.B(n_1131),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1551),
.B(n_788),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1590),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1594),
.B(n_1260),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_SL g1833 ( 
.A(n_1661),
.B(n_1166),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1594),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1687),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1711),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1703),
.B(n_1602),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1690),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1724),
.B(n_1685),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1677),
.B(n_1602),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1679),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1728),
.A2(n_1218),
.B1(n_1223),
.B2(n_1166),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1690),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1706),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1708),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1688),
.B(n_1615),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1729),
.B(n_1615),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1679),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1697),
.B(n_956),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1692),
.A2(n_1223),
.B1(n_1231),
.B2(n_1218),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1725),
.B(n_1231),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1767),
.B(n_991),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1772),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1761),
.B(n_1011),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1721),
.B(n_1082),
.C(n_1078),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1772),
.B(n_1125),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1742),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1710),
.B(n_1235),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1681),
.B(n_1235),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1771),
.A2(n_1246),
.B(n_1152),
.C(n_1050),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1732),
.A2(n_1691),
.B1(n_1695),
.B2(n_1735),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1712),
.B(n_1236),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1691),
.B(n_1667),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_SL g1864 ( 
.A(n_1777),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1773),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1773),
.B(n_1036),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1730),
.B(n_1058),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1698),
.Y(n_1868)
);

BUFx5_ASAP7_75t_L g1869 ( 
.A(n_1815),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1779),
.B(n_1061),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1809),
.A2(n_1267),
.B(n_1270),
.C(n_1262),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1680),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1782),
.B(n_1063),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1702),
.B(n_1068),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1700),
.B(n_1236),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1713),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1780),
.B(n_1696),
.C(n_1744),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1787),
.A2(n_1619),
.B(n_844),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1689),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1714),
.B(n_1070),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1709),
.B(n_1240),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1786),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1746),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1695),
.A2(n_1244),
.B1(n_1245),
.B2(n_1240),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1750),
.B(n_1075),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1679),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1757),
.B(n_1076),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1762),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1781),
.B(n_1077),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1741),
.B(n_1244),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1752),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1738),
.B(n_1245),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1675),
.A2(n_932),
.B(n_934),
.C(n_921),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1684),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1759),
.B(n_1667),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1759),
.B(n_1667),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1716),
.B(n_1084),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1745),
.B(n_1093),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1693),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1694),
.B(n_1096),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1699),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1704),
.B(n_1269),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1817),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1764),
.A2(n_960),
.B1(n_980),
.B2(n_952),
.Y(n_1904)
);

O2A1O1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1765),
.A2(n_1107),
.B(n_1108),
.C(n_1097),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1701),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1715),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1785),
.B(n_1120),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1759),
.B(n_790),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1764),
.A2(n_999),
.B1(n_1006),
.B2(n_995),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1720),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1678),
.B(n_791),
.Y(n_1912)
);

INVx5_ASAP7_75t_L g1913 ( 
.A(n_1794),
.Y(n_1913)
);

INVxp67_ASAP7_75t_SL g1914 ( 
.A(n_1682),
.Y(n_1914)
);

A2O1A1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1678),
.A2(n_1016),
.B(n_1021),
.C(n_1015),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1815),
.A2(n_1619),
.B(n_744),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1739),
.B(n_1121),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1821),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1722),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1727),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1828),
.B(n_792),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1828),
.B(n_794),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1736),
.B(n_1791),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1733),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1825),
.B(n_795),
.Y(n_1925)
);

NOR2xp67_ASAP7_75t_L g1926 ( 
.A(n_1821),
.B(n_1030),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1754),
.B(n_1124),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1717),
.B(n_798),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1795),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1775),
.B(n_1126),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1737),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1717),
.B(n_800),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1775),
.B(n_1137),
.Y(n_1933)
);

A2O1A1Ixp33_ASAP7_75t_L g1934 ( 
.A1(n_1769),
.A2(n_1069),
.B(n_1090),
.C(n_1033),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1743),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1751),
.B(n_1143),
.C(n_1138),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1748),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1795),
.Y(n_1938)
);

NOR2xp67_ASAP7_75t_L g1939 ( 
.A(n_1821),
.B(n_1092),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1718),
.A2(n_803),
.B1(n_811),
.B2(n_805),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1755),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1682),
.B(n_1146),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_1814),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1707),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1707),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1723),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1731),
.B(n_831),
.C(n_818),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1723),
.B(n_1147),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1718),
.B(n_812),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1797),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1726),
.B(n_814),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1800),
.B(n_817),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_1760),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1827),
.B(n_1155),
.Y(n_1954)
);

NAND2xp33_ASAP7_75t_L g1955 ( 
.A(n_1794),
.B(n_1705),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1740),
.A2(n_1263),
.B1(n_850),
.B2(n_927),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1769),
.B(n_1157),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1798),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1770),
.B(n_1158),
.Y(n_1959)
);

NAND2xp33_ASAP7_75t_L g1960 ( 
.A(n_1794),
.B(n_822),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1770),
.A2(n_823),
.B1(n_828),
.B2(n_827),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1807),
.A2(n_838),
.B1(n_927),
.B2(n_850),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1801),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1833),
.B(n_832),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1804),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1758),
.B(n_1763),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1676),
.B(n_1160),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1784),
.Y(n_1968)
);

NOR2xp67_ASAP7_75t_SL g1969 ( 
.A(n_1790),
.B(n_845),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1813),
.B(n_848),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1676),
.B(n_1165),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1683),
.B(n_1167),
.Y(n_1972)
);

AND2x6_ASAP7_75t_SL g1973 ( 
.A(n_1829),
.B(n_1169),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1683),
.B(n_1734),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1734),
.B(n_1753),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1806),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1800),
.B(n_852),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1686),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1793),
.Y(n_1979)
);

INVx8_ASAP7_75t_L g1980 ( 
.A(n_1756),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1753),
.B(n_1170),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1802),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1778),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1822),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1808),
.B(n_1186),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1803),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1811),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1749),
.A2(n_855),
.B1(n_857),
.B2(n_854),
.Y(n_1988)
);

INVx8_ASAP7_75t_L g1989 ( 
.A(n_1756),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1686),
.B(n_858),
.Y(n_1990)
);

NOR2x1p5_ASAP7_75t_L g1991 ( 
.A(n_1783),
.B(n_1789),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1808),
.B(n_1188),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1774),
.B(n_1190),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1823),
.B(n_838),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1719),
.B(n_850),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1776),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1783),
.B(n_1196),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1686),
.B(n_866),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1766),
.Y(n_1999)
);

INVx2_ASAP7_75t_SL g2000 ( 
.A(n_1796),
.Y(n_2000)
);

BUFx8_ASAP7_75t_L g2001 ( 
.A(n_1766),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1766),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1799),
.B(n_1198),
.Y(n_2003)
);

INVx4_ASAP7_75t_L g2004 ( 
.A(n_1799),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1831),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1799),
.B(n_1834),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1788),
.B(n_1210),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1836),
.Y(n_2008)
);

NAND2x1p5_ASAP7_75t_L g2009 ( 
.A(n_1903),
.B(n_1747),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1857),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1892),
.B(n_1812),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1853),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1963),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1875),
.A2(n_1792),
.B1(n_1820),
.B2(n_1816),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1862),
.A2(n_1805),
.B1(n_1818),
.B2(n_1794),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1965),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1839),
.B(n_1810),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1984),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1839),
.B(n_1830),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1861),
.B(n_1768),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1865),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_2001),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1837),
.B(n_1826),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1841),
.Y(n_2024)
);

BUFx8_ASAP7_75t_L g2025 ( 
.A(n_1864),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1845),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1923),
.B(n_1768),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1966),
.B(n_1832),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_2001),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1902),
.A2(n_938),
.B1(n_986),
.B2(n_927),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1842),
.A2(n_873),
.B1(n_876),
.B2(n_869),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1991),
.B(n_1824),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1911),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1859),
.B(n_938),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1852),
.B(n_1251),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1924),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_1888),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1931),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1929),
.B(n_1938),
.Y(n_2039)
);

OR2x6_ASAP7_75t_L g2040 ( 
.A(n_1980),
.B(n_1213),
.Y(n_2040)
);

AND3x1_ASAP7_75t_L g2041 ( 
.A(n_1850),
.B(n_1224),
.C(n_1217),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1844),
.B(n_938),
.Y(n_2042)
);

INVx5_ASAP7_75t_L g2043 ( 
.A(n_1913),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1879),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_R g2045 ( 
.A(n_1882),
.B(n_1819),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1851),
.B(n_878),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1980),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_SL g2048 ( 
.A(n_1835),
.B(n_986),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1858),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1840),
.B(n_1268),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1868),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1876),
.Y(n_2052)
);

NOR2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1838),
.B(n_880),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_SL g2054 ( 
.A1(n_1881),
.A2(n_1083),
.B1(n_1214),
.B2(n_986),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1843),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1883),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_SL g2057 ( 
.A(n_1855),
.B(n_885),
.C(n_884),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1989),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1849),
.B(n_1239),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1884),
.B(n_881),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1899),
.Y(n_2061)
);

INVx3_ASAP7_75t_SL g2062 ( 
.A(n_1943),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1937),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1950),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1890),
.B(n_886),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1841),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1958),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_R g2068 ( 
.A(n_1989),
.B(n_1918),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1856),
.B(n_1249),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1891),
.B(n_1257),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1898),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1913),
.B(n_887),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1983),
.B(n_1261),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1976),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1936),
.A2(n_1214),
.B1(n_1237),
.B2(n_1083),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1914),
.B(n_1264),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_1898),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1908),
.B(n_1266),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1867),
.B(n_888),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1919),
.Y(n_2080)
);

AO22x1_ASAP7_75t_L g2081 ( 
.A1(n_1964),
.A2(n_890),
.B1(n_897),
.B2(n_891),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1955),
.A2(n_1824),
.B(n_1222),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1920),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_2000),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1935),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1925),
.A2(n_900),
.B1(n_902),
.B2(n_901),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1913),
.B(n_1233),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1945),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2002),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1944),
.A2(n_904),
.B1(n_906),
.B2(n_903),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1946),
.Y(n_2091)
);

INVxp67_ASAP7_75t_L g2092 ( 
.A(n_1970),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1872),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1993),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_1918),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1994),
.A2(n_1214),
.B1(n_1237),
.B2(n_1083),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1841),
.Y(n_2097)
);

NOR3xp33_ASAP7_75t_L g2098 ( 
.A(n_1988),
.B(n_1271),
.C(n_1250),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1953),
.A2(n_1222),
.B(n_760),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1941),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1894),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1848),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_SL g2103 ( 
.A1(n_1951),
.A2(n_910),
.B1(n_913),
.B2(n_907),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1877),
.B(n_914),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1846),
.B(n_1219),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1901),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1848),
.B(n_915),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_1930),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_SL g2109 ( 
.A(n_1848),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1886),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1906),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2004),
.B(n_911),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1886),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1947),
.A2(n_1237),
.B1(n_918),
.B2(n_922),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_1995),
.A2(n_926),
.B1(n_933),
.B2(n_916),
.Y(n_2115)
);

BUFx2_ASAP7_75t_L g2116 ( 
.A(n_1886),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1854),
.B(n_941),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1978),
.B(n_942),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1907),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_1978),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_1933),
.B(n_946),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1968),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1979),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1967),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1973),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1971),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1986),
.B(n_947),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1978),
.B(n_948),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1999),
.B(n_911),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1917),
.B(n_957),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1982),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1972),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1981),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1985),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1974),
.Y(n_2135)
);

BUFx3_ASAP7_75t_L g2136 ( 
.A(n_1996),
.Y(n_2136)
);

AND3x1_ASAP7_75t_SL g2137 ( 
.A(n_2005),
.B(n_965),
.C(n_959),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1992),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1927),
.B(n_1225),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_1956),
.A2(n_968),
.B1(n_970),
.B2(n_967),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1961),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_1987),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_R g2143 ( 
.A(n_1960),
.B(n_971),
.Y(n_2143)
);

INVxp67_ASAP7_75t_SL g2144 ( 
.A(n_1847),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1940),
.B(n_973),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2006),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_2003),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1921),
.B(n_1229),
.Y(n_2148)
);

OR2x2_ASAP7_75t_SL g2149 ( 
.A(n_1997),
.B(n_892),
.Y(n_2149)
);

AND2x6_ASAP7_75t_L g2150 ( 
.A(n_1975),
.B(n_937),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1870),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1922),
.B(n_1230),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1954),
.B(n_1234),
.Y(n_2153)
);

O2A1O1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_1860),
.A2(n_1191),
.B(n_1195),
.C(n_1141),
.Y(n_2154)
);

AND3x1_ASAP7_75t_L g2155 ( 
.A(n_1962),
.B(n_1199),
.C(n_1197),
.Y(n_2155)
);

INVxp67_ASAP7_75t_SL g2156 ( 
.A(n_1869),
.Y(n_2156)
);

INVx5_ASAP7_75t_L g2157 ( 
.A(n_1869),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1904),
.B(n_974),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1910),
.B(n_1209),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1957),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2007),
.B(n_978),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1866),
.B(n_1212),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_2092),
.B(n_1952),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2011),
.B(n_1977),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_2044),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2108),
.B(n_1897),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2141),
.B(n_1990),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2034),
.B(n_1874),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2013),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_2043),
.B(n_1869),
.Y(n_2170)
);

AND3x1_ASAP7_75t_SL g2171 ( 
.A(n_2053),
.B(n_982),
.C(n_981),
.Y(n_2171)
);

OR2x6_ASAP7_75t_L g2172 ( 
.A(n_2022),
.B(n_1926),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2084),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2160),
.B(n_1880),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2051),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_2008),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_2029),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_2043),
.B(n_1869),
.Y(n_2178)
);

BUFx2_ASAP7_75t_L g2179 ( 
.A(n_2156),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2018),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2052),
.Y(n_2181)
);

INVxp67_ASAP7_75t_SL g2182 ( 
.A(n_2074),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2049),
.B(n_2151),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2016),
.Y(n_2184)
);

CKINVDCx20_ASAP7_75t_R g2185 ( 
.A(n_2025),
.Y(n_2185)
);

CKINVDCx20_ASAP7_75t_R g2186 ( 
.A(n_2025),
.Y(n_2186)
);

CKINVDCx8_ASAP7_75t_R g2187 ( 
.A(n_2010),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_2068),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2124),
.B(n_1885),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2126),
.B(n_1887),
.Y(n_2190)
);

INVx6_ASAP7_75t_L g2191 ( 
.A(n_2040),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_2026),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2060),
.A2(n_1939),
.B1(n_1912),
.B2(n_1998),
.Y(n_2193)
);

NAND2x1p5_ASAP7_75t_L g2194 ( 
.A(n_2043),
.B(n_1895),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2056),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_2032),
.B(n_1915),
.Y(n_2196)
);

NAND2x1p5_ASAP7_75t_L g2197 ( 
.A(n_2037),
.B(n_1896),
.Y(n_2197)
);

INVx5_ASAP7_75t_L g2198 ( 
.A(n_2024),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2065),
.B(n_1889),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2080),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2148),
.A2(n_1942),
.B1(n_1948),
.B2(n_1900),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2088),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2132),
.B(n_1873),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2091),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_2055),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2062),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2154),
.A2(n_1905),
.B(n_1871),
.C(n_1934),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_2109),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2041),
.B(n_983),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2133),
.B(n_1959),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2134),
.B(n_1969),
.Y(n_2211)
);

INVx4_ASAP7_75t_L g2212 ( 
.A(n_2024),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2033),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2064),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2138),
.B(n_1909),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2067),
.Y(n_2216)
);

OR2x6_ASAP7_75t_L g2217 ( 
.A(n_2040),
.B(n_1863),
.Y(n_2217)
);

NOR2xp67_ASAP7_75t_L g2218 ( 
.A(n_2047),
.B(n_1928),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_2089),
.Y(n_2219)
);

BUFx8_ASAP7_75t_L g2220 ( 
.A(n_2071),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2036),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2032),
.B(n_1932),
.Y(n_2222)
);

NAND2x1p5_ASAP7_75t_L g2223 ( 
.A(n_2058),
.B(n_1949),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2145),
.A2(n_987),
.B1(n_990),
.B2(n_984),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2061),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2113),
.Y(n_2226)
);

BUFx2_ASAP7_75t_L g2227 ( 
.A(n_2135),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_2046),
.B(n_996),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2077),
.B(n_2039),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2120),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2038),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2094),
.B(n_998),
.Y(n_2232)
);

BUFx2_ASAP7_75t_L g2233 ( 
.A(n_2135),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2083),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_2015),
.B(n_1893),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_2135),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2161),
.B(n_1242),
.Y(n_2237)
);

BUFx4f_ASAP7_75t_L g2238 ( 
.A(n_2009),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2045),
.Y(n_2239)
);

NAND2x1_ASAP7_75t_L g2240 ( 
.A(n_2024),
.B(n_1878),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2147),
.B(n_1004),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2127),
.B(n_1005),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2014),
.B(n_2012),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2103),
.B(n_1007),
.Y(n_2244)
);

BUFx2_ASAP7_75t_L g2245 ( 
.A(n_2097),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2039),
.B(n_1916),
.Y(n_2246)
);

CKINVDCx20_ASAP7_75t_R g2247 ( 
.A(n_2125),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2085),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_2066),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2021),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2031),
.B(n_1008),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2019),
.B(n_1211),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2078),
.B(n_1009),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2066),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2042),
.B(n_1207),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_2102),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2100),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2063),
.Y(n_2258)
);

NAND2x1p5_ASAP7_75t_L g2259 ( 
.A(n_2157),
.B(n_937),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2153),
.B(n_1017),
.Y(n_2260)
);

BUFx3_ASAP7_75t_L g2261 ( 
.A(n_2116),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2144),
.B(n_1018),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2066),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_SL g2264 ( 
.A1(n_2081),
.A2(n_1024),
.B1(n_1025),
.B2(n_1019),
.Y(n_2264)
);

INVxp67_ASAP7_75t_L g2265 ( 
.A(n_2028),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2079),
.B(n_1027),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2017),
.B(n_1101),
.Y(n_2267)
);

CKINVDCx8_ASAP7_75t_R g2268 ( 
.A(n_2087),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2121),
.B(n_1228),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2106),
.Y(n_2270)
);

INVx4_ASAP7_75t_L g2271 ( 
.A(n_2110),
.Y(n_2271)
);

BUFx4f_ASAP7_75t_SL g2272 ( 
.A(n_2136),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2119),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2093),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2162),
.B(n_1028),
.Y(n_2275)
);

NOR2xp67_ASAP7_75t_L g2276 ( 
.A(n_2095),
.B(n_546),
.Y(n_2276)
);

AOI22x1_ASAP7_75t_L g2277 ( 
.A1(n_2099),
.A2(n_1032),
.B1(n_1035),
.B2(n_1029),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2057),
.B(n_2152),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2101),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_2157),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2157),
.Y(n_2281)
);

AND2x6_ASAP7_75t_L g2282 ( 
.A(n_2110),
.B(n_1202),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2111),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2122),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2117),
.B(n_1044),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2123),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2131),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2110),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2086),
.B(n_1203),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2142),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2087),
.Y(n_2291)
);

BUFx3_ASAP7_75t_L g2292 ( 
.A(n_2129),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2146),
.Y(n_2293)
);

AOI221xp5_ASAP7_75t_L g2294 ( 
.A1(n_2098),
.A2(n_1052),
.B1(n_1054),
.B2(n_1049),
.C(n_1048),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2129),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2112),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2143),
.B(n_1221),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_2112),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2130),
.B(n_1055),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2149),
.Y(n_2300)
);

OR2x6_ASAP7_75t_SL g2301 ( 
.A(n_2090),
.B(n_1059),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2155),
.A2(n_2048),
.B1(n_2115),
.B2(n_2054),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2027),
.B(n_1101),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2139),
.B(n_1060),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2030),
.B(n_1065),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2023),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2035),
.B(n_1074),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2104),
.Y(n_2308)
);

BUFx2_ASAP7_75t_L g2309 ( 
.A(n_2150),
.Y(n_2309)
);

AOI21xp33_ASAP7_75t_L g2310 ( 
.A1(n_2158),
.A2(n_1208),
.B(n_1140),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2076),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2069),
.B(n_1085),
.Y(n_2312)
);

INVx2_ASAP7_75t_SL g2313 ( 
.A(n_2107),
.Y(n_2313)
);

INVx1_ASAP7_75t_SL g2314 ( 
.A(n_2118),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2059),
.B(n_1089),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2070),
.B(n_1095),
.Y(n_2316)
);

BUFx4f_ASAP7_75t_L g2317 ( 
.A(n_2150),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2073),
.Y(n_2318)
);

AOI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2201),
.A2(n_2082),
.B(n_2020),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2199),
.B(n_2050),
.Y(n_2320)
);

OAI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2242),
.A2(n_2105),
.B(n_2159),
.Y(n_2321)
);

CKINVDCx11_ASAP7_75t_R g2322 ( 
.A(n_2185),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_2165),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2179),
.A2(n_2072),
.B(n_2128),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2200),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2164),
.A2(n_2114),
.B(n_2140),
.Y(n_2326)
);

OAI21x1_ASAP7_75t_L g2327 ( 
.A1(n_2240),
.A2(n_2150),
.B(n_2096),
.Y(n_2327)
);

AOI21x1_ASAP7_75t_L g2328 ( 
.A1(n_2235),
.A2(n_2150),
.B(n_2137),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2168),
.B(n_2075),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2169),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2175),
.Y(n_2331)
);

OAI21x1_ASAP7_75t_L g2332 ( 
.A1(n_2170),
.A2(n_1177),
.B(n_549),
.Y(n_2332)
);

AO31x2_ASAP7_75t_L g2333 ( 
.A1(n_2309),
.A2(n_1140),
.A3(n_1208),
.B(n_1177),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_2178),
.A2(n_1177),
.B(n_550),
.Y(n_2334)
);

AO21x1_ASAP7_75t_L g2335 ( 
.A1(n_2278),
.A2(n_1177),
.B(n_1099),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2306),
.B(n_1098),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2181),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2189),
.B(n_2190),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_2261),
.Y(n_2339)
);

AOI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2179),
.A2(n_892),
.B(n_824),
.Y(n_2340)
);

NAND3xp33_ASAP7_75t_L g2341 ( 
.A(n_2244),
.B(n_1103),
.C(n_1100),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2195),
.Y(n_2342)
);

OAI21x1_ASAP7_75t_SL g2343 ( 
.A1(n_2211),
.A2(n_1),
.B(n_2),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2280),
.A2(n_953),
.B(n_892),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_2165),
.Y(n_2345)
);

OAI21x1_ASAP7_75t_L g2346 ( 
.A1(n_2250),
.A2(n_1177),
.B(n_552),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2301),
.A2(n_1113),
.B1(n_1114),
.B2(n_1106),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2280),
.A2(n_953),
.B(n_892),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2281),
.A2(n_975),
.B(n_953),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2188),
.B(n_953),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2182),
.B(n_1115),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_2186),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2281),
.A2(n_1000),
.B(n_975),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_SL g2354 ( 
.A1(n_2243),
.A2(n_1),
.B(n_2),
.Y(n_2354)
);

NAND3xp33_ASAP7_75t_L g2355 ( 
.A(n_2264),
.B(n_1118),
.C(n_1116),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2265),
.B(n_1119),
.Y(n_2356)
);

OAI21x1_ASAP7_75t_SL g2357 ( 
.A1(n_2193),
.A2(n_3),
.B(n_4),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_L g2358 ( 
.A1(n_2234),
.A2(n_1177),
.B(n_553),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2174),
.B(n_1127),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_SL g2360 ( 
.A(n_2238),
.B(n_742),
.Y(n_2360)
);

OAI21x1_ASAP7_75t_L g2361 ( 
.A1(n_2248),
.A2(n_1177),
.B(n_555),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2224),
.A2(n_2251),
.B(n_2207),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2289),
.A2(n_1241),
.B(n_1179),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2318),
.B(n_1130),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2205),
.Y(n_2365)
);

AO31x2_ASAP7_75t_L g2366 ( 
.A1(n_2309),
.A2(n_829),
.A3(n_556),
.B(n_560),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2166),
.B(n_1132),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2209),
.A2(n_975),
.B1(n_1010),
.B2(n_1000),
.Y(n_2368)
);

AO31x2_ASAP7_75t_L g2369 ( 
.A1(n_2270),
.A2(n_829),
.A3(n_561),
.B(n_565),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2205),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2214),
.B(n_975),
.Y(n_2371)
);

AO31x2_ASAP7_75t_L g2372 ( 
.A1(n_2273),
.A2(n_2257),
.A3(n_2233),
.B(n_2236),
.Y(n_2372)
);

BUFx2_ASAP7_75t_L g2373 ( 
.A(n_2272),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2260),
.A2(n_1194),
.B(n_1180),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2203),
.B(n_1133),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_L g2376 ( 
.A1(n_2216),
.A2(n_567),
.B(n_547),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2311),
.B(n_2210),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2225),
.B(n_1000),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2196),
.A2(n_2246),
.B(n_2222),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2176),
.B(n_1135),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2180),
.B(n_1139),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2192),
.B(n_1142),
.Y(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2259),
.A2(n_571),
.B(n_570),
.Y(n_2383)
);

AOI21xp33_ASAP7_75t_L g2384 ( 
.A1(n_2310),
.A2(n_1145),
.B(n_1144),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2183),
.B(n_1148),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_SL g2386 ( 
.A(n_2187),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2167),
.B(n_1150),
.Y(n_2387)
);

AO31x2_ASAP7_75t_L g2388 ( 
.A1(n_2227),
.A2(n_574),
.A3(n_575),
.B(n_573),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2317),
.A2(n_1010),
.B(n_1000),
.Y(n_2389)
);

OAI21xp33_ASAP7_75t_L g2390 ( 
.A1(n_2228),
.A2(n_1153),
.B(n_1151),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2293),
.Y(n_2391)
);

OAI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2302),
.A2(n_2163),
.B1(n_2314),
.B2(n_2275),
.Y(n_2392)
);

OAI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2253),
.A2(n_1226),
.B(n_1171),
.Y(n_2393)
);

INVx1_ASAP7_75t_SL g2394 ( 
.A(n_2191),
.Y(n_2394)
);

AO21x1_ASAP7_75t_L g2395 ( 
.A1(n_2215),
.A2(n_1161),
.B(n_1154),
.Y(n_2395)
);

OAI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2266),
.A2(n_1175),
.B(n_1168),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2237),
.B(n_1162),
.Y(n_2397)
);

OAI21x1_ASAP7_75t_L g2398 ( 
.A1(n_2194),
.A2(n_578),
.B(n_577),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2184),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2202),
.Y(n_2400)
);

OAI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2299),
.A2(n_1215),
.B(n_1193),
.Y(n_2401)
);

NOR2x1_ASAP7_75t_SL g2402 ( 
.A(n_2198),
.B(n_1010),
.Y(n_2402)
);

AO31x2_ASAP7_75t_L g2403 ( 
.A1(n_2227),
.A2(n_580),
.A3(n_581),
.B(n_579),
.Y(n_2403)
);

AOI21x1_ASAP7_75t_L g2404 ( 
.A1(n_2233),
.A2(n_1014),
.B(n_1010),
.Y(n_2404)
);

OAI21x1_ASAP7_75t_L g2405 ( 
.A1(n_2308),
.A2(n_583),
.B(n_582),
.Y(n_2405)
);

NAND3xp33_ASAP7_75t_SL g2406 ( 
.A(n_2294),
.B(n_1173),
.C(n_1172),
.Y(n_2406)
);

OAI21x1_ASAP7_75t_L g2407 ( 
.A1(n_2197),
.A2(n_587),
.B(n_585),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2198),
.A2(n_1248),
.B(n_1014),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2204),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2198),
.A2(n_1248),
.B(n_1014),
.Y(n_2410)
);

BUFx12f_ASAP7_75t_L g2411 ( 
.A(n_2206),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2252),
.A2(n_1248),
.B(n_1014),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2274),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2304),
.A2(n_1248),
.B(n_759),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2300),
.A2(n_590),
.B(n_589),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2239),
.B(n_3),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2298),
.B(n_1176),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2219),
.B(n_1178),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2291),
.B(n_1181),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2173),
.B(n_1182),
.Y(n_2420)
);

AOI21x1_ASAP7_75t_L g2421 ( 
.A1(n_2236),
.A2(n_771),
.B(n_750),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2245),
.B(n_4),
.Y(n_2422)
);

AO21x1_ASAP7_75t_L g2423 ( 
.A1(n_2297),
.A2(n_5),
.B(n_7),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2245),
.B(n_5),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2191),
.Y(n_2425)
);

OAI21x1_ASAP7_75t_L g2426 ( 
.A1(n_2283),
.A2(n_595),
.B(n_593),
.Y(n_2426)
);

INVx5_ASAP7_75t_L g2427 ( 
.A(n_2208),
.Y(n_2427)
);

INVx5_ASAP7_75t_L g2428 ( 
.A(n_2282),
.Y(n_2428)
);

CKINVDCx8_ASAP7_75t_R g2429 ( 
.A(n_2206),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2286),
.Y(n_2430)
);

INVxp67_ASAP7_75t_L g2431 ( 
.A(n_2226),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2262),
.A2(n_774),
.B(n_773),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2305),
.A2(n_787),
.B1(n_797),
.B2(n_775),
.Y(n_2433)
);

BUFx4_ASAP7_75t_SL g2434 ( 
.A(n_2247),
.Y(n_2434)
);

OAI21x1_ASAP7_75t_L g2435 ( 
.A1(n_2213),
.A2(n_601),
.B(n_598),
.Y(n_2435)
);

OAI21xp33_ASAP7_75t_L g2436 ( 
.A1(n_2315),
.A2(n_2312),
.B(n_2316),
.Y(n_2436)
);

OAI21xp33_ASAP7_75t_L g2437 ( 
.A1(n_2307),
.A2(n_808),
.B(n_806),
.Y(n_2437)
);

OAI21x1_ASAP7_75t_L g2438 ( 
.A1(n_2221),
.A2(n_604),
.B(n_603),
.Y(n_2438)
);

OAI21x1_ASAP7_75t_L g2439 ( 
.A1(n_2231),
.A2(n_607),
.B(n_605),
.Y(n_2439)
);

AO21x1_ASAP7_75t_L g2440 ( 
.A1(n_2303),
.A2(n_9),
.B(n_10),
.Y(n_2440)
);

A2O1A1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_2313),
.A2(n_819),
.B(n_847),
.C(n_815),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2296),
.B(n_2282),
.Y(n_2442)
);

OAI21x1_ASAP7_75t_L g2443 ( 
.A1(n_2258),
.A2(n_610),
.B(n_609),
.Y(n_2443)
);

AOI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2276),
.A2(n_860),
.B(n_853),
.Y(n_2444)
);

BUFx5_ASAP7_75t_L g2445 ( 
.A(n_2282),
.Y(n_2445)
);

INVxp67_ASAP7_75t_L g2446 ( 
.A(n_2230),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2295),
.B(n_9),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2292),
.B(n_11),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2229),
.B(n_12),
.Y(n_2449)
);

AO31x2_ASAP7_75t_L g2450 ( 
.A1(n_2279),
.A2(n_2284),
.A3(n_2287),
.B(n_2290),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2269),
.B(n_12),
.Y(n_2451)
);

OAI21x1_ASAP7_75t_L g2452 ( 
.A1(n_2223),
.A2(n_612),
.B(n_611),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2249),
.B(n_863),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2288),
.A2(n_870),
.B(n_865),
.Y(n_2454)
);

OAI21x1_ASAP7_75t_L g2455 ( 
.A1(n_2277),
.A2(n_615),
.B(n_614),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2249),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2268),
.B(n_13),
.Y(n_2457)
);

OAI21x1_ASAP7_75t_L g2458 ( 
.A1(n_2218),
.A2(n_623),
.B(n_618),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2256),
.B(n_2255),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2232),
.B(n_13),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2177),
.B(n_16),
.Y(n_2461)
);

A2O1A1Ixp33_ASAP7_75t_L g2462 ( 
.A1(n_2285),
.A2(n_879),
.B(n_883),
.C(n_875),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2241),
.A2(n_920),
.B(n_899),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2320),
.B(n_2254),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2319),
.A2(n_2263),
.B(n_2254),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2431),
.B(n_2217),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2386),
.Y(n_2467)
);

O2A1O1Ixp5_ASAP7_75t_L g2468 ( 
.A1(n_2362),
.A2(n_2212),
.B(n_2271),
.C(n_2267),
.Y(n_2468)
);

BUFx8_ASAP7_75t_SL g2469 ( 
.A(n_2352),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2446),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2339),
.B(n_2263),
.Y(n_2471)
);

OR2x6_ASAP7_75t_L g2472 ( 
.A(n_2379),
.B(n_2217),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2331),
.Y(n_2473)
);

OR2x2_ASAP7_75t_L g2474 ( 
.A(n_2337),
.B(n_2172),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2394),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2338),
.B(n_2220),
.Y(n_2476)
);

INVx3_ASAP7_75t_L g2477 ( 
.A(n_2365),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2451),
.B(n_2172),
.Y(n_2478)
);

AO21x2_ASAP7_75t_L g2479 ( 
.A1(n_2404),
.A2(n_2171),
.B(n_1189),
.Y(n_2479)
);

OR2x6_ASAP7_75t_L g2480 ( 
.A(n_2411),
.B(n_625),
.Y(n_2480)
);

INVx1_ASAP7_75t_SL g2481 ( 
.A(n_2425),
.Y(n_2481)
);

O2A1O1Ixp5_ASAP7_75t_SL g2482 ( 
.A1(n_2342),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2482)
);

AOI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2324),
.A2(n_925),
.B(n_893),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2370),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2340),
.A2(n_930),
.B(n_929),
.Y(n_2485)
);

AOI21xp5_ASAP7_75t_L g2486 ( 
.A1(n_2321),
.A2(n_962),
.B(n_939),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2377),
.B(n_2392),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2335),
.A2(n_969),
.B(n_966),
.Y(n_2488)
);

AOI221xp5_ASAP7_75t_L g2489 ( 
.A1(n_2326),
.A2(n_994),
.B1(n_1002),
.B2(n_977),
.C(n_976),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_2429),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2456),
.B(n_17),
.Y(n_2491)
);

A2O1A1Ixp33_ASAP7_75t_SL g2492 ( 
.A1(n_2420),
.A2(n_2387),
.B(n_2393),
.C(n_2374),
.Y(n_2492)
);

BUFx3_ASAP7_75t_L g2493 ( 
.A(n_2373),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2413),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2430),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2428),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2372),
.B(n_631),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2422),
.B(n_18),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_2344),
.A2(n_1026),
.B(n_1023),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2372),
.B(n_21),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2391),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2436),
.A2(n_1040),
.B1(n_1041),
.B2(n_1038),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2348),
.A2(n_1043),
.B(n_1042),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2349),
.A2(n_1047),
.B(n_1046),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_SL g2505 ( 
.A(n_2428),
.B(n_2360),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2450),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2450),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2427),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2351),
.B(n_21),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2353),
.A2(n_1057),
.B(n_1053),
.Y(n_2510)
);

CKINVDCx20_ASAP7_75t_R g2511 ( 
.A(n_2322),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2428),
.A2(n_1183),
.B1(n_1184),
.B2(n_1163),
.Y(n_2512)
);

OR2x6_ASAP7_75t_L g2513 ( 
.A(n_2442),
.B(n_634),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2427),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2323),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2327),
.A2(n_1064),
.B(n_1062),
.Y(n_2516)
);

NAND2x1p5_ASAP7_75t_L g2517 ( 
.A(n_2427),
.B(n_637),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_2459),
.Y(n_2518)
);

AOI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2389),
.A2(n_1081),
.B(n_1080),
.Y(n_2519)
);

OR2x6_ASAP7_75t_L g2520 ( 
.A(n_2345),
.B(n_639),
.Y(n_2520)
);

AOI21xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2347),
.A2(n_24),
.B(n_23),
.Y(n_2521)
);

CKINVDCx20_ASAP7_75t_R g2522 ( 
.A(n_2397),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2424),
.B(n_22),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2325),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2408),
.A2(n_1105),
.B(n_1087),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2330),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2329),
.B(n_23),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2449),
.B(n_24),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2399),
.Y(n_2529)
);

O2A1O1Ixp5_ASAP7_75t_L g2530 ( 
.A1(n_2328),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2371),
.B(n_26),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2400),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2350),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2409),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2378),
.Y(n_2535)
);

O2A1O1Ixp5_ASAP7_75t_L g2536 ( 
.A1(n_2423),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2375),
.B(n_29),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2367),
.B(n_30),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2410),
.A2(n_1111),
.B(n_1110),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2359),
.B(n_32),
.Y(n_2540)
);

OAI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2433),
.A2(n_1247),
.B1(n_1256),
.B2(n_1128),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2445),
.B(n_2440),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2434),
.Y(n_2543)
);

INVx3_ASAP7_75t_SL g2544 ( 
.A(n_2461),
.Y(n_2544)
);

A2O1A1Ixp33_ASAP7_75t_L g2545 ( 
.A1(n_2437),
.A2(n_1117),
.B(n_1123),
.C(n_1112),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2333),
.Y(n_2546)
);

A2O1A1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2341),
.A2(n_1159),
.B(n_1185),
.C(n_1149),
.Y(n_2547)
);

O2A1O1Ixp5_ASAP7_75t_SL g2548 ( 
.A1(n_2453),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_2548)
);

O2A1O1Ixp33_ASAP7_75t_L g2549 ( 
.A1(n_2363),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2333),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2416),
.B(n_36),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2445),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2445),
.B(n_37),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2445),
.B(n_38),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2448),
.B(n_38),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2457),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2381),
.Y(n_2557)
);

OR2x2_ASAP7_75t_SL g2558 ( 
.A(n_2355),
.B(n_39),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2380),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2447),
.Y(n_2560)
);

AOI222xp33_ASAP7_75t_L g2561 ( 
.A1(n_2390),
.A2(n_1220),
.B1(n_1205),
.B2(n_1216),
.C1(n_1204),
.C2(n_41),
.Y(n_2561)
);

NAND2x1_ASAP7_75t_L g2562 ( 
.A(n_2354),
.B(n_39),
.Y(n_2562)
);

A2O1A1Ixp33_ASAP7_75t_L g2563 ( 
.A1(n_2414),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2369),
.Y(n_2564)
);

BUFx4f_ASAP7_75t_L g2565 ( 
.A(n_2402),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2366),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2460),
.B(n_42),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2336),
.B(n_43),
.Y(n_2568)
);

INVx5_ASAP7_75t_L g2569 ( 
.A(n_2458),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2406),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2570)
);

HB1xp67_ASAP7_75t_L g2571 ( 
.A(n_2369),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2343),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2471),
.B(n_2464),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2470),
.B(n_2385),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2494),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2487),
.B(n_2364),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_2552),
.B(n_2388),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2473),
.Y(n_2578)
);

A2O1A1Ixp33_ASAP7_75t_L g2579 ( 
.A1(n_2492),
.A2(n_2384),
.B(n_2401),
.C(n_2396),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2495),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2501),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2518),
.B(n_2382),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2543),
.B(n_2418),
.Y(n_2583)
);

O2A1O1Ixp33_ASAP7_75t_L g2584 ( 
.A1(n_2521),
.A2(n_2462),
.B(n_2357),
.C(n_2463),
.Y(n_2584)
);

AOI21x1_ASAP7_75t_SL g2585 ( 
.A1(n_2523),
.A2(n_2419),
.B(n_2356),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_2469),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2560),
.B(n_2395),
.Y(n_2587)
);

A2O1A1Ixp33_ASAP7_75t_L g2588 ( 
.A1(n_2549),
.A2(n_2441),
.B(n_2432),
.C(n_2368),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2514),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2478),
.B(n_2493),
.Y(n_2590)
);

HB1xp67_ASAP7_75t_L g2591 ( 
.A(n_2474),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2500),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2535),
.B(n_2417),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2527),
.B(n_46),
.Y(n_2594)
);

BUFx3_ASAP7_75t_L g2595 ( 
.A(n_2511),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2526),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2559),
.B(n_47),
.Y(n_2597)
);

OAI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2570),
.A2(n_2421),
.B1(n_2454),
.B2(n_2444),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2508),
.B(n_2388),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2472),
.B(n_2403),
.Y(n_2600)
);

AOI21xp5_ASAP7_75t_SL g2601 ( 
.A1(n_2513),
.A2(n_2412),
.B(n_2366),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2556),
.B(n_48),
.Y(n_2602)
);

INVx2_ASAP7_75t_SL g2603 ( 
.A(n_2515),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2477),
.B(n_2452),
.Y(n_2604)
);

AND2x4_ASAP7_75t_L g2605 ( 
.A(n_2472),
.B(n_2497),
.Y(n_2605)
);

BUFx12f_ASAP7_75t_L g2606 ( 
.A(n_2533),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2466),
.B(n_48),
.Y(n_2607)
);

NOR2xp67_ASAP7_75t_L g2608 ( 
.A(n_2476),
.B(n_2465),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2544),
.B(n_2498),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2484),
.B(n_2403),
.Y(n_2610)
);

OAI22xp5_ASAP7_75t_SL g2611 ( 
.A1(n_2558),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2572),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2497),
.B(n_2415),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2532),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2524),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2555),
.B(n_2467),
.Y(n_2616)
);

OR2x2_ASAP7_75t_SL g2617 ( 
.A(n_2496),
.B(n_2553),
.Y(n_2617)
);

HB1xp67_ASAP7_75t_L g2618 ( 
.A(n_2571),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2475),
.B(n_2407),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2481),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2567),
.B(n_50),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2491),
.B(n_51),
.Y(n_2622)
);

OA22x2_ASAP7_75t_L g2623 ( 
.A1(n_2513),
.A2(n_2358),
.B1(n_2361),
.B2(n_2346),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2496),
.B(n_2398),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2568),
.B(n_53),
.Y(n_2625)
);

O2A1O1Ixp5_ASAP7_75t_L g2626 ( 
.A1(n_2542),
.A2(n_64),
.B(n_73),
.C(n_53),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2490),
.B(n_2376),
.Y(n_2627)
);

AND2x4_ASAP7_75t_L g2628 ( 
.A(n_2496),
.B(n_2566),
.Y(n_2628)
);

AND2x2_ASAP7_75t_L g2629 ( 
.A(n_2528),
.B(n_2332),
.Y(n_2629)
);

INVxp67_ASAP7_75t_L g2630 ( 
.A(n_2557),
.Y(n_2630)
);

OA21x2_ASAP7_75t_L g2631 ( 
.A1(n_2564),
.A2(n_2426),
.B(n_2405),
.Y(n_2631)
);

CKINVDCx11_ASAP7_75t_R g2632 ( 
.A(n_2522),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2534),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2551),
.B(n_2334),
.Y(n_2634)
);

OR2x6_ASAP7_75t_L g2635 ( 
.A(n_2480),
.B(n_2383),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2529),
.Y(n_2636)
);

INVx2_ASAP7_75t_SL g2637 ( 
.A(n_2533),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2507),
.Y(n_2638)
);

OA21x2_ASAP7_75t_L g2639 ( 
.A1(n_2550),
.A2(n_2455),
.B(n_2438),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2509),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2480),
.B(n_54),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2506),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2546),
.B(n_2435),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2505),
.B(n_2439),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2516),
.A2(n_2443),
.B(n_56),
.Y(n_2645)
);

NAND2x1p5_ASAP7_75t_L g2646 ( 
.A(n_2565),
.B(n_640),
.Y(n_2646)
);

HB1xp67_ASAP7_75t_L g2647 ( 
.A(n_2531),
.Y(n_2647)
);

BUFx4f_ASAP7_75t_L g2648 ( 
.A(n_2517),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2554),
.Y(n_2649)
);

O2A1O1Ixp33_ASAP7_75t_L g2650 ( 
.A1(n_2563),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2569),
.B(n_57),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2520),
.B(n_58),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2540),
.B(n_59),
.Y(n_2653)
);

A2O1A1Ixp33_ASAP7_75t_L g2654 ( 
.A1(n_2536),
.A2(n_63),
.B(n_59),
.C(n_61),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2562),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2569),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2590),
.B(n_2538),
.Y(n_2657)
);

OAI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2576),
.A2(n_2520),
.B1(n_2537),
.B2(n_2569),
.Y(n_2658)
);

CKINVDCx6p67_ASAP7_75t_R g2659 ( 
.A(n_2632),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2575),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2575),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_SL g2662 ( 
.A(n_2595),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2578),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2580),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2603),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2648),
.Y(n_2666)
);

INVxp67_ASAP7_75t_L g2667 ( 
.A(n_2612),
.Y(n_2667)
);

AOI21x1_ASAP7_75t_L g2668 ( 
.A1(n_2587),
.A2(n_2486),
.B(n_2483),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2573),
.B(n_2468),
.Y(n_2669)
);

BUFx12f_ASAP7_75t_L g2670 ( 
.A(n_2586),
.Y(n_2670)
);

AOI21x1_ASAP7_75t_L g2671 ( 
.A1(n_2608),
.A2(n_2488),
.B(n_2485),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2606),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2589),
.Y(n_2673)
);

INVx6_ASAP7_75t_L g2674 ( 
.A(n_2609),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2636),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2618),
.Y(n_2676)
);

OAI21x1_ASAP7_75t_L g2677 ( 
.A1(n_2623),
.A2(n_2482),
.B(n_2530),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2596),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2581),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2649),
.B(n_2479),
.Y(n_2680)
);

OAI21x1_ASAP7_75t_L g2681 ( 
.A1(n_2656),
.A2(n_2548),
.B(n_2503),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2614),
.Y(n_2682)
);

OA21x2_ASAP7_75t_L g2683 ( 
.A1(n_2656),
.A2(n_2502),
.B(n_2512),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_SL g2684 ( 
.A1(n_2611),
.A2(n_2561),
.B1(n_2541),
.B2(n_2499),
.Y(n_2684)
);

INVx3_ASAP7_75t_L g2685 ( 
.A(n_2589),
.Y(n_2685)
);

OAI21x1_ASAP7_75t_L g2686 ( 
.A1(n_2644),
.A2(n_2510),
.B(n_2504),
.Y(n_2686)
);

OAI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2601),
.A2(n_2642),
.B(n_2639),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2591),
.B(n_61),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2616),
.B(n_64),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2633),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2615),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2592),
.A2(n_2489),
.B1(n_2519),
.B2(n_2525),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2652),
.A2(n_2545),
.B1(n_2547),
.B2(n_2539),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2620),
.Y(n_2694)
);

AO31x2_ASAP7_75t_L g2695 ( 
.A1(n_2638),
.A2(n_67),
.A3(n_65),
.B(n_66),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2593),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2610),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2647),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2599),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2599),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2617),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2640),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2583),
.Y(n_2703)
);

OR2x6_ASAP7_75t_L g2704 ( 
.A(n_2605),
.B(n_641),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2577),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2628),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2577),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2619),
.Y(n_2708)
);

INVx4_ASAP7_75t_SL g2709 ( 
.A(n_2600),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2628),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2574),
.Y(n_2711)
);

HB1xp67_ASAP7_75t_L g2712 ( 
.A(n_2639),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2600),
.Y(n_2713)
);

OAI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2626),
.A2(n_65),
.B(n_66),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2605),
.Y(n_2715)
);

OAI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2579),
.A2(n_68),
.B(n_69),
.Y(n_2716)
);

AO22x2_ASAP7_75t_L g2717 ( 
.A1(n_2582),
.A2(n_71),
.B1(n_68),
.B2(n_69),
.Y(n_2717)
);

OAI21x1_ASAP7_75t_L g2718 ( 
.A1(n_2631),
.A2(n_71),
.B(n_72),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2655),
.Y(n_2719)
);

HB1xp67_ASAP7_75t_L g2720 ( 
.A(n_2631),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2643),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2653),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2630),
.B(n_74),
.Y(n_2723)
);

OAI21x1_ASAP7_75t_L g2724 ( 
.A1(n_2585),
.A2(n_76),
.B(n_79),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2643),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2604),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2602),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_2597),
.B(n_80),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2613),
.Y(n_2729)
);

OAI21x1_ASAP7_75t_L g2730 ( 
.A1(n_2627),
.A2(n_81),
.B(n_82),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2613),
.Y(n_2731)
);

AO21x1_ASAP7_75t_SL g2732 ( 
.A1(n_2607),
.A2(n_81),
.B(n_82),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2629),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2651),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2733),
.B(n_2634),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2720),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2719),
.B(n_2621),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2660),
.Y(n_2738)
);

INVxp67_ASAP7_75t_L g2739 ( 
.A(n_2662),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2733),
.B(n_2641),
.Y(n_2740)
);

INVx6_ASAP7_75t_L g2741 ( 
.A(n_2670),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2711),
.B(n_2594),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2661),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2727),
.B(n_2651),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2669),
.B(n_2637),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2673),
.Y(n_2746)
);

BUFx2_ASAP7_75t_L g2747 ( 
.A(n_2673),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2667),
.B(n_2622),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2676),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2676),
.B(n_2625),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2667),
.B(n_2624),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2720),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2709),
.B(n_2624),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2659),
.Y(n_2754)
);

NOR2x1_ASAP7_75t_L g2755 ( 
.A(n_2701),
.B(n_2635),
.Y(n_2755)
);

INVx1_ASAP7_75t_SL g2756 ( 
.A(n_2662),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2729),
.B(n_2635),
.Y(n_2757)
);

NOR3xp33_ASAP7_75t_L g2758 ( 
.A(n_2716),
.B(n_2650),
.C(n_2598),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2674),
.B(n_2648),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2698),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2712),
.Y(n_2761)
);

HB1xp67_ASAP7_75t_L g2762 ( 
.A(n_2712),
.Y(n_2762)
);

OR2x6_ASAP7_75t_L g2763 ( 
.A(n_2704),
.B(n_2646),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2708),
.B(n_2654),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2663),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2687),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2696),
.B(n_2731),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2674),
.B(n_2645),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2685),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2679),
.Y(n_2770)
);

BUFx2_ASAP7_75t_L g2771 ( 
.A(n_2685),
.Y(n_2771)
);

INVxp67_ASAP7_75t_SL g2772 ( 
.A(n_2680),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2726),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2709),
.B(n_2588),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2716),
.A2(n_2584),
.B1(n_85),
.B2(n_83),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2691),
.Y(n_2776)
);

INVxp67_ASAP7_75t_SL g2777 ( 
.A(n_2680),
.Y(n_2777)
);

INVxp67_ASAP7_75t_SL g2778 ( 
.A(n_2658),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2706),
.B(n_83),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2739),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2738),
.Y(n_2781)
);

OR2x2_ASAP7_75t_L g2782 ( 
.A(n_2749),
.B(n_2694),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2735),
.B(n_2665),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2740),
.B(n_2706),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2750),
.B(n_2688),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2755),
.B(n_2709),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2736),
.Y(n_2787)
);

BUFx2_ASAP7_75t_L g2788 ( 
.A(n_2754),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2736),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2752),
.Y(n_2790)
);

OR2x2_ASAP7_75t_L g2791 ( 
.A(n_2748),
.B(n_2742),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2743),
.Y(n_2792)
);

INVxp67_ASAP7_75t_L g2793 ( 
.A(n_2750),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2745),
.B(n_2657),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2747),
.B(n_2707),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2737),
.B(n_2658),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2765),
.Y(n_2797)
);

HB1xp67_ASAP7_75t_L g2798 ( 
.A(n_2761),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2768),
.B(n_2710),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2771),
.B(n_2700),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2754),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2770),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2760),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2752),
.Y(n_2804)
);

OR2x2_ASAP7_75t_L g2805 ( 
.A(n_2767),
.B(n_2734),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2776),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2759),
.B(n_2702),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2746),
.B(n_2705),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2746),
.B(n_2699),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2753),
.B(n_2713),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2776),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2746),
.B(n_2697),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2751),
.B(n_2664),
.Y(n_2813)
);

BUFx8_ASAP7_75t_SL g2814 ( 
.A(n_2779),
.Y(n_2814)
);

BUFx3_ASAP7_75t_L g2815 ( 
.A(n_2741),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2737),
.B(n_2728),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2797),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2780),
.B(n_2756),
.Y(n_2818)
);

AND2x2_ASAP7_75t_SL g2819 ( 
.A(n_2786),
.B(n_2758),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2802),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2793),
.B(n_2778),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2794),
.B(n_2784),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2786),
.B(n_2774),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2787),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2794),
.B(n_2769),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2815),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2786),
.B(n_2774),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2798),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2781),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2791),
.B(n_2764),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2784),
.B(n_2769),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2783),
.B(n_2769),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2783),
.B(n_2757),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2792),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2787),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2795),
.B(n_2757),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_SL g2837 ( 
.A1(n_2796),
.A2(n_2717),
.B1(n_2774),
.B2(n_2763),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2795),
.B(n_2741),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2803),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2798),
.Y(n_2840)
);

AND2x4_ASAP7_75t_L g2841 ( 
.A(n_2815),
.B(n_2810),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2789),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2789),
.Y(n_2843)
);

NAND2x1p5_ASAP7_75t_L g2844 ( 
.A(n_2801),
.B(n_2666),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2810),
.B(n_2790),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2800),
.B(n_2741),
.Y(n_2846)
);

HB1xp67_ASAP7_75t_L g2847 ( 
.A(n_2790),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2788),
.B(n_2703),
.Y(n_2848)
);

INVxp67_ASAP7_75t_SL g2849 ( 
.A(n_2804),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2804),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2814),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2805),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2813),
.Y(n_2853)
);

HB1xp67_ASAP7_75t_L g2854 ( 
.A(n_2785),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2782),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2800),
.B(n_2753),
.Y(n_2856)
);

OAI221xp5_ASAP7_75t_SL g2857 ( 
.A1(n_2837),
.A2(n_2775),
.B1(n_2722),
.B2(n_2816),
.C(n_2684),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2854),
.B(n_2772),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2851),
.Y(n_2859)
);

NAND2x1_ASAP7_75t_L g2860 ( 
.A(n_2841),
.B(n_2810),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2845),
.Y(n_2861)
);

INVx1_ASAP7_75t_SL g2862 ( 
.A(n_2819),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2822),
.B(n_2838),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2818),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2845),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2828),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2845),
.Y(n_2867)
);

INVx2_ASAP7_75t_SL g2868 ( 
.A(n_2846),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2828),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2836),
.Y(n_2870)
);

AOI211xp5_ASAP7_75t_L g2871 ( 
.A1(n_2821),
.A2(n_2823),
.B(n_2827),
.C(n_2819),
.Y(n_2871)
);

AOI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_2830),
.A2(n_2775),
.B1(n_2717),
.B2(n_2684),
.Y(n_2872)
);

NAND3xp33_ASAP7_75t_SL g2873 ( 
.A(n_2826),
.B(n_2722),
.C(n_2714),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2849),
.A2(n_2763),
.B(n_2714),
.Y(n_2874)
);

OA21x2_ASAP7_75t_L g2875 ( 
.A1(n_2849),
.A2(n_2766),
.B(n_2762),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2841),
.B(n_2801),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2833),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2817),
.Y(n_2878)
);

NAND4xp25_ASAP7_75t_L g2879 ( 
.A(n_2848),
.B(n_2807),
.C(n_2723),
.D(n_2693),
.Y(n_2879)
);

OAI211xp5_ASAP7_75t_SL g2880 ( 
.A1(n_2840),
.A2(n_2848),
.B(n_2829),
.C(n_2834),
.Y(n_2880)
);

BUFx3_ASAP7_75t_L g2881 ( 
.A(n_2844),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2841),
.B(n_2812),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2820),
.Y(n_2883)
);

AO21x2_ASAP7_75t_L g2884 ( 
.A1(n_2843),
.A2(n_2762),
.B(n_2761),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2839),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2844),
.B(n_2814),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2856),
.B(n_2812),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2825),
.Y(n_2888)
);

OA21x2_ASAP7_75t_L g2889 ( 
.A1(n_2824),
.A2(n_2766),
.B(n_2777),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2854),
.B(n_2808),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2823),
.A2(n_2763),
.B1(n_2689),
.B2(n_2704),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2863),
.B(n_2855),
.Y(n_2892)
);

OAI21xp5_ASAP7_75t_L g2893 ( 
.A1(n_2874),
.A2(n_2827),
.B(n_2823),
.Y(n_2893)
);

OR2x2_ASAP7_75t_L g2894 ( 
.A(n_2864),
.B(n_2852),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2866),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2876),
.B(n_2827),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2862),
.B(n_2853),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2859),
.Y(n_2898)
);

INVx3_ASAP7_75t_SL g2899 ( 
.A(n_2876),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2882),
.B(n_2832),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2869),
.Y(n_2901)
);

INVxp67_ASAP7_75t_SL g2902 ( 
.A(n_2886),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2860),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_L g2904 ( 
.A(n_2886),
.B(n_2672),
.Y(n_2904)
);

AND2x4_ASAP7_75t_SL g2905 ( 
.A(n_2868),
.B(n_2666),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2858),
.B(n_2853),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2861),
.Y(n_2907)
);

NAND2x1p5_ASAP7_75t_L g2908 ( 
.A(n_2881),
.B(n_2666),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2881),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2877),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2878),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2890),
.B(n_2831),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2872),
.B(n_2843),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2861),
.B(n_2831),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2867),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2883),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2870),
.B(n_2847),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2885),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2872),
.B(n_2847),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2867),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2865),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2873),
.B(n_2842),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2873),
.B(n_2824),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2874),
.B(n_2835),
.Y(n_2924)
);

OAI22xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2857),
.A2(n_2835),
.B1(n_2850),
.B2(n_2744),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2887),
.B(n_2808),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2888),
.B(n_2809),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2884),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2871),
.B(n_2850),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2891),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2884),
.B(n_2809),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2889),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2875),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2889),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2875),
.Y(n_2935)
);

AND3x2_ASAP7_75t_L g2936 ( 
.A(n_2857),
.B(n_2753),
.C(n_2732),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2875),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2909),
.Y(n_2938)
);

OR2x2_ASAP7_75t_L g2939 ( 
.A(n_2906),
.B(n_2879),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2933),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2933),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2892),
.B(n_2891),
.Y(n_2942)
);

OR2x2_ASAP7_75t_L g2943 ( 
.A(n_2894),
.B(n_2724),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2936),
.B(n_2799),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2909),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2911),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2903),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2899),
.B(n_2880),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2911),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2916),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2916),
.Y(n_2951)
);

INVxp67_ASAP7_75t_L g2952 ( 
.A(n_2902),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2918),
.Y(n_2953)
);

OR2x2_ASAP7_75t_L g2954 ( 
.A(n_2917),
.B(n_2880),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2910),
.B(n_2889),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2896),
.B(n_2677),
.Y(n_2956)
);

INVx3_ASAP7_75t_L g2957 ( 
.A(n_2896),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2918),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2898),
.B(n_2806),
.Y(n_2959)
);

NAND2xp33_ASAP7_75t_L g2960 ( 
.A(n_2908),
.B(n_2693),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2907),
.B(n_2811),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2935),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2903),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2912),
.B(n_2730),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2915),
.B(n_2773),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2897),
.B(n_2773),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2900),
.B(n_2715),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2904),
.B(n_2668),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2905),
.B(n_2704),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2926),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2935),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_L g2972 ( 
.A(n_2930),
.B(n_2671),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2914),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2914),
.B(n_2683),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2937),
.Y(n_2975)
);

AND2x4_ASAP7_75t_L g2976 ( 
.A(n_2901),
.B(n_2718),
.Y(n_2976)
);

INVx1_ASAP7_75t_SL g2977 ( 
.A(n_2929),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2927),
.B(n_2683),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2921),
.B(n_2920),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2895),
.B(n_2681),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2895),
.B(n_2686),
.Y(n_2981)
);

AOI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2913),
.A2(n_2692),
.B1(n_2721),
.B2(n_2725),
.Y(n_2982)
);

OR2x2_ASAP7_75t_L g2983 ( 
.A(n_2922),
.B(n_2695),
.Y(n_2983)
);

INVx3_ASAP7_75t_L g2984 ( 
.A(n_2931),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2923),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2932),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2919),
.A2(n_2692),
.B1(n_2675),
.B2(n_2682),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2893),
.B(n_84),
.Y(n_2988)
);

INVx2_ASAP7_75t_SL g2989 ( 
.A(n_2928),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2925),
.B(n_2924),
.Y(n_2990)
);

OR2x2_ASAP7_75t_L g2991 ( 
.A(n_2937),
.B(n_2934),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2906),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2909),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2906),
.Y(n_2994)
);

OR2x2_ASAP7_75t_L g2995 ( 
.A(n_2906),
.B(n_2695),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2899),
.B(n_84),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2906),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2909),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2909),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2933),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2899),
.B(n_85),
.Y(n_3001)
);

NOR2xp33_ASAP7_75t_L g3002 ( 
.A(n_2899),
.B(n_86),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2909),
.Y(n_3003)
);

OR2x2_ASAP7_75t_L g3004 ( 
.A(n_2906),
.B(n_2695),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2957),
.B(n_88),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2991),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2957),
.B(n_88),
.Y(n_3007)
);

OR2x2_ASAP7_75t_L g3008 ( 
.A(n_2952),
.B(n_89),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2996),
.B(n_91),
.Y(n_3009)
);

NAND2xp33_ASAP7_75t_SL g3010 ( 
.A(n_2954),
.B(n_91),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_3001),
.B(n_92),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2940),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2940),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2941),
.Y(n_3014)
);

INVxp67_ASAP7_75t_SL g3015 ( 
.A(n_3002),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2985),
.B(n_92),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2973),
.B(n_93),
.Y(n_3017)
);

NAND4xp25_ASAP7_75t_L g3018 ( 
.A(n_2948),
.B(n_2945),
.C(n_2993),
.D(n_2938),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2941),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2998),
.B(n_94),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2970),
.B(n_94),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2999),
.B(n_95),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2962),
.Y(n_3023)
);

NAND2x1p5_ASAP7_75t_L g3024 ( 
.A(n_2988),
.B(n_96),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2977),
.B(n_96),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2962),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_3003),
.B(n_97),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2971),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2992),
.B(n_2994),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2947),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2971),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2968),
.B(n_2963),
.Y(n_3032)
);

CKINVDCx16_ASAP7_75t_R g3033 ( 
.A(n_2939),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2997),
.B(n_97),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2975),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2975),
.Y(n_3036)
);

OR2x2_ASAP7_75t_L g3037 ( 
.A(n_2942),
.B(n_99),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2956),
.B(n_100),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2944),
.B(n_2969),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_3000),
.Y(n_3040)
);

NAND2x1p5_ASAP7_75t_L g3041 ( 
.A(n_2979),
.B(n_2984),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2974),
.Y(n_3042)
);

BUFx2_ASAP7_75t_L g3043 ( 
.A(n_2984),
.Y(n_3043)
);

INVx5_ASAP7_75t_L g3044 ( 
.A(n_2989),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2978),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2964),
.B(n_101),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2967),
.B(n_101),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_3000),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2980),
.B(n_103),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2986),
.Y(n_3050)
);

OR2x6_ASAP7_75t_L g3051 ( 
.A(n_2990),
.B(n_104),
.Y(n_3051)
);

INVxp67_ASAP7_75t_L g3052 ( 
.A(n_2983),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2946),
.B(n_104),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2949),
.B(n_105),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2960),
.B(n_105),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2950),
.B(n_106),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2951),
.B(n_109),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2953),
.B(n_111),
.Y(n_3058)
);

NAND2xp33_ASAP7_75t_R g3059 ( 
.A(n_2955),
.B(n_111),
.Y(n_3059)
);

INVx5_ASAP7_75t_L g3060 ( 
.A(n_2976),
.Y(n_3060)
);

OR2x2_ASAP7_75t_L g3061 ( 
.A(n_2959),
.B(n_112),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_2943),
.B(n_112),
.Y(n_3062)
);

BUFx3_ASAP7_75t_L g3063 ( 
.A(n_2958),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2981),
.B(n_2976),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2961),
.B(n_113),
.Y(n_3065)
);

INVxp67_ASAP7_75t_L g3066 ( 
.A(n_2972),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2966),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2981),
.B(n_2982),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2995),
.B(n_115),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3004),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2965),
.Y(n_3071)
);

OR2x2_ASAP7_75t_L g3072 ( 
.A(n_2987),
.B(n_117),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2957),
.B(n_117),
.Y(n_3073)
);

INVx1_ASAP7_75t_SL g3074 ( 
.A(n_2996),
.Y(n_3074)
);

BUFx3_ASAP7_75t_L g3075 ( 
.A(n_2996),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2991),
.Y(n_3076)
);

INVx5_ASAP7_75t_L g3077 ( 
.A(n_2996),
.Y(n_3077)
);

OR2x2_ASAP7_75t_L g3078 ( 
.A(n_2952),
.B(n_119),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2957),
.Y(n_3079)
);

NOR3xp33_ASAP7_75t_L g3080 ( 
.A(n_2990),
.B(n_2690),
.C(n_2678),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2957),
.Y(n_3081)
);

NAND4xp75_ASAP7_75t_L g3082 ( 
.A(n_2990),
.B(n_121),
.C(n_119),
.D(n_120),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2952),
.B(n_122),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2996),
.B(n_124),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2996),
.B(n_124),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2996),
.B(n_125),
.Y(n_3086)
);

NOR2x1_ASAP7_75t_SL g3087 ( 
.A(n_2996),
.B(n_125),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2952),
.B(n_126),
.Y(n_3088)
);

INVx3_ASAP7_75t_L g3089 ( 
.A(n_2957),
.Y(n_3089)
);

INVx1_ASAP7_75t_SL g3090 ( 
.A(n_2996),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2991),
.Y(n_3091)
);

OR2x2_ASAP7_75t_L g3092 ( 
.A(n_2952),
.B(n_126),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2990),
.A2(n_127),
.B(n_128),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2957),
.B(n_128),
.Y(n_3094)
);

NOR4xp25_ASAP7_75t_SL g3095 ( 
.A(n_2985),
.B(n_135),
.C(n_129),
.D(n_131),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2957),
.B(n_131),
.Y(n_3096)
);

O2A1O1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2985),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_3097)
);

NAND2x1_ASAP7_75t_SL g3098 ( 
.A(n_3089),
.B(n_136),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3079),
.B(n_139),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3043),
.Y(n_3100)
);

OR2x2_ASAP7_75t_L g3101 ( 
.A(n_3033),
.B(n_139),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3054),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_3077),
.Y(n_3103)
);

INVx1_ASAP7_75t_SL g3104 ( 
.A(n_3074),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3057),
.Y(n_3105)
);

OR2x2_ASAP7_75t_L g3106 ( 
.A(n_3006),
.B(n_140),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_3090),
.B(n_140),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_3081),
.B(n_142),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3047),
.B(n_142),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3058),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3087),
.B(n_143),
.Y(n_3111)
);

AND2x4_ASAP7_75t_L g3112 ( 
.A(n_3077),
.B(n_144),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3034),
.Y(n_3113)
);

NAND4xp25_ASAP7_75t_SL g3114 ( 
.A(n_3029),
.B(n_148),
.C(n_146),
.D(n_147),
.Y(n_3114)
);

INVx1_ASAP7_75t_SL g3115 ( 
.A(n_3077),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3037),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_3041),
.B(n_3032),
.Y(n_3117)
);

OR2x2_ASAP7_75t_L g3118 ( 
.A(n_3076),
.B(n_147),
.Y(n_3118)
);

NAND3xp33_ASAP7_75t_L g3119 ( 
.A(n_3010),
.B(n_3059),
.C(n_3093),
.Y(n_3119)
);

OAI33xp33_ASAP7_75t_L g3120 ( 
.A1(n_3050),
.A2(n_3091),
.A3(n_3018),
.B1(n_3012),
.B2(n_3019),
.B3(n_3013),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_3030),
.B(n_148),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_3055),
.B(n_150),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_3009),
.B(n_3005),
.Y(n_3123)
);

AND2x4_ASAP7_75t_L g3124 ( 
.A(n_3075),
.B(n_150),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3025),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_3007),
.B(n_152),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3011),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_3024),
.B(n_152),
.Y(n_3128)
);

AND2x4_ASAP7_75t_L g3129 ( 
.A(n_3073),
.B(n_153),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_3038),
.B(n_154),
.Y(n_3130)
);

INVxp67_ASAP7_75t_L g3131 ( 
.A(n_3051),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_3049),
.B(n_156),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_3094),
.B(n_156),
.Y(n_3133)
);

OR3x2_ASAP7_75t_L g3134 ( 
.A(n_3062),
.B(n_3061),
.C(n_3008),
.Y(n_3134)
);

INVxp67_ASAP7_75t_L g3135 ( 
.A(n_3051),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3069),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3078),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3092),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_3039),
.B(n_157),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3016),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3096),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_3060),
.B(n_157),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_3022),
.B(n_158),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3014),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_3066),
.B(n_159),
.Y(n_3145)
);

NAND4xp25_ASAP7_75t_SL g3146 ( 
.A(n_3042),
.B(n_162),
.C(n_160),
.D(n_161),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3023),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_3015),
.B(n_160),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_3017),
.B(n_161),
.Y(n_3149)
);

AOI31xp33_ASAP7_75t_SL g3150 ( 
.A1(n_3045),
.A2(n_165),
.A3(n_163),
.B(n_164),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3026),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3046),
.B(n_166),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3028),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3031),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3060),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3035),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_3063),
.B(n_166),
.Y(n_3157)
);

OAI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3044),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3158)
);

BUFx3_ASAP7_75t_L g3159 ( 
.A(n_3084),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3036),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_3020),
.B(n_167),
.Y(n_3161)
);

CKINVDCx16_ASAP7_75t_R g3162 ( 
.A(n_3095),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3067),
.B(n_169),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3060),
.B(n_171),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3044),
.B(n_172),
.Y(n_3165)
);

HB1xp67_ASAP7_75t_L g3166 ( 
.A(n_3044),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3040),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3083),
.B(n_174),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3048),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_3088),
.B(n_174),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3064),
.B(n_175),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_3027),
.B(n_176),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3085),
.B(n_176),
.Y(n_3173)
);

NOR2x1_ASAP7_75t_L g3174 ( 
.A(n_3021),
.B(n_177),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_3086),
.B(n_177),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3082),
.B(n_178),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3065),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3071),
.B(n_180),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3053),
.B(n_181),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3056),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_3068),
.B(n_182),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_3097),
.B(n_182),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_3052),
.B(n_183),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3070),
.Y(n_3184)
);

NAND2x1p5_ASAP7_75t_L g3185 ( 
.A(n_3072),
.B(n_183),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_3080),
.B(n_185),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3089),
.B(n_185),
.Y(n_3187)
);

INVxp67_ASAP7_75t_SL g3188 ( 
.A(n_3087),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3043),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3089),
.B(n_186),
.Y(n_3190)
);

OR2x2_ASAP7_75t_L g3191 ( 
.A(n_3033),
.B(n_186),
.Y(n_3191)
);

INVx1_ASAP7_75t_SL g3192 ( 
.A(n_3074),
.Y(n_3192)
);

OAI21xp33_ASAP7_75t_L g3193 ( 
.A1(n_3075),
.A2(n_188),
.B(n_189),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3043),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_3087),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3089),
.B(n_188),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3089),
.B(n_189),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_SL g3198 ( 
.A(n_3074),
.B(n_190),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3074),
.B(n_190),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3010),
.A2(n_191),
.B(n_192),
.Y(n_3200)
);

AND2x2_ASAP7_75t_L g3201 ( 
.A(n_3089),
.B(n_192),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_3087),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3074),
.B(n_193),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3074),
.B(n_193),
.Y(n_3204)
);

NOR2x1_ASAP7_75t_L g3205 ( 
.A(n_3089),
.B(n_195),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_3077),
.B(n_195),
.Y(n_3206)
);

INVxp67_ASAP7_75t_L g3207 ( 
.A(n_3087),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3074),
.B(n_196),
.Y(n_3208)
);

HB1xp67_ASAP7_75t_L g3209 ( 
.A(n_3077),
.Y(n_3209)
);

NOR2x1_ASAP7_75t_L g3210 ( 
.A(n_3089),
.B(n_196),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3043),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3043),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_3087),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3033),
.B(n_197),
.Y(n_3214)
);

HB1xp67_ASAP7_75t_L g3215 ( 
.A(n_3077),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3043),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3043),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3033),
.B(n_198),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_3087),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3043),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3074),
.B(n_199),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3043),
.Y(n_3222)
);

NAND2x1p5_ASAP7_75t_L g3223 ( 
.A(n_3077),
.B(n_199),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3077),
.B(n_200),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3074),
.B(n_202),
.Y(n_3225)
);

NAND3xp33_ASAP7_75t_SL g3226 ( 
.A(n_3093),
.B(n_205),
.C(n_206),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3074),
.B(n_208),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3074),
.B(n_209),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3087),
.Y(n_3229)
);

NAND3xp33_ASAP7_75t_L g3230 ( 
.A(n_3010),
.B(n_209),
.C(n_210),
.Y(n_3230)
);

OR2x2_ASAP7_75t_L g3231 ( 
.A(n_3033),
.B(n_210),
.Y(n_3231)
);

INVx2_ASAP7_75t_SL g3232 ( 
.A(n_3077),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_3010),
.A2(n_212),
.B(n_213),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3074),
.B(n_212),
.Y(n_3234)
);

INVx1_ASAP7_75t_SL g3235 ( 
.A(n_3074),
.Y(n_3235)
);

AND2x2_ASAP7_75t_SL g3236 ( 
.A(n_3033),
.B(n_215),
.Y(n_3236)
);

OAI221xp5_ASAP7_75t_L g3237 ( 
.A1(n_3010),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_221),
.Y(n_3237)
);

INVx2_ASAP7_75t_SL g3238 ( 
.A(n_3077),
.Y(n_3238)
);

OR2x2_ASAP7_75t_L g3239 ( 
.A(n_3033),
.B(n_217),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3074),
.B(n_219),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_3089),
.B(n_221),
.Y(n_3241)
);

INVx1_ASAP7_75t_SL g3242 ( 
.A(n_3074),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_3077),
.B(n_222),
.Y(n_3243)
);

INVx1_ASAP7_75t_SL g3244 ( 
.A(n_3074),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3074),
.B(n_223),
.Y(n_3245)
);

NAND3xp33_ASAP7_75t_L g3246 ( 
.A(n_3010),
.B(n_224),
.C(n_225),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3074),
.B(n_224),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3043),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3089),
.B(n_225),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3077),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3087),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3074),
.B(n_226),
.Y(n_3252)
);

INVx1_ASAP7_75t_SL g3253 ( 
.A(n_3074),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3243),
.A2(n_3142),
.B(n_3236),
.Y(n_3254)
);

OAI221xp5_ASAP7_75t_L g3255 ( 
.A1(n_3207),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.C(n_230),
.Y(n_3255)
);

AOI31xp33_ASAP7_75t_SL g3256 ( 
.A1(n_3195),
.A2(n_230),
.A3(n_228),
.B(n_229),
.Y(n_3256)
);

OAI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3162),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3257)
);

NAND3x1_ASAP7_75t_L g3258 ( 
.A(n_3117),
.B(n_232),
.C(n_236),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3129),
.B(n_236),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3104),
.B(n_237),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3101),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3191),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3192),
.B(n_237),
.Y(n_3263)
);

HB1xp67_ASAP7_75t_L g3264 ( 
.A(n_3103),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3214),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3235),
.B(n_238),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_SL g3267 ( 
.A1(n_3119),
.A2(n_3188),
.B1(n_3213),
.B2(n_3202),
.Y(n_3267)
);

OA21x2_ASAP7_75t_L g3268 ( 
.A1(n_3165),
.A2(n_238),
.B(n_239),
.Y(n_3268)
);

OAI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_3198),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3218),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_3098),
.B(n_240),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3242),
.B(n_241),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3219),
.A2(n_246),
.B1(n_243),
.B2(n_244),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3231),
.Y(n_3274)
);

INVx1_ASAP7_75t_SL g3275 ( 
.A(n_3239),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3121),
.Y(n_3276)
);

INVx2_ASAP7_75t_SL g3277 ( 
.A(n_3223),
.Y(n_3277)
);

AOI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3229),
.A2(n_247),
.B1(n_243),
.B2(n_246),
.Y(n_3278)
);

NAND2x1p5_ASAP7_75t_L g3279 ( 
.A(n_3157),
.B(n_248),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3134),
.Y(n_3280)
);

INVxp67_ASAP7_75t_L g3281 ( 
.A(n_3209),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3129),
.B(n_249),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3133),
.B(n_250),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3244),
.B(n_250),
.Y(n_3284)
);

OAI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_3205),
.A2(n_251),
.B(n_253),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3215),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3250),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3133),
.B(n_254),
.Y(n_3288)
);

AOI222xp33_ASAP7_75t_L g3289 ( 
.A1(n_3181),
.A2(n_257),
.B1(n_259),
.B2(n_255),
.C1(n_256),
.C2(n_258),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3132),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_3251),
.B(n_255),
.Y(n_3291)
);

AOI222xp33_ASAP7_75t_L g3292 ( 
.A1(n_3131),
.A2(n_259),
.B1(n_261),
.B2(n_257),
.C1(n_258),
.C2(n_260),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3130),
.B(n_261),
.Y(n_3293)
);

INVxp67_ASAP7_75t_L g3294 ( 
.A(n_3166),
.Y(n_3294)
);

AOI21xp33_ASAP7_75t_L g3295 ( 
.A1(n_3135),
.A2(n_263),
.B(n_264),
.Y(n_3295)
);

INVx1_ASAP7_75t_SL g3296 ( 
.A(n_3253),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3112),
.B(n_265),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3185),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3159),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3127),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3112),
.B(n_267),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3224),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_3100),
.B(n_268),
.Y(n_3303)
);

AOI22xp5_ASAP7_75t_L g3304 ( 
.A1(n_3226),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3189),
.B(n_3194),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3224),
.B(n_269),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_3211),
.B(n_270),
.Y(n_3307)
);

CKINVDCx14_ASAP7_75t_R g3308 ( 
.A(n_3141),
.Y(n_3308)
);

OAI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_3115),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_3309)
);

NOR2x1_ASAP7_75t_L g3310 ( 
.A(n_3206),
.B(n_272),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_3210),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3124),
.B(n_3143),
.Y(n_3312)
);

INVxp67_ASAP7_75t_L g3313 ( 
.A(n_3128),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3124),
.B(n_273),
.Y(n_3314)
);

OAI21xp5_ASAP7_75t_L g3315 ( 
.A1(n_3200),
.A2(n_3233),
.B(n_3230),
.Y(n_3315)
);

OAI32xp33_ASAP7_75t_L g3316 ( 
.A1(n_3212),
.A2(n_276),
.A3(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_3114),
.B(n_274),
.Y(n_3317)
);

O2A1O1Ixp33_ASAP7_75t_L g3318 ( 
.A1(n_3150),
.A2(n_278),
.B(n_275),
.C(n_276),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3106),
.Y(n_3319)
);

NAND3xp33_ASAP7_75t_L g3320 ( 
.A(n_3216),
.B(n_278),
.C(n_279),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3116),
.B(n_280),
.Y(n_3321)
);

AOI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3125),
.A2(n_3136),
.B1(n_3113),
.B2(n_3182),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3118),
.Y(n_3323)
);

AOI211xp5_ASAP7_75t_L g3324 ( 
.A1(n_3232),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3152),
.Y(n_3325)
);

BUFx3_ASAP7_75t_L g3326 ( 
.A(n_3099),
.Y(n_3326)
);

AOI21xp33_ASAP7_75t_SL g3327 ( 
.A1(n_3238),
.A2(n_282),
.B(n_283),
.Y(n_3327)
);

AOI221xp5_ASAP7_75t_L g3328 ( 
.A1(n_3120),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.C(n_287),
.Y(n_3328)
);

AOI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_3177),
.A2(n_288),
.B1(n_285),
.B2(n_286),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3140),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_3330)
);

OAI22xp5_ASAP7_75t_L g3331 ( 
.A1(n_3217),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3174),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_3332)
);

HB1xp67_ASAP7_75t_L g3333 ( 
.A(n_3164),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3108),
.B(n_295),
.Y(n_3334)
);

OAI22xp5_ASAP7_75t_L g3335 ( 
.A1(n_3220),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3109),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_3111),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3123),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3173),
.Y(n_3339)
);

NAND2x1_ASAP7_75t_L g3340 ( 
.A(n_3155),
.B(n_298),
.Y(n_3340)
);

OAI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3246),
.A2(n_299),
.B(n_300),
.Y(n_3341)
);

NOR2xp33_ASAP7_75t_L g3342 ( 
.A(n_3146),
.B(n_300),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3102),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3105),
.B(n_301),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3110),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3345)
);

XNOR2xp5_ASAP7_75t_L g3346 ( 
.A(n_3139),
.B(n_302),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3149),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3172),
.B(n_303),
.Y(n_3348)
);

AOI21xp33_ASAP7_75t_SL g3349 ( 
.A1(n_3222),
.A2(n_304),
.B(n_305),
.Y(n_3349)
);

OR2x2_ASAP7_75t_L g3350 ( 
.A(n_3248),
.B(n_305),
.Y(n_3350)
);

AOI321xp33_ASAP7_75t_SL g3351 ( 
.A1(n_3183),
.A2(n_306),
.A3(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_3351)
);

OR2x2_ASAP7_75t_L g3352 ( 
.A(n_3107),
.B(n_307),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3148),
.Y(n_3353)
);

INVxp67_ASAP7_75t_L g3354 ( 
.A(n_3175),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3126),
.Y(n_3355)
);

XNOR2xp5_ASAP7_75t_L g3356 ( 
.A(n_3158),
.B(n_308),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3176),
.A2(n_3203),
.B(n_3199),
.Y(n_3357)
);

OAI21xp33_ASAP7_75t_L g3358 ( 
.A1(n_3180),
.A2(n_310),
.B(n_311),
.Y(n_3358)
);

NAND3xp33_ASAP7_75t_L g3359 ( 
.A(n_3186),
.B(n_312),
.C(n_313),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3187),
.B(n_312),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3179),
.Y(n_3361)
);

AOI221xp5_ASAP7_75t_L g3362 ( 
.A1(n_3184),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.C(n_316),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3190),
.Y(n_3363)
);

OR2x2_ASAP7_75t_L g3364 ( 
.A(n_3204),
.B(n_315),
.Y(n_3364)
);

AOI221xp5_ASAP7_75t_L g3365 ( 
.A1(n_3137),
.A2(n_3138),
.B1(n_3163),
.B2(n_3144),
.C(n_3151),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3208),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3193),
.A2(n_320),
.B1(n_317),
.B2(n_318),
.Y(n_3367)
);

OAI21x1_ASAP7_75t_L g3368 ( 
.A1(n_3221),
.A2(n_3227),
.B(n_3225),
.Y(n_3368)
);

AOI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3122),
.A2(n_326),
.B1(n_322),
.B2(n_324),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3228),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3234),
.A2(n_3245),
.B1(n_3247),
.B2(n_3240),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_3196),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3171),
.A2(n_327),
.B1(n_322),
.B2(n_324),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3252),
.Y(n_3374)
);

A2O1A1Ixp33_ASAP7_75t_L g3375 ( 
.A1(n_3237),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3197),
.B(n_3201),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3145),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3296),
.B(n_3241),
.Y(n_3378)
);

NAND2x1p5_ASAP7_75t_L g3379 ( 
.A(n_3340),
.B(n_3277),
.Y(n_3379)
);

AND3x1_ASAP7_75t_L g3380 ( 
.A(n_3328),
.B(n_3249),
.C(n_3153),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3271),
.B(n_3161),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3333),
.Y(n_3382)
);

AOI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3275),
.A2(n_3178),
.B1(n_3170),
.B2(n_3168),
.Y(n_3383)
);

OR2x2_ASAP7_75t_L g3384 ( 
.A(n_3299),
.B(n_3147),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3260),
.B(n_3154),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3279),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3372),
.B(n_3156),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3350),
.B(n_3160),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3264),
.Y(n_3389)
);

OAI21xp33_ASAP7_75t_L g3390 ( 
.A1(n_3267),
.A2(n_3169),
.B(n_3167),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3293),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3268),
.Y(n_3392)
);

OR2x2_ASAP7_75t_L g3393 ( 
.A(n_3300),
.B(n_328),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3258),
.Y(n_3394)
);

INVx1_ASAP7_75t_SL g3395 ( 
.A(n_3312),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3311),
.B(n_330),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3263),
.B(n_332),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_3266),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3268),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3290),
.B(n_332),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3348),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3272),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3326),
.Y(n_3403)
);

INVxp67_ASAP7_75t_L g3404 ( 
.A(n_3310),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3254),
.B(n_333),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3284),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_L g3407 ( 
.A(n_3327),
.B(n_335),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3308),
.B(n_335),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3302),
.B(n_336),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3305),
.B(n_3303),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3307),
.B(n_338),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3310),
.Y(n_3412)
);

OR2x2_ASAP7_75t_L g3413 ( 
.A(n_3343),
.B(n_338),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3349),
.B(n_339),
.Y(n_3414)
);

HB1xp67_ASAP7_75t_L g3415 ( 
.A(n_3346),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3259),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3282),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3361),
.B(n_340),
.Y(n_3418)
);

INVxp67_ASAP7_75t_SL g3419 ( 
.A(n_3376),
.Y(n_3419)
);

O2A1O1Ixp5_ASAP7_75t_L g3420 ( 
.A1(n_3286),
.A2(n_343),
.B(n_340),
.C(n_341),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3294),
.B(n_343),
.Y(n_3421)
);

INVx1_ASAP7_75t_SL g3422 ( 
.A(n_3352),
.Y(n_3422)
);

INVxp67_ASAP7_75t_L g3423 ( 
.A(n_3342),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3364),
.Y(n_3424)
);

NOR2x1_ASAP7_75t_L g3425 ( 
.A(n_3320),
.B(n_344),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3281),
.B(n_344),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3283),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3288),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3297),
.Y(n_3429)
);

INVx2_ASAP7_75t_SL g3430 ( 
.A(n_3291),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3261),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3298),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3289),
.B(n_345),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3301),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3262),
.B(n_346),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3265),
.B(n_347),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3306),
.Y(n_3437)
);

AND2x4_ASAP7_75t_SL g3438 ( 
.A(n_3363),
.B(n_347),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3334),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3270),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3274),
.B(n_348),
.Y(n_3441)
);

INVx1_ASAP7_75t_SL g3442 ( 
.A(n_3360),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3287),
.B(n_348),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3365),
.B(n_349),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3276),
.B(n_349),
.Y(n_3445)
);

BUFx12f_ASAP7_75t_L g3446 ( 
.A(n_3313),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3354),
.B(n_350),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3318),
.B(n_350),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3314),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3319),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3323),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_SL g3452 ( 
.A(n_3317),
.B(n_351),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3377),
.B(n_351),
.Y(n_3453)
);

OR2x2_ASAP7_75t_L g3454 ( 
.A(n_3344),
.B(n_3321),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3337),
.A2(n_356),
.B1(n_352),
.B2(n_353),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3324),
.B(n_353),
.Y(n_3456)
);

INVx1_ASAP7_75t_SL g3457 ( 
.A(n_3280),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3257),
.B(n_357),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3269),
.B(n_358),
.Y(n_3459)
);

INVx1_ASAP7_75t_SL g3460 ( 
.A(n_3356),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3256),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3292),
.B(n_359),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3347),
.Y(n_3463)
);

HB1xp67_ASAP7_75t_L g3464 ( 
.A(n_3285),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3315),
.B(n_359),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3368),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3341),
.B(n_360),
.Y(n_3467)
);

HB1xp67_ASAP7_75t_L g3468 ( 
.A(n_3309),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_3331),
.B(n_360),
.Y(n_3469)
);

HB1xp67_ASAP7_75t_L g3470 ( 
.A(n_3325),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_3336),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3355),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3339),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3304),
.B(n_3332),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3353),
.Y(n_3475)
);

INVx2_ASAP7_75t_SL g3476 ( 
.A(n_3335),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3273),
.B(n_363),
.Y(n_3477)
);

OR2x2_ASAP7_75t_L g3478 ( 
.A(n_3322),
.B(n_363),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3370),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3374),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3373),
.B(n_3357),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3338),
.Y(n_3482)
);

OR2x2_ASAP7_75t_L g3483 ( 
.A(n_3358),
.B(n_364),
.Y(n_3483)
);

OR2x2_ASAP7_75t_L g3484 ( 
.A(n_3366),
.B(n_364),
.Y(n_3484)
);

O2A1O1Ixp5_ASAP7_75t_L g3485 ( 
.A1(n_3371),
.A2(n_368),
.B(n_365),
.C(n_367),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3369),
.B(n_365),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3278),
.B(n_367),
.Y(n_3487)
);

HB1xp67_ASAP7_75t_L g3488 ( 
.A(n_3255),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3367),
.B(n_368),
.Y(n_3489)
);

NAND2x1p5_ASAP7_75t_L g3490 ( 
.A(n_3345),
.B(n_370),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3375),
.B(n_370),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3329),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3316),
.Y(n_3493)
);

INVxp67_ASAP7_75t_L g3494 ( 
.A(n_3359),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3330),
.B(n_371),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3362),
.B(n_372),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3295),
.B(n_3351),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3271),
.B(n_372),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3296),
.B(n_373),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3296),
.B(n_373),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3271),
.B(n_375),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3271),
.B(n_376),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3296),
.B(n_378),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3279),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3333),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_3296),
.B(n_378),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3333),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3296),
.B(n_379),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3271),
.B(n_379),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3271),
.B(n_380),
.Y(n_3510)
);

INVx3_ASAP7_75t_L g3511 ( 
.A(n_3340),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3271),
.B(n_381),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3271),
.B(n_381),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3333),
.Y(n_3514)
);

OAI21xp33_ASAP7_75t_L g3515 ( 
.A1(n_3296),
.A2(n_382),
.B(n_383),
.Y(n_3515)
);

INVx2_ASAP7_75t_SL g3516 ( 
.A(n_3260),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3271),
.B(n_382),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_SL g3518 ( 
.A(n_3296),
.B(n_383),
.Y(n_3518)
);

INVx3_ASAP7_75t_SL g3519 ( 
.A(n_3296),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3271),
.B(n_384),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3333),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3296),
.B(n_385),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3333),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3333),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3271),
.B(n_386),
.Y(n_3525)
);

INVx1_ASAP7_75t_SL g3526 ( 
.A(n_3296),
.Y(n_3526)
);

INVxp67_ASAP7_75t_L g3527 ( 
.A(n_3311),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3271),
.B(n_386),
.Y(n_3528)
);

NOR2xp67_ASAP7_75t_L g3529 ( 
.A(n_3277),
.B(n_387),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3271),
.B(n_389),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3318),
.A2(n_389),
.B(n_390),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3279),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3379),
.Y(n_3533)
);

AOI311xp33_ASAP7_75t_L g3534 ( 
.A1(n_3389),
.A2(n_391),
.A3(n_392),
.B(n_393),
.C(n_394),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3519),
.B(n_392),
.Y(n_3535)
);

AOI21xp33_ASAP7_75t_L g3536 ( 
.A1(n_3404),
.A2(n_3399),
.B(n_3392),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3410),
.B(n_393),
.Y(n_3537)
);

NOR3xp33_ASAP7_75t_SL g3538 ( 
.A(n_3390),
.B(n_394),
.C(n_395),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3526),
.B(n_396),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3398),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3511),
.B(n_396),
.Y(n_3541)
);

INVxp67_ASAP7_75t_L g3542 ( 
.A(n_3518),
.Y(n_3542)
);

OAI21xp33_ASAP7_75t_SL g3543 ( 
.A1(n_3378),
.A2(n_397),
.B(n_399),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3408),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3415),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3499),
.B(n_3500),
.Y(n_3546)
);

OAI311xp33_ASAP7_75t_L g3547 ( 
.A1(n_3527),
.A2(n_397),
.A3(n_399),
.B1(n_400),
.C1(n_401),
.Y(n_3547)
);

OAI221xp5_ASAP7_75t_L g3548 ( 
.A1(n_3505),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.C(n_405),
.Y(n_3548)
);

INVxp67_ASAP7_75t_SL g3549 ( 
.A(n_3511),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3461),
.B(n_3395),
.Y(n_3550)
);

HB1xp67_ASAP7_75t_L g3551 ( 
.A(n_3461),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3412),
.Y(n_3552)
);

INVx1_ASAP7_75t_SL g3553 ( 
.A(n_3411),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3516),
.B(n_402),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3446),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_3403),
.B(n_405),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3397),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3503),
.B(n_406),
.Y(n_3558)
);

INVx1_ASAP7_75t_SL g3559 ( 
.A(n_3508),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3394),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3522),
.B(n_407),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3385),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3388),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3453),
.Y(n_3564)
);

NOR2xp67_ASAP7_75t_SL g3565 ( 
.A(n_3470),
.B(n_3505),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3529),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3445),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3393),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3438),
.Y(n_3569)
);

NOR3xp33_ASAP7_75t_SL g3570 ( 
.A(n_3387),
.B(n_407),
.C(n_408),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_3386),
.B(n_408),
.Y(n_3571)
);

AOI221xp5_ASAP7_75t_L g3572 ( 
.A1(n_3380),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.C(n_414),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3413),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3419),
.B(n_410),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3443),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3465),
.Y(n_3576)
);

NAND4xp25_ASAP7_75t_L g3577 ( 
.A(n_3382),
.B(n_415),
.C(n_411),
.D(n_414),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3468),
.Y(n_3578)
);

XOR2xp5_ASAP7_75t_L g3579 ( 
.A(n_3383),
.B(n_415),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3464),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3504),
.B(n_416),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3532),
.B(n_417),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3454),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3430),
.B(n_417),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3448),
.Y(n_3585)
);

NOR2xp67_ASAP7_75t_L g3586 ( 
.A(n_3507),
.B(n_418),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3402),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3406),
.B(n_419),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3514),
.B(n_420),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3422),
.B(n_420),
.Y(n_3590)
);

AOI21xp33_ASAP7_75t_L g3591 ( 
.A1(n_3457),
.A2(n_421),
.B(n_422),
.Y(n_3591)
);

OAI211xp5_ASAP7_75t_L g3592 ( 
.A1(n_3521),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3466),
.A2(n_427),
.B1(n_424),
.B2(n_426),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3424),
.B(n_426),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3433),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3407),
.B(n_427),
.Y(n_3596)
);

INVx2_ASAP7_75t_SL g3597 ( 
.A(n_3384),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3531),
.B(n_429),
.Y(n_3598)
);

AOI221xp5_ASAP7_75t_L g3599 ( 
.A1(n_3497),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.C(n_433),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3414),
.B(n_430),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3442),
.B(n_431),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3523),
.B(n_432),
.Y(n_3602)
);

NOR4xp25_ASAP7_75t_SL g3603 ( 
.A(n_3431),
.B(n_435),
.C(n_433),
.D(n_434),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3396),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3524),
.B(n_434),
.Y(n_3605)
);

HB1xp67_ASAP7_75t_L g3606 ( 
.A(n_3431),
.Y(n_3606)
);

AOI221xp5_ASAP7_75t_L g3607 ( 
.A1(n_3444),
.A2(n_3423),
.B1(n_3429),
.B2(n_3437),
.C(n_3434),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3490),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3421),
.Y(n_3609)
);

INVx2_ASAP7_75t_SL g3610 ( 
.A(n_3426),
.Y(n_3610)
);

NAND3xp33_ASAP7_75t_L g3611 ( 
.A(n_3485),
.B(n_436),
.C(n_438),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3467),
.B(n_436),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3420),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3440),
.B(n_439),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3498),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3501),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3502),
.Y(n_3617)
);

O2A1O1Ixp5_ASAP7_75t_L g3618 ( 
.A1(n_3471),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3509),
.Y(n_3619)
);

OAI211xp5_ASAP7_75t_SL g3620 ( 
.A1(n_3450),
.A2(n_445),
.B(n_443),
.C(n_444),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3401),
.B(n_443),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3460),
.B(n_444),
.Y(n_3622)
);

OAI211xp5_ASAP7_75t_L g3623 ( 
.A1(n_3451),
.A2(n_3472),
.B(n_3473),
.C(n_3463),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3510),
.Y(n_3624)
);

NAND2xp67_ASAP7_75t_SL g3625 ( 
.A(n_3589),
.B(n_3602),
.Y(n_3625)
);

NOR3x1_ASAP7_75t_L g3626 ( 
.A(n_3549),
.B(n_3405),
.C(n_3506),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_3543),
.B(n_3452),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3606),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3578),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3533),
.B(n_3537),
.Y(n_3630)
);

AOI221xp5_ASAP7_75t_L g3631 ( 
.A1(n_3536),
.A2(n_3381),
.B1(n_3449),
.B2(n_3416),
.C(n_3417),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3533),
.B(n_3391),
.Y(n_3632)
);

NAND4xp25_ASAP7_75t_L g3633 ( 
.A(n_3580),
.B(n_3493),
.C(n_3432),
.D(n_3475),
.Y(n_3633)
);

OAI21xp5_ASAP7_75t_SL g3634 ( 
.A1(n_3613),
.A2(n_3479),
.B(n_3425),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_3597),
.B(n_3476),
.Y(n_3635)
);

INVxp33_ASAP7_75t_L g3636 ( 
.A(n_3565),
.Y(n_3636)
);

NOR2xp67_ASAP7_75t_SL g3637 ( 
.A(n_3555),
.B(n_3463),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3550),
.A2(n_3400),
.B(n_3418),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3546),
.B(n_3439),
.Y(n_3639)
);

XOR2x2_ASAP7_75t_L g3640 ( 
.A(n_3553),
.B(n_3481),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3586),
.B(n_3458),
.Y(n_3641)
);

NAND3xp33_ASAP7_75t_L g3642 ( 
.A(n_3572),
.B(n_3478),
.C(n_3462),
.Y(n_3642)
);

AOI211xp5_ASAP7_75t_L g3643 ( 
.A1(n_3551),
.A2(n_3480),
.B(n_3515),
.C(n_3494),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3535),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3558),
.Y(n_3645)
);

OAI22xp5_ASAP7_75t_L g3646 ( 
.A1(n_3540),
.A2(n_3563),
.B1(n_3562),
.B2(n_3555),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3534),
.B(n_3538),
.Y(n_3647)
);

INVx1_ASAP7_75t_SL g3648 ( 
.A(n_3561),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3559),
.B(n_3477),
.Y(n_3649)
);

OAI22xp33_ASAP7_75t_L g3650 ( 
.A1(n_3544),
.A2(n_3435),
.B1(n_3441),
.B2(n_3436),
.Y(n_3650)
);

NAND4xp25_ASAP7_75t_L g3651 ( 
.A(n_3545),
.B(n_3474),
.C(n_3492),
.D(n_3482),
.Y(n_3651)
);

NOR4xp25_ASAP7_75t_SL g3652 ( 
.A(n_3552),
.B(n_3427),
.C(n_3428),
.D(n_3488),
.Y(n_3652)
);

NAND4xp75_ASAP7_75t_L g3653 ( 
.A(n_3607),
.B(n_3409),
.C(n_3447),
.D(n_3512),
.Y(n_3653)
);

AOI221x1_ASAP7_75t_L g3654 ( 
.A1(n_3560),
.A2(n_3530),
.B1(n_3528),
.B2(n_3525),
.C(n_3520),
.Y(n_3654)
);

INVxp67_ASAP7_75t_SL g3655 ( 
.A(n_3541),
.Y(n_3655)
);

OAI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3542),
.A2(n_3469),
.B1(n_3517),
.B2(n_3513),
.Y(n_3656)
);

NOR3xp33_ASAP7_75t_L g3657 ( 
.A(n_3623),
.B(n_3491),
.C(n_3456),
.Y(n_3657)
);

NOR3xp33_ASAP7_75t_L g3658 ( 
.A(n_3539),
.B(n_3496),
.C(n_3486),
.Y(n_3658)
);

NOR3xp33_ASAP7_75t_SL g3659 ( 
.A(n_3587),
.B(n_3459),
.C(n_3487),
.Y(n_3659)
);

OAI211xp5_ASAP7_75t_L g3660 ( 
.A1(n_3574),
.A2(n_3455),
.B(n_3484),
.C(n_3483),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3556),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3554),
.A2(n_3489),
.B(n_3495),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3605),
.B(n_445),
.Y(n_3663)
);

OAI21xp33_ASAP7_75t_L g3664 ( 
.A1(n_3583),
.A2(n_446),
.B(n_447),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3557),
.Y(n_3665)
);

NOR4xp25_ASAP7_75t_L g3666 ( 
.A(n_3595),
.B(n_449),
.C(n_447),
.D(n_448),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3614),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3577),
.B(n_448),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3579),
.Y(n_3669)
);

NOR2xp67_ASAP7_75t_SL g3670 ( 
.A(n_3590),
.B(n_451),
.Y(n_3670)
);

INVxp33_ASAP7_75t_L g3671 ( 
.A(n_3570),
.Y(n_3671)
);

OAI211xp5_ASAP7_75t_L g3672 ( 
.A1(n_3593),
.A2(n_451),
.B(n_453),
.C(n_454),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3592),
.B(n_453),
.Y(n_3673)
);

NAND4xp25_ASAP7_75t_L g3674 ( 
.A(n_3585),
.B(n_454),
.C(n_457),
.D(n_459),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3612),
.Y(n_3675)
);

NAND4xp25_ASAP7_75t_L g3676 ( 
.A(n_3569),
.B(n_459),
.C(n_460),
.D(n_461),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3603),
.B(n_460),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3564),
.B(n_462),
.Y(n_3678)
);

NAND3xp33_ASAP7_75t_L g3679 ( 
.A(n_3618),
.B(n_463),
.C(n_464),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_SL g3680 ( 
.A(n_3610),
.B(n_465),
.Y(n_3680)
);

NOR3xp33_ASAP7_75t_L g3681 ( 
.A(n_3622),
.B(n_465),
.C(n_467),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3566),
.Y(n_3682)
);

INVx3_ASAP7_75t_L g3683 ( 
.A(n_3609),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3575),
.B(n_468),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3666),
.B(n_3611),
.Y(n_3685)
);

NAND3x1_ASAP7_75t_L g3686 ( 
.A(n_3630),
.B(n_3584),
.C(n_3588),
.Y(n_3686)
);

INVx2_ASAP7_75t_SL g3687 ( 
.A(n_3640),
.Y(n_3687)
);

NOR5xp2_ASAP7_75t_L g3688 ( 
.A(n_3634),
.B(n_3548),
.C(n_3576),
.D(n_3604),
.E(n_3573),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3663),
.B(n_3567),
.Y(n_3689)
);

OAI211xp5_ASAP7_75t_SL g3690 ( 
.A1(n_3643),
.A2(n_3568),
.B(n_3616),
.C(n_3615),
.Y(n_3690)
);

NAND4xp25_ASAP7_75t_L g3691 ( 
.A(n_3633),
.B(n_3608),
.C(n_3619),
.D(n_3617),
.Y(n_3691)
);

HB1xp67_ASAP7_75t_L g3692 ( 
.A(n_3677),
.Y(n_3692)
);

NAND4xp25_ASAP7_75t_L g3693 ( 
.A(n_3626),
.B(n_3624),
.C(n_3594),
.D(n_3599),
.Y(n_3693)
);

NAND3xp33_ASAP7_75t_SL g3694 ( 
.A(n_3652),
.B(n_3601),
.C(n_3621),
.Y(n_3694)
);

OAI211xp5_ASAP7_75t_SL g3695 ( 
.A1(n_3631),
.A2(n_3582),
.B(n_3581),
.C(n_3571),
.Y(n_3695)
);

NAND3xp33_ASAP7_75t_L g3696 ( 
.A(n_3637),
.B(n_3591),
.C(n_3598),
.Y(n_3696)
);

INVx2_ASAP7_75t_SL g3697 ( 
.A(n_3684),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_SL g3698 ( 
.A(n_3629),
.B(n_3684),
.Y(n_3698)
);

INVx1_ASAP7_75t_SL g3699 ( 
.A(n_3632),
.Y(n_3699)
);

NOR3xp33_ASAP7_75t_L g3700 ( 
.A(n_3651),
.B(n_3596),
.C(n_3600),
.Y(n_3700)
);

OAI32xp33_ASAP7_75t_L g3701 ( 
.A1(n_3636),
.A2(n_3620),
.A3(n_3547),
.B1(n_470),
.B2(n_471),
.Y(n_3701)
);

INVxp67_ASAP7_75t_L g3702 ( 
.A(n_3627),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_3628),
.B(n_468),
.Y(n_3703)
);

NAND4xp25_ASAP7_75t_SL g3704 ( 
.A(n_3638),
.B(n_469),
.C(n_470),
.D(n_471),
.Y(n_3704)
);

NAND3xp33_ASAP7_75t_SL g3705 ( 
.A(n_3648),
.B(n_472),
.C(n_473),
.Y(n_3705)
);

NAND3xp33_ASAP7_75t_SL g3706 ( 
.A(n_3657),
.B(n_473),
.C(n_474),
.Y(n_3706)
);

OA22x2_ASAP7_75t_L g3707 ( 
.A1(n_3635),
.A2(n_3647),
.B1(n_3682),
.B2(n_3665),
.Y(n_3707)
);

NAND3xp33_ASAP7_75t_L g3708 ( 
.A(n_3681),
.B(n_474),
.C(n_476),
.Y(n_3708)
);

OA211x2_ASAP7_75t_L g3709 ( 
.A1(n_3664),
.A2(n_477),
.B(n_479),
.C(n_480),
.Y(n_3709)
);

OAI221xp5_ASAP7_75t_L g3710 ( 
.A1(n_3639),
.A2(n_3683),
.B1(n_3659),
.B2(n_3644),
.C(n_3679),
.Y(n_3710)
);

AOI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3680),
.A2(n_479),
.B(n_481),
.Y(n_3711)
);

NOR5xp2_ASAP7_75t_L g3712 ( 
.A(n_3642),
.B(n_482),
.C(n_484),
.D(n_485),
.E(n_486),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_SL g3713 ( 
.A(n_3683),
.B(n_482),
.Y(n_3713)
);

NAND3xp33_ASAP7_75t_L g3714 ( 
.A(n_3670),
.B(n_484),
.C(n_485),
.Y(n_3714)
);

NOR2x1_ASAP7_75t_L g3715 ( 
.A(n_3646),
.B(n_486),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3668),
.A2(n_3678),
.B(n_3676),
.Y(n_3716)
);

AOI221x1_ASAP7_75t_L g3717 ( 
.A1(n_3669),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.C(n_490),
.Y(n_3717)
);

AOI22x1_ASAP7_75t_L g3718 ( 
.A1(n_3662),
.A2(n_487),
.B1(n_489),
.B2(n_490),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3671),
.B(n_492),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3667),
.B(n_492),
.Y(n_3720)
);

NAND3xp33_ASAP7_75t_L g3721 ( 
.A(n_3700),
.B(n_3654),
.C(n_3649),
.Y(n_3721)
);

A2O1A1Ixp33_ASAP7_75t_L g3722 ( 
.A1(n_3687),
.A2(n_3673),
.B(n_3655),
.C(n_3645),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3699),
.A2(n_3653),
.B1(n_3641),
.B2(n_3675),
.Y(n_3723)
);

AOI31xp33_ASAP7_75t_L g3724 ( 
.A1(n_3698),
.A2(n_3661),
.A3(n_3660),
.B(n_3650),
.Y(n_3724)
);

AND2x4_ASAP7_75t_L g3725 ( 
.A(n_3697),
.B(n_3658),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3719),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3707),
.B(n_3672),
.Y(n_3727)
);

AOI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3694),
.A2(n_3656),
.B1(n_3674),
.B2(n_3625),
.Y(n_3728)
);

INVxp67_ASAP7_75t_L g3729 ( 
.A(n_3715),
.Y(n_3729)
);

NAND4xp25_ASAP7_75t_SL g3730 ( 
.A(n_3710),
.B(n_493),
.C(n_494),
.D(n_495),
.Y(n_3730)
);

XNOR2xp5_ASAP7_75t_L g3731 ( 
.A(n_3686),
.B(n_3709),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3692),
.A2(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_3732)
);

OAI21xp33_ASAP7_75t_SL g3733 ( 
.A1(n_3691),
.A2(n_496),
.B(n_497),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3689),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3718),
.Y(n_3735)
);

A2O1A1Ixp33_ASAP7_75t_L g3736 ( 
.A1(n_3696),
.A2(n_497),
.B(n_498),
.C(n_499),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_3685),
.Y(n_3737)
);

OAI21xp33_ASAP7_75t_L g3738 ( 
.A1(n_3690),
.A2(n_500),
.B(n_501),
.Y(n_3738)
);

NOR2x1_ASAP7_75t_L g3739 ( 
.A(n_3703),
.B(n_501),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_3737),
.B(n_3701),
.Y(n_3740)
);

NOR3xp33_ASAP7_75t_L g3741 ( 
.A(n_3721),
.B(n_3702),
.C(n_3695),
.Y(n_3741)
);

AOI21xp33_ASAP7_75t_SL g3742 ( 
.A1(n_3724),
.A2(n_3713),
.B(n_3714),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3727),
.Y(n_3743)
);

CKINVDCx20_ASAP7_75t_R g3744 ( 
.A(n_3726),
.Y(n_3744)
);

NOR3xp33_ASAP7_75t_L g3745 ( 
.A(n_3723),
.B(n_3720),
.C(n_3693),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3725),
.Y(n_3746)
);

NAND3xp33_ASAP7_75t_SL g3747 ( 
.A(n_3728),
.B(n_3688),
.C(n_3712),
.Y(n_3747)
);

NOR2x1_ASAP7_75t_L g3748 ( 
.A(n_3730),
.B(n_3704),
.Y(n_3748)
);

NOR2x1_ASAP7_75t_L g3749 ( 
.A(n_3734),
.B(n_3706),
.Y(n_3749)
);

NOR2x1_ASAP7_75t_L g3750 ( 
.A(n_3735),
.B(n_3705),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3731),
.B(n_3717),
.Y(n_3751)
);

NAND4xp75_ASAP7_75t_L g3752 ( 
.A(n_3739),
.B(n_3716),
.C(n_3711),
.D(n_3708),
.Y(n_3752)
);

NOR3xp33_ASAP7_75t_L g3753 ( 
.A(n_3746),
.B(n_3722),
.C(n_3725),
.Y(n_3753)
);

NAND3xp33_ASAP7_75t_L g3754 ( 
.A(n_3741),
.B(n_3745),
.C(n_3740),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3750),
.B(n_3729),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3748),
.B(n_3738),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3744),
.A2(n_3733),
.B1(n_3732),
.B2(n_3736),
.Y(n_3757)
);

NAND2x1p5_ASAP7_75t_L g3758 ( 
.A(n_3749),
.B(n_502),
.Y(n_3758)
);

NAND3xp33_ASAP7_75t_L g3759 ( 
.A(n_3742),
.B(n_502),
.C(n_503),
.Y(n_3759)
);

AOI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3751),
.A2(n_504),
.B1(n_506),
.B2(n_507),
.Y(n_3760)
);

AOI21xp33_ASAP7_75t_SL g3761 ( 
.A1(n_3743),
.A2(n_506),
.B(n_508),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3752),
.B(n_508),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3758),
.B(n_3747),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3755),
.Y(n_3764)
);

INVxp67_ASAP7_75t_SL g3765 ( 
.A(n_3753),
.Y(n_3765)
);

INVxp33_ASAP7_75t_L g3766 ( 
.A(n_3762),
.Y(n_3766)
);

NOR2x1_ASAP7_75t_L g3767 ( 
.A(n_3754),
.B(n_509),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3765),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3763),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3764),
.A2(n_3756),
.B1(n_3757),
.B2(n_3759),
.Y(n_3770)
);

NAND3xp33_ASAP7_75t_L g3771 ( 
.A(n_3767),
.B(n_3761),
.C(n_3760),
.Y(n_3771)
);

AOI21xp33_ASAP7_75t_L g3772 ( 
.A1(n_3768),
.A2(n_3766),
.B(n_510),
.Y(n_3772)
);

OAI211xp5_ASAP7_75t_SL g3773 ( 
.A1(n_3772),
.A2(n_3770),
.B(n_3769),
.C(n_3771),
.Y(n_3773)
);

AOI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3773),
.A2(n_511),
.B(n_512),
.Y(n_3774)
);

O2A1O1Ixp33_ASAP7_75t_L g3775 ( 
.A1(n_3774),
.A2(n_512),
.B(n_514),
.C(n_515),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3775),
.Y(n_3776)
);

OAI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3776),
.A2(n_514),
.B(n_515),
.Y(n_3777)
);

AOI222xp33_ASAP7_75t_SL g3778 ( 
.A1(n_3777),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.C1(n_519),
.C2(n_521),
.Y(n_3778)
);

HB1xp67_ASAP7_75t_L g3779 ( 
.A(n_3778),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3778),
.Y(n_3780)
);

AOI21xp33_ASAP7_75t_SL g3781 ( 
.A1(n_3780),
.A2(n_519),
.B(n_521),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3781),
.A2(n_3779),
.B(n_523),
.Y(n_3782)
);

AOI211xp5_ASAP7_75t_L g3783 ( 
.A1(n_3782),
.A2(n_523),
.B(n_524),
.C(n_525),
.Y(n_3783)
);


endmodule