module fake_jpeg_19647_n_344 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_43),
.B1(n_48),
.B2(n_45),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_62),
.B1(n_25),
.B2(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_19),
.B1(n_15),
.B2(n_22),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_99),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_35),
.B1(n_36),
.B2(n_22),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_48),
.B1(n_41),
.B2(n_22),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_81),
.B1(n_84),
.B2(n_88),
.Y(n_107)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_35),
.B1(n_15),
.B2(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_93),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_49),
.B1(n_15),
.B2(n_35),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_16),
.B1(n_24),
.B2(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_91),
.B1(n_97),
.B2(n_100),
.Y(n_108)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_86),
.Y(n_134)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_36),
.B1(n_41),
.B2(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_26),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_28),
.B1(n_29),
.B2(n_26),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_26),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_25),
.B1(n_47),
.B2(n_44),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_47),
.B1(n_46),
.B2(n_44),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_23),
.B(n_26),
.C(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_123)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_23),
.B1(n_18),
.B2(n_30),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_95),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_77),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_111),
.B(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_133),
.B1(n_136),
.B2(n_107),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_23),
.B1(n_32),
.B2(n_18),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_101),
.B1(n_93),
.B2(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_34),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_SL g135 ( 
.A(n_78),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_135),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_71),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_157),
.C(n_128),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_117),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_147),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_102),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_87),
.B1(n_79),
.B2(n_70),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_152),
.B(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_66),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_100),
.B1(n_110),
.B2(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_158),
.B1(n_133),
.B2(n_125),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_67),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_120),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_161),
.B1(n_125),
.B2(n_137),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_106),
.B(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_108),
.A2(n_98),
.B1(n_75),
.B2(n_65),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_98),
.B1(n_89),
.B2(n_2),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_73),
.A3(n_69),
.B1(n_18),
.B2(n_74),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_164),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_104),
.B(n_74),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_142),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_118),
.B(n_111),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_179),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_171),
.B1(n_189),
.B2(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_125),
.B1(n_132),
.B2(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_181),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_178),
.B1(n_184),
.B2(n_194),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_125),
.B1(n_130),
.B2(n_121),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_131),
.B(n_121),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_112),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_130),
.B1(n_117),
.B2(n_128),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_192),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_124),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_134),
.B1(n_116),
.B2(n_124),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_141),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_23),
.B(n_104),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_1),
.B(n_3),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_116),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_34),
.B(n_33),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_152),
.B(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_116),
.B1(n_34),
.B2(n_33),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_33),
.B1(n_30),
.B2(n_2),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_152),
.B1(n_143),
.B2(n_2),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_198),
.A2(n_215),
.B1(n_222),
.B2(n_184),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_209),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_147),
.B(n_162),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_203),
.B(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_225),
.B1(n_176),
.B2(n_182),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_219),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_157),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_143),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_0),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_0),
.C(n_1),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_166),
.C(n_172),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_168),
.B(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_169),
.B1(n_188),
.B2(n_189),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_4),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_4),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_227),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_188),
.B1(n_193),
.B2(n_165),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_239),
.C(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_245),
.C(n_252),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_168),
.C(n_173),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_251),
.Y(n_274)
);

XNOR2x2_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_173),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_166),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_194),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_198),
.B1(n_210),
.B2(n_223),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_257),
.A2(n_270),
.B1(n_273),
.B2(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_263),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_201),
.CI(n_197),
.CON(n_263),
.SN(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_272),
.Y(n_281)
);

BUFx12f_ASAP7_75t_SL g269 ( 
.A(n_238),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_269),
.A2(n_271),
.B(n_203),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_197),
.B1(n_199),
.B2(n_215),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_219),
.B(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_216),
.B1(n_243),
.B2(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_252),
.C(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_283),
.C(n_279),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_280),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_230),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_225),
.B1(n_228),
.B2(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_240),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_237),
.B(n_242),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_289),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_292),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_229),
.B1(n_211),
.B2(n_244),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_239),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_280),
.C(n_288),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_293),
.B(n_294),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_228),
.C(n_263),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_275),
.A2(n_208),
.B1(n_257),
.B2(n_270),
.Y(n_295)
);

AOI22x1_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_176),
.B1(n_211),
.B2(n_207),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_234),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_277),
.B1(n_291),
.B2(n_172),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_263),
.C(n_254),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_214),
.C(n_200),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_273),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_262),
.C(n_261),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_5),
.C(n_6),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_285),
.B1(n_262),
.B2(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_310),
.A2(n_313),
.B1(n_315),
.B2(n_304),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_318),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_276),
.B1(n_220),
.B2(n_200),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_295),
.B1(n_307),
.B2(n_301),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_220),
.B1(n_226),
.B2(n_195),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_182),
.C(n_6),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_6),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_298),
.B(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_316),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_302),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_314),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_304),
.B(n_8),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_318),
.C(n_312),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_7),
.B(n_8),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_334),
.B(n_330),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_331),
.Y(n_339)
);

NOR4xp25_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_333),
.C(n_336),
.D(n_10),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_8),
.B(n_9),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_344)
);


endmodule