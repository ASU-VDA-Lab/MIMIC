module fake_ariane_2752_n_1863 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1863);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1863;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_91),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_24),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_47),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_24),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_116),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_67),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_29),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_115),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

BUFx8_ASAP7_75t_SL g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_124),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_137),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_117),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_145),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_94),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_164),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_102),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_0),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_1),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_59),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_150),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_40),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_136),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_146),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_144),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_33),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_40),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_60),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_87),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_37),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_73),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_109),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_68),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_22),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_75),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_43),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_76),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_33),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

BUFx2_ASAP7_75t_SL g269 ( 
.A(n_147),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_127),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_39),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_99),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_169),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_82),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_112),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_178),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_89),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_28),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_77),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_32),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_172),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_132),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_27),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_41),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_36),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_59),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_64),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_103),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_41),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_83),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_182),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_52),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_93),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_170),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_119),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_151),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_110),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_86),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_174),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_179),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_56),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_166),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_29),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_0),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_98),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_111),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_18),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_2),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_27),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_50),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_22),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_80),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_70),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_168),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_74),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_23),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_54),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_26),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_92),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_152),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_45),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_44),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_107),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_32),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_9),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_159),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_19),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_26),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_58),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_13),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_8),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_21),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_3),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_13),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_18),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_30),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_165),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_43),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_35),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_154),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_58),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_21),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_148),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_121),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_175),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_139),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_23),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_17),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_173),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_31),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_31),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_11),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_50),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_214),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_212),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_286),
.B(n_2),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_221),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_240),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_277),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_277),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_264),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_277),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_267),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_314),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_206),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_247),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_206),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_353),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_228),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_231),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_206),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_192),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_232),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_206),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_3),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_220),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_199),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_241),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_206),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_4),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_236),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_282),
.B(n_7),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_297),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_185),
.B(n_9),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_237),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_312),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_340),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_192),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_194),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_244),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_249),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_239),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_254),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_239),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_339),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_251),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_258),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_266),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_268),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_315),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_259),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_259),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_351),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_270),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_340),
.B(n_10),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_348),
.B(n_12),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_348),
.B(n_12),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_227),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_326),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_227),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_326),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_227),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_329),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_313),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_329),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_313),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_313),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_357),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_224),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_272),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_273),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_285),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_224),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_291),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_307),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_295),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_305),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_307),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_188),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_317),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_357),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_357),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_191),
.B(n_20),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_318),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_211),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_213),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_385),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_196),
.B(n_193),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_389),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_376),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_379),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_399),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_400),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_382),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_384),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_413),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_422),
.B(n_431),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_210),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_436),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_368),
.Y(n_496)
);

NAND2x1_ASAP7_75t_L g497 ( 
.A(n_377),
.B(n_210),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_420),
.B(n_186),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_436),
.B(n_198),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_372),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_375),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_392),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_R g507 ( 
.A(n_409),
.B(n_197),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_417),
.B(n_262),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_420),
.B(n_186),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_377),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_262),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_R g513 ( 
.A(n_373),
.B(n_418),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_378),
.B(n_234),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_388),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_454),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_383),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_378),
.B(n_235),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_381),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_381),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_462),
.A2(n_278),
.B(n_255),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_425),
.B(n_226),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_428),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_371),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_426),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_419),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_427),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_432),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_414),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_471),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_493),
.B(n_508),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_428),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_511),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_536),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_507),
.A2(n_374),
.B1(n_443),
.B2(n_439),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_449),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_525),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_533),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_496),
.B(n_450),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_535),
.B(n_539),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_453),
.C(n_451),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_498),
.B(n_455),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_484),
.B(n_443),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_496),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_516),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_516),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_509),
.B(n_456),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_544),
.B(n_518),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_518),
.B(n_459),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_532),
.B(n_220),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_532),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_513),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_532),
.B(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_525),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_484),
.B(n_386),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_523),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_516),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_510),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_524),
.B(n_445),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_526),
.B(n_446),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_505),
.B(n_386),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_482),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_472),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_527),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_499),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_512),
.B(n_465),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_470),
.B(n_394),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_505),
.B(n_390),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_469),
.B(n_433),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_473),
.A2(n_397),
.B1(n_341),
.B2(n_369),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_525),
.B(n_280),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_501),
.B(n_415),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_434),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_478),
.B(n_380),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_469),
.A2(n_403),
.B1(n_435),
.B2(n_342),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_528),
.B(n_458),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_515),
.B(n_281),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_528),
.B(n_220),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_541),
.B(n_458),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_515),
.B(n_284),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_530),
.B(n_287),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_528),
.B(n_220),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_497),
.B(n_464),
.Y(n_623)
);

INVx4_ASAP7_75t_SL g624 ( 
.A(n_500),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_530),
.B(n_293),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_469),
.A2(n_534),
.B1(n_542),
.B2(n_499),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_542),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_467),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_497),
.B(n_464),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

INVx4_ASAP7_75t_SL g631 ( 
.A(n_500),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_469),
.A2(n_261),
.B1(n_265),
.B2(n_257),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_488),
.B(n_197),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_534),
.A2(n_248),
.B1(n_325),
.B2(n_310),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_534),
.Y(n_635)
);

INVx4_ASAP7_75t_SL g636 ( 
.A(n_500),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_474),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_534),
.B(n_195),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_542),
.B(n_301),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_542),
.B(n_304),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_542),
.B(n_276),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_537),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_421),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_542),
.B(n_323),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_476),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_540),
.A2(n_253),
.B1(n_319),
.B2(n_330),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_500),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_540),
.B(n_421),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_479),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_479),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_486),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_486),
.B(n_306),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_468),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_481),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_481),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_485),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_485),
.B(n_429),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_500),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_480),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_500),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_489),
.B(n_187),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_489),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_492),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_429),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_468),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_504),
.A2(n_334),
.B1(n_208),
.B2(n_203),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_468),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_506),
.B(n_187),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_468),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_506),
.B(n_514),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_514),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_517),
.B(n_437),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_468),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_520),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_520),
.B(n_189),
.Y(n_680)
);

INVx4_ASAP7_75t_SL g681 ( 
.A(n_521),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_521),
.B(n_441),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_522),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_529),
.B(n_405),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_522),
.B(n_447),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_480),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_480),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_483),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_480),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_475),
.A2(n_346),
.B1(n_300),
.B2(n_361),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_490),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_475),
.B(n_460),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_475),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_477),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_477),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_604),
.B(n_189),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_575),
.B(n_502),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_679),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_566),
.A2(n_201),
.B1(n_223),
.B2(n_222),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_549),
.A2(n_208),
.B(n_203),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_559),
.B(n_320),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_566),
.A2(n_200),
.B1(n_223),
.B2(n_222),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_597),
.B(n_548),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_551),
.B(n_190),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_574),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_604),
.B(n_679),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_545),
.B(n_629),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_545),
.B(n_619),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_550),
.B(n_321),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_591),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_576),
.B(n_328),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_679),
.B(n_190),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_619),
.B(n_200),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_679),
.B(n_201),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_556),
.B(n_202),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_547),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_562),
.A2(n_570),
.B1(n_589),
.B2(n_586),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_202),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_555),
.A2(n_332),
.B1(n_218),
.B2(n_216),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_600),
.A2(n_332),
.B1(n_218),
.B2(n_216),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_565),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_547),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_503),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_563),
.A2(n_289),
.B(n_296),
.C(n_229),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_578),
.B(n_204),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_581),
.B(n_204),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_611),
.B(n_217),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_630),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_584),
.B(n_205),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_557),
.B(n_205),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_632),
.A2(n_405),
.B1(n_292),
.B2(n_246),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_557),
.B(n_207),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_646),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_575),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_583),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_588),
.B(n_207),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_634),
.A2(n_290),
.B1(n_368),
.B2(n_444),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_592),
.B(n_215),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_595),
.A2(n_598),
.B1(n_602),
.B2(n_596),
.Y(n_742)
);

AND2x6_ASAP7_75t_SL g743 ( 
.A(n_645),
.B(n_593),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_646),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_593),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_217),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_660),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_633),
.A2(n_225),
.B1(n_334),
.B2(n_336),
.C(n_343),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_603),
.B(n_215),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_583),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_557),
.B(n_279),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_565),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_279),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_617),
.B(n_335),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_630),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_637),
.B(n_461),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_617),
.B(n_335),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_688),
.B(n_430),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_623),
.A2(n_358),
.B1(n_360),
.B2(n_362),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_553),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_620),
.B(n_358),
.Y(n_762)
);

AND3x1_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_440),
.C(n_430),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_557),
.B(n_360),
.Y(n_764)
);

INVxp33_ASAP7_75t_L g765 ( 
.A(n_613),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_620),
.B(n_362),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_585),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_684),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_645),
.B(n_561),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_691),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_585),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_590),
.B(n_491),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_668),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_668),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_621),
.B(n_219),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_554),
.B(n_219),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_621),
.B(n_225),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_661),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_564),
.B(n_338),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_SL g783 ( 
.A(n_682),
.B(n_685),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_587),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_625),
.B(n_283),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_628),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_599),
.B(n_612),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_587),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_594),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_625),
.B(n_283),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_571),
.B(n_336),
.C(n_344),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_590),
.B(n_491),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_690),
.A2(n_365),
.B1(n_343),
.B2(n_349),
.C(n_352),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_560),
.B(n_440),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_614),
.A2(n_352),
.B1(n_344),
.B2(n_347),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_594),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_564),
.B(n_350),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_601),
.B(n_347),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_684),
.Y(n_799)
);

OAI221xp5_ASAP7_75t_L g800 ( 
.A1(n_649),
.A2(n_355),
.B1(n_349),
.B2(n_365),
.C(n_367),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_651),
.B(n_355),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_651),
.A2(n_368),
.B1(n_444),
.B2(n_442),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_648),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_692),
.B(n_364),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_651),
.B(n_364),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_686),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_653),
.B(n_367),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_370),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_670),
.B(n_370),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_658),
.B(n_230),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_623),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_659),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_686),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_675),
.B(n_233),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_672),
.B(n_356),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_571),
.B(n_442),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_623),
.A2(n_269),
.B1(n_359),
.B2(n_242),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_238),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_680),
.B(n_567),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_623),
.A2(n_294),
.B1(n_243),
.B2(n_245),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_689),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_689),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_560),
.B(n_250),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_609),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_609),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_643),
.B(n_25),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_633),
.A2(n_302),
.B1(n_252),
.B2(n_256),
.C(n_327),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_643),
.B(n_654),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_567),
.B(n_260),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_643),
.B(n_30),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_568),
.B(n_288),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_568),
.B(n_288),
.Y(n_832)
);

NOR3x1_ASAP7_75t_L g833 ( 
.A(n_572),
.B(n_34),
.C(n_36),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_572),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_635),
.A2(n_220),
.B1(n_366),
.B2(n_288),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_610),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_582),
.B(n_674),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_582),
.B(n_288),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_654),
.B(n_288),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_635),
.B(n_303),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_569),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_610),
.B(n_38),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_654),
.B(n_299),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_639),
.B(n_38),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_569),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_662),
.B(n_308),
.Y(n_846)
);

BUFx5_ASAP7_75t_L g847 ( 
.A(n_573),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_662),
.B(n_42),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_638),
.B(n_298),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_642),
.A2(n_366),
.B1(n_288),
.B2(n_495),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_642),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_652),
.B(n_309),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_652),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_657),
.B(n_263),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_665),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_665),
.B(n_288),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_666),
.B(n_311),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_644),
.B(n_42),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_666),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_667),
.B(n_288),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_667),
.B(n_324),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_683),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_683),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_647),
.B(n_687),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_783),
.A2(n_655),
.B1(n_569),
.B2(n_579),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_745),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_730),
.A2(n_655),
.B(n_640),
.C(n_641),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_704),
.A2(n_607),
.B(n_669),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_738),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_839),
.A2(n_607),
.B(n_669),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_839),
.A2(n_669),
.B(n_671),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_837),
.A2(n_819),
.B(n_828),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_787),
.B(n_626),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_787),
.B(n_627),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_730),
.A2(n_608),
.B(n_640),
.C(n_641),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_726),
.B(n_693),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_786),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_771),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_707),
.A2(n_694),
.B(n_477),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_779),
.B(n_579),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_864),
.B(n_832),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_765),
.B(n_579),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_719),
.A2(n_742),
.B1(n_709),
.B2(n_804),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_742),
.A2(n_656),
.B1(n_671),
.B2(n_650),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_708),
.B(n_693),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_811),
.B(n_650),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_696),
.A2(n_656),
.B(n_693),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_804),
.B(n_663),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_747),
.A2(n_656),
.B1(n_663),
.B2(n_661),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_815),
.A2(n_661),
.B(n_695),
.C(n_678),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_759),
.A2(n_661),
.B1(n_678),
.B2(n_673),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_803),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_701),
.A2(n_681),
.B1(n_573),
.B2(n_274),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_812),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_723),
.B(n_678),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_824),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_774),
.A2(n_678),
.B1(n_673),
.B2(n_546),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_697),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_831),
.A2(n_673),
.B(n_546),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_843),
.A2(n_702),
.B(n_731),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_711),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_712),
.B(n_681),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_775),
.A2(n_673),
.B1(n_546),
.B2(n_695),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_752),
.B(n_695),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_809),
.B(n_722),
.C(n_748),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_825),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_777),
.B(n_681),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_755),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_701),
.A2(n_695),
.B1(n_316),
.B2(n_275),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_808),
.A2(n_271),
.B(n_495),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_712),
.B(n_636),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_773),
.B(n_573),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_767),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_838),
.A2(n_495),
.B(n_366),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_834),
.B(n_45),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_761),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_697),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_838),
.A2(n_366),
.B(n_631),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_707),
.A2(n_717),
.B(n_856),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_799),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_710),
.B(n_636),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_856),
.A2(n_366),
.B(n_631),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_756),
.B(n_710),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_800),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_755),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_860),
.A2(n_636),
.B(n_631),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_860),
.A2(n_624),
.B(n_573),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_817),
.B(n_624),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_792),
.B(n_51),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_781),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_760),
.B(n_624),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_808),
.B(n_736),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_836),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_725),
.B(n_798),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_744),
.B(n_573),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_781),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_705),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_829),
.A2(n_622),
.B(n_618),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_R g939 ( 
.A(n_761),
.B(n_622),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_715),
.B(n_53),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_816),
.B(n_55),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_815),
.B(n_57),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_802),
.B(n_57),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_802),
.B(n_740),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_758),
.B(n_62),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_700),
.B(n_63),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_758),
.B(n_65),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_770),
.A2(n_622),
.B1(n_618),
.B2(n_71),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_758),
.B(n_622),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_740),
.B(n_734),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_734),
.B(n_618),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_794),
.B(n_725),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_791),
.B(n_622),
.C(n_618),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_746),
.B(n_618),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_699),
.B(n_66),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_770),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_789),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_789),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_750),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_713),
.A2(n_69),
.B(n_72),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_796),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_851),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_746),
.B(n_778),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_725),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_768),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_743),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_713),
.A2(n_79),
.B(n_84),
.Y(n_967)
);

OAI21xp33_ASAP7_75t_L g968 ( 
.A1(n_703),
.A2(n_88),
.B(n_97),
.Y(n_968)
);

OR2x2_ASAP7_75t_SL g969 ( 
.A(n_768),
.B(n_100),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_820),
.B(n_101),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_858),
.A2(n_104),
.B(n_108),
.C(n_113),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_795),
.A2(n_114),
.B(n_120),
.C(n_122),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_SL g973 ( 
.A1(n_826),
.A2(n_129),
.B(n_130),
.C(n_133),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_855),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_716),
.A2(n_134),
.B(n_141),
.Y(n_975)
);

OAI321xp33_ASAP7_75t_L g976 ( 
.A1(n_721),
.A2(n_142),
.A3(n_158),
.B1(n_161),
.B2(n_163),
.C(n_167),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_793),
.A2(n_171),
.B(n_183),
.C(n_807),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_718),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_716),
.A2(n_764),
.B(n_751),
.C(n_733),
.Y(n_979)
);

AOI33xp33_ASAP7_75t_L g980 ( 
.A1(n_727),
.A2(n_706),
.A3(n_714),
.B1(n_842),
.B2(n_859),
.B3(n_827),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_794),
.B(n_776),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_796),
.B(n_718),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_778),
.B(n_826),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_733),
.A2(n_764),
.B(n_751),
.C(n_735),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_861),
.B(n_857),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_731),
.A2(n_830),
.B1(n_835),
.B2(n_848),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_794),
.B(n_801),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_805),
.B(n_763),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_830),
.A2(n_735),
.B(n_814),
.C(n_818),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_769),
.B(n_823),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_781),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_844),
.A2(n_858),
.B(n_840),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_781),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_780),
.B(n_790),
.C(n_785),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_835),
.A2(n_848),
.B1(n_720),
.B2(n_739),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_SL g996 ( 
.A(n_844),
.B(n_724),
.Y(n_996)
);

AND2x4_ASAP7_75t_SL g997 ( 
.A(n_698),
.B(n_862),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_833),
.B(n_766),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_754),
.B(n_757),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_852),
.A2(n_854),
.B(n_863),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_853),
.A2(n_806),
.B(n_813),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_762),
.B(n_728),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_729),
.B(n_732),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_821),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_SL g1005 ( 
.A(n_847),
.B(n_741),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_841),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_822),
.A2(n_810),
.B(n_846),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_772),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_749),
.A2(n_753),
.B(n_788),
.C(n_784),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_845),
.B(n_782),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_797),
.B(n_850),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_847),
.B(n_549),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_847),
.A2(n_734),
.B1(n_740),
.B2(n_604),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_847),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_847),
.A2(n_783),
.B1(n_804),
.B2(n_730),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_847),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_787),
.B(n_549),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_783),
.B(n_719),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_737),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_787),
.B(n_549),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_704),
.A2(n_839),
.B(n_837),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_783),
.B(n_719),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_828),
.A2(n_704),
.B(n_839),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_704),
.A2(n_549),
.B1(n_779),
.B2(n_719),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_787),
.B(n_549),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_726),
.B(n_777),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_783),
.B(n_719),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_786),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_726),
.B(n_777),
.Y(n_1029)
);

O2A1O1Ixp5_ASAP7_75t_L g1030 ( 
.A1(n_719),
.A2(n_549),
.B(n_716),
.C(n_713),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_779),
.B(n_783),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_704),
.A2(n_549),
.B1(n_779),
.B2(n_719),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_786),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_787),
.B(n_549),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_811),
.B(n_737),
.Y(n_1035)
);

AOI22x1_ASAP7_75t_L g1036 ( 
.A1(n_731),
.A2(n_706),
.B1(n_714),
.B2(n_702),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_787),
.B(n_549),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_704),
.A2(n_839),
.B(n_837),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_704),
.A2(n_549),
.B1(n_779),
.B2(n_719),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_783),
.B(n_719),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_726),
.B(n_777),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_730),
.A2(n_549),
.B(n_779),
.C(n_719),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_704),
.A2(n_839),
.B(n_837),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_704),
.A2(n_839),
.B(n_837),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_787),
.B(n_549),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_SL g1046 ( 
.A(n_725),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_964),
.B(n_878),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_901),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1035),
.B(n_1019),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_919),
.A2(n_887),
.B(n_870),
.Y(n_1052)
);

AOI221xp5_ASAP7_75t_L g1053 ( 
.A1(n_929),
.A2(n_883),
.B1(n_905),
.B2(n_1025),
.C(n_1034),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_SL g1054 ( 
.A1(n_1031),
.A2(n_1042),
.B(n_1037),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_877),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_L g1056 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_1027),
.C(n_1040),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1045),
.A2(n_872),
.B(n_986),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_963),
.B(n_1024),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_992),
.A2(n_881),
.B(n_872),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1035),
.B(n_1019),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1030),
.A2(n_983),
.B(n_995),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1032),
.B(n_1039),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_881),
.A2(n_1007),
.B(n_1000),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_866),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1015),
.A2(n_946),
.B(n_942),
.C(n_924),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_993),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1012),
.A2(n_874),
.B(n_1023),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_SL g1068 ( 
.A(n_916),
.B(n_917),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_SL g1069 ( 
.A1(n_1007),
.A2(n_972),
.B(n_985),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_950),
.A2(n_944),
.B(n_1013),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_868),
.A2(n_1001),
.B(n_871),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1026),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_920),
.A2(n_923),
.B1(n_1041),
.B2(n_1029),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_873),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_898),
.Y(n_1075)
);

INVx5_ASAP7_75t_L g1076 ( 
.A(n_1014),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1001),
.A2(n_871),
.B(n_922),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_934),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_876),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_888),
.A2(n_900),
.B(n_1043),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_902),
.B(n_911),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_922),
.A2(n_918),
.B(n_914),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_908),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_932),
.B(n_1003),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_SL g1085 ( 
.A1(n_985),
.A2(n_960),
.B(n_975),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1021),
.A2(n_1043),
.B(n_1038),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_945),
.B(n_988),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_987),
.B(n_907),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_965),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1044),
.A2(n_989),
.B(n_921),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_938),
.A2(n_954),
.B(n_889),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1002),
.A2(n_979),
.B(n_1009),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_867),
.A2(n_875),
.B(n_981),
.C(n_968),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_926),
.A2(n_927),
.B(n_899),
.Y(n_1094)
);

BUFx5_ASAP7_75t_L g1095 ( 
.A(n_1008),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_966),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_984),
.A2(n_885),
.B(n_884),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1005),
.A2(n_890),
.B(n_891),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_938),
.A2(n_1011),
.A3(n_975),
.B(n_967),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_952),
.A2(n_947),
.B1(n_915),
.B2(n_990),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_994),
.A2(n_940),
.B(n_935),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_980),
.A2(n_943),
.B(n_937),
.C(n_977),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_913),
.Y(n_1103)
);

OAI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_951),
.A2(n_941),
.B1(n_925),
.B2(n_999),
.C1(n_896),
.C2(n_933),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_930),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_892),
.B(n_894),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_955),
.A2(n_976),
.B(n_970),
.C(n_967),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_912),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_880),
.A2(n_897),
.B(n_903),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_957),
.B(n_961),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_906),
.A2(n_962),
.B(n_974),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_928),
.A2(n_931),
.B(n_960),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1028),
.B(n_1033),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_959),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_998),
.B(n_895),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_971),
.A2(n_1004),
.A3(n_1010),
.B(n_948),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_865),
.A2(n_910),
.B(n_893),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_882),
.B(n_1006),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_949),
.B(n_958),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_886),
.A2(n_991),
.B(n_982),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_957),
.B(n_958),
.Y(n_1121)
);

AO32x2_ASAP7_75t_L g1122 ( 
.A1(n_978),
.A2(n_909),
.A3(n_1016),
.B1(n_956),
.B2(n_908),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_996),
.A2(n_978),
.B(n_973),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_904),
.B(n_1006),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_930),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_939),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1046),
.A2(n_997),
.B1(n_953),
.B2(n_886),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1014),
.A2(n_936),
.A3(n_969),
.B(n_1046),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_936),
.B(n_1015),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1017),
.A2(n_1020),
.B1(n_1034),
.B2(n_1025),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1035),
.B(n_811),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_878),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1035),
.B(n_811),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_877),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_883),
.A2(n_919),
.B(n_1015),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_877),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1035),
.B(n_811),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_878),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_869),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_1018),
.A2(n_1027),
.B(n_1040),
.C(n_1022),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1026),
.B(n_726),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_993),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1017),
.A2(n_1020),
.B1(n_1034),
.B2(n_1025),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_993),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_SL g1153 ( 
.A1(n_883),
.A2(n_919),
.B(n_1015),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1017),
.A2(n_1020),
.B1(n_1034),
.B2(n_1025),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1035),
.B(n_811),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1035),
.B(n_811),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_SL g1159 ( 
.A1(n_883),
.A2(n_919),
.B(n_1015),
.Y(n_1159)
);

AOI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_983),
.A2(n_783),
.B(n_484),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1034),
.C(n_1020),
.Y(n_1161)
);

AND3x4_ASAP7_75t_L g1162 ( 
.A(n_866),
.B(n_923),
.C(n_791),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_905),
.A2(n_783),
.B1(n_779),
.B2(n_593),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_877),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_916),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1034),
.C(n_1020),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_983),
.A2(n_783),
.B(n_484),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_869),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1026),
.B(n_726),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1042),
.B(n_783),
.C(n_779),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_993),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_869),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1035),
.B(n_811),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_869),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_901),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_869),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1017),
.B(n_1020),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1026),
.B(n_726),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_877),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_879),
.A2(n_1036),
.B(n_919),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1020),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1058),
.B(n_1062),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1105),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1058),
.A2(n_1057),
.B(n_1061),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1147),
.A2(n_1170),
.B(n_1165),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1055),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1049),
.B(n_1126),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1114),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1198)
);

OR2x2_ASAP7_75t_SL g1199 ( 
.A(n_1047),
.B(n_1142),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1053),
.A2(n_1130),
.B1(n_1155),
.B2(n_1150),
.Y(n_1200)
);

AOI21xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1163),
.A2(n_1162),
.B(n_1149),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1146),
.B(n_1154),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1066),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1056),
.A2(n_1144),
.B(n_1161),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1161),
.A2(n_1167),
.B1(n_1177),
.B2(n_1183),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1064),
.Y(n_1207)
);

INVx6_ASAP7_75t_SL g1208 ( 
.A(n_1049),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1160),
.A2(n_1168),
.B1(n_1070),
.B2(n_1084),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1091),
.A2(n_1081),
.B(n_1059),
.Y(n_1210)
);

AOI222xp33_ASAP7_75t_L g1211 ( 
.A1(n_1140),
.A2(n_1190),
.B1(n_1087),
.B2(n_1072),
.C1(n_1184),
.C2(n_1167),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1136),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1078),
.B(n_1050),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_1166),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_1172),
.B1(n_1189),
.B2(n_1188),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1080),
.A2(n_1067),
.B(n_1090),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1105),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1162),
.A2(n_1073),
.B1(n_1100),
.B2(n_1115),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1166),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1066),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1066),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1086),
.A2(n_1123),
.B(n_1109),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1138),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1180),
.B(n_1079),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1079),
.B(n_1134),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1066),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1074),
.B(n_1118),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1056),
.B(n_1144),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1068),
.A2(n_1089),
.B1(n_1118),
.B2(n_1141),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1096),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1065),
.A2(n_1093),
.B(n_1104),
.C(n_1102),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1051),
.A2(n_1060),
.B1(n_1108),
.B2(n_1088),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1085),
.A2(n_1098),
.B(n_1107),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1096),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1076),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1076),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1074),
.A2(n_1088),
.B1(n_1185),
.B2(n_1164),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1107),
.A2(n_1069),
.B(n_1153),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1129),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1137),
.A2(n_1159),
.B(n_1097),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1076),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1048),
.A2(n_1187),
.B(n_1186),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1065),
.A2(n_1092),
.B(n_1093),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1088),
.B(n_1075),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1152),
.Y(n_1245)
);

OAI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1102),
.A2(n_1101),
.B(n_1106),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1113),
.B(n_1049),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1117),
.A2(n_1111),
.B1(n_1131),
.B2(n_1178),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1148),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1148),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1103),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1131),
.B(n_1139),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1076),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1131),
.B(n_1157),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_1051),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1152),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1173),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1095),
.B(n_1124),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1135),
.A2(n_1156),
.B1(n_1139),
.B2(n_1157),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1060),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1104),
.B(n_1119),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1132),
.A2(n_1158),
.B(n_1133),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1135),
.B(n_1156),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1135),
.B(n_1178),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1052),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1139),
.B(n_1156),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1071),
.A2(n_1151),
.B(n_1181),
.Y(n_1268)
);

BUFx4_ASAP7_75t_SL g1269 ( 
.A(n_1173),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1157),
.A2(n_1178),
.B1(n_1127),
.B2(n_1095),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1083),
.A2(n_1110),
.B1(n_1121),
.B2(n_1127),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1095),
.B(n_1110),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1120),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1125),
.B(n_1095),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1128),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1112),
.A2(n_1094),
.B(n_1082),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1128),
.Y(n_1277)
);

NOR2xp67_ASAP7_75t_L g1278 ( 
.A(n_1143),
.B(n_1182),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1169),
.A2(n_1182),
.A3(n_1179),
.B(n_1175),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1122),
.A2(n_1179),
.B(n_1175),
.C(n_1169),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1128),
.B(n_1122),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1095),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1077),
.A2(n_1063),
.B(n_1122),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1128),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1122),
.B(n_1095),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1116),
.B(n_1099),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1055),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1105),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1072),
.B(n_777),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1050),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1057),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1055),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1066),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1055),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1058),
.A2(n_1062),
.B(n_983),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1055),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1300)
);

INVx4_ASAP7_75t_SL g1301 ( 
.A(n_1128),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1055),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1049),
.B(n_964),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1064),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1055),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1066),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1057),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1064),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1058),
.A2(n_1062),
.B1(n_1017),
.B2(n_1025),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1057),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1055),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1064),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1057),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1058),
.A2(n_1062),
.B1(n_1017),
.B2(n_1025),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1105),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1053),
.A2(n_1058),
.B1(n_950),
.B2(n_883),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1064),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1105),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1055),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1130),
.A2(n_1155),
.B1(n_1150),
.B2(n_1053),
.C(n_783),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1062),
.A2(n_1058),
.B(n_1057),
.Y(n_1330)
);

CKINVDCx6p67_ASAP7_75t_R g1331 ( 
.A(n_1166),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1048),
.A2(n_1133),
.B(n_1132),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1055),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1255),
.B(n_1256),
.Y(n_1335)
);

BUFx2_ASAP7_75t_R g1336 ( 
.A(n_1219),
.Y(n_1336)
);

INVx8_ASAP7_75t_L g1337 ( 
.A(n_1261),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1329),
.A2(n_1321),
.B1(n_1200),
.B2(n_1314),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1212),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1223),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1216),
.A2(n_1283),
.B(n_1222),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1198),
.B(n_1299),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1255),
.B(n_1256),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1242),
.A2(n_1332),
.B(n_1263),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1262),
.A2(n_1319),
.B1(n_1334),
.B2(n_1322),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1262),
.A2(n_1296),
.B1(n_1325),
.B2(n_1289),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1305),
.B(n_1310),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1300),
.A2(n_1328),
.B1(n_1206),
.B2(n_1297),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1255),
.B(n_1307),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1224),
.B(n_1291),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1287),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1201),
.B(n_1191),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1279),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1329),
.A2(n_1321),
.B1(n_1211),
.B2(n_1191),
.Y(n_1355)
);

INVx6_ASAP7_75t_L g1356 ( 
.A(n_1309),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1290),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1230),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1213),
.Y(n_1359)
);

BUFx4f_ASAP7_75t_L g1360 ( 
.A(n_1331),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1202),
.A2(n_1205),
.B1(n_1199),
.B2(n_1231),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1293),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1295),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1208),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1298),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1209),
.A2(n_1243),
.B1(n_1246),
.B2(n_1218),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1292),
.A2(n_1330),
.B(n_1312),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1302),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1235),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1308),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1316),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1327),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1214),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1333),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1209),
.A2(n_1243),
.B1(n_1248),
.B2(n_1237),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1231),
.A2(n_1193),
.B1(n_1330),
.B2(n_1318),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1215),
.A2(n_1204),
.B(n_1228),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1251),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1235),
.Y(n_1379)
);

CKINVDCx6p67_ASAP7_75t_R g1380 ( 
.A(n_1234),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1248),
.A2(n_1237),
.B1(n_1227),
.B2(n_1225),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1216),
.A2(n_1283),
.B(n_1222),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1232),
.A2(n_1247),
.B1(n_1270),
.B2(n_1303),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1267),
.A2(n_1193),
.B1(n_1252),
.B2(n_1254),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1264),
.B(n_1267),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1315),
.A2(n_1318),
.B1(n_1240),
.B2(n_1238),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1197),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1217),
.B(n_1324),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1282),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1239),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1210),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1239),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1244),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1260),
.A2(n_1264),
.B1(n_1228),
.B2(n_1265),
.Y(n_1395)
);

INVx4_ASAP7_75t_SL g1396 ( 
.A(n_1277),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1306),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1240),
.A2(n_1238),
.B1(n_1229),
.B2(n_1317),
.Y(n_1398)
);

NOR2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1257),
.B(n_1313),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1285),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1278),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1234),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1284),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1303),
.A2(n_1196),
.B1(n_1260),
.B2(n_1271),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1324),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1207),
.B(n_1323),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1192),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1192),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1220),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1288),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1288),
.Y(n_1411)
);

BUFx4f_ASAP7_75t_SL g1412 ( 
.A(n_1208),
.Y(n_1412)
);

BUFx8_ASAP7_75t_SL g1413 ( 
.A(n_1249),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1273),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1276),
.A2(n_1280),
.B(n_1233),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1320),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1320),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1303),
.A2(n_1196),
.B1(n_1326),
.B2(n_1304),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1269),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1274),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1250),
.A2(n_1258),
.B1(n_1304),
.B2(n_1326),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1236),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1236),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1203),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1241),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1274),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1266),
.A2(n_1272),
.B(n_1259),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1268),
.A2(n_1273),
.B(n_1266),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1281),
.A2(n_1275),
.B1(n_1301),
.B2(n_1259),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1241),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1221),
.B(n_1311),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1280),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1253),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1301),
.A2(n_1245),
.B1(n_1294),
.B2(n_1226),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1290),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1329),
.A2(n_1053),
.B1(n_1058),
.B2(n_783),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1255),
.B(n_1256),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1200),
.B(n_1058),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1195),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1194),
.A2(n_1085),
.B(n_1069),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1208),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1235),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1261),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1195),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1234),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1262),
.A2(n_783),
.B1(n_372),
.B2(n_383),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1329),
.A2(n_783),
.B1(n_730),
.B2(n_905),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1329),
.A2(n_1053),
.B1(n_1058),
.B2(n_783),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1195),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1195),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1242),
.A2(n_1332),
.B(n_1263),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1282),
.Y(n_1452)
);

CKINVDCx6p67_ASAP7_75t_R g1453 ( 
.A(n_1402),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1403),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1391),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1400),
.B(n_1420),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1393),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1402),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1344),
.A2(n_1451),
.B(n_1367),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1378),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1432),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1390),
.B(n_1426),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1445),
.Y(n_1463)
);

AND2x6_ASAP7_75t_L g1464 ( 
.A(n_1335),
.B(n_1404),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1427),
.Y(n_1465)
);

AO31x2_ASAP7_75t_L g1466 ( 
.A1(n_1376),
.A2(n_1377),
.A3(n_1386),
.B(n_1354),
.Y(n_1466)
);

AOI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1438),
.A2(n_1366),
.B(n_1447),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1359),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1350),
.B(n_1394),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1339),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1340),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1351),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1414),
.Y(n_1473)
);

INVxp33_ASAP7_75t_L g1474 ( 
.A(n_1413),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1362),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1451),
.A2(n_1428),
.B(n_1392),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1363),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1365),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1368),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1414),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1346),
.B(n_1345),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1370),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1440),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1413),
.B(n_1406),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1374),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1439),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1415),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1444),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1411),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1436),
.A2(n_1448),
.B(n_1338),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1384),
.B(n_1348),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1342),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1384),
.B(n_1347),
.Y(n_1495)
);

INVxp33_ASAP7_75t_L g1496 ( 
.A(n_1424),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1353),
.B(n_1375),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1353),
.B(n_1375),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1405),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1430),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1381),
.B(n_1357),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1361),
.B(n_1338),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1503)
);

NOR2x1_ASAP7_75t_SL g1504 ( 
.A(n_1398),
.B(n_1379),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1452),
.A2(n_1382),
.B(n_1341),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1452),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1436),
.A2(n_1448),
.B(n_1355),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1397),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1341),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1405),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1383),
.A2(n_1401),
.B(n_1387),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1382),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1407),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1408),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1429),
.B(n_1382),
.Y(n_1515)
);

BUFx4f_ASAP7_75t_SL g1516 ( 
.A(n_1380),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1435),
.B(n_1355),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1381),
.B(n_1429),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1395),
.B(n_1410),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1434),
.A2(n_1425),
.B(n_1417),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1446),
.A2(n_1395),
.B(n_1421),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1416),
.B(n_1425),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1423),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1423),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1433),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1433),
.B(n_1352),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1515),
.B(n_1422),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1497),
.B(n_1383),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1515),
.B(n_1422),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1466),
.B(n_1422),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1469),
.B(n_1380),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1454),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1483),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1500),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1454),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1460),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1491),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1498),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1467),
.B(n_1405),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1509),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1466),
.B(n_1369),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1466),
.B(n_1369),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1466),
.B(n_1369),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1507),
.A2(n_1418),
.B1(n_1337),
.B2(n_1441),
.C(n_1364),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1465),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1492),
.A2(n_1356),
.B1(n_1443),
.B2(n_1337),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1509),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1465),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1388),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1500),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1456),
.B(n_1385),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1455),
.B(n_1409),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1455),
.B(n_1457),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1488),
.B(n_1399),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1502),
.B(n_1424),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1481),
.A2(n_1409),
.B1(n_1419),
.B2(n_1437),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1483),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1457),
.B(n_1431),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1476),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1521),
.A2(n_1443),
.B1(n_1360),
.B2(n_1349),
.C(n_1343),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1513),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1558),
.B(n_1496),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1528),
.A2(n_1518),
.B1(n_1493),
.B2(n_1501),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1551),
.B(n_1456),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_SL g1568 ( 
.A(n_1558),
.B(n_1493),
.C(n_1545),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1538),
.B(n_1468),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1539),
.A2(n_1517),
.B(n_1508),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1539),
.A2(n_1520),
.B(n_1519),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1564),
.B(n_1514),
.C(n_1501),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1473),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1534),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1529),
.B(n_1480),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1528),
.A2(n_1518),
.B1(n_1453),
.B2(n_1494),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1541),
.A2(n_1474),
.B(n_1484),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1537),
.B(n_1519),
.C(n_1523),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1504),
.B(n_1506),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1541),
.A2(n_1543),
.B(n_1542),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1534),
.B(n_1553),
.C(n_1533),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1541),
.B(n_1542),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1562),
.A2(n_1505),
.B(n_1459),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1559),
.B(n_1545),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1544),
.B(n_1523),
.C(n_1524),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1555),
.B(n_1458),
.C(n_1373),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_SL g1588 ( 
.A(n_1559),
.B(n_1373),
.C(n_1490),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1543),
.B(n_1506),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1470),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1470),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1530),
.A2(n_1503),
.B(n_1526),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1563),
.B(n_1499),
.C(n_1510),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1557),
.A2(n_1511),
.B1(n_1464),
.B2(n_1462),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1556),
.B(n_1471),
.Y(n_1595)
);

NOR2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1531),
.B(n_1453),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1471),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1544),
.B(n_1524),
.C(n_1461),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1546),
.B(n_1461),
.C(n_1478),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1522),
.C(n_1482),
.D(n_1479),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1547),
.A2(n_1487),
.B1(n_1482),
.B2(n_1479),
.C(n_1478),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1546),
.B(n_1477),
.C(n_1475),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1530),
.A2(n_1503),
.B(n_1526),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1533),
.B(n_1525),
.C(n_1522),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1532),
.B(n_1472),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1557),
.A2(n_1511),
.B1(n_1464),
.B2(n_1462),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1532),
.B(n_1472),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1530),
.A2(n_1489),
.B(n_1477),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_1475),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1535),
.B(n_1486),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1536),
.B(n_1486),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1583),
.B(n_1540),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1605),
.Y(n_1613)
);

OAI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1578),
.A2(n_1580),
.B(n_1572),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1574),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1607),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1569),
.B(n_1554),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1609),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1567),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1610),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1584),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1608),
.B(n_1547),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1568),
.A2(n_1548),
.B1(n_1464),
.B2(n_1552),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1611),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_L g1630 ( 
.A(n_1586),
.B(n_1549),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1595),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1567),
.B(n_1581),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1589),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1597),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1608),
.B(n_1550),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1591),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1573),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1572),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1639),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1613),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1614),
.A2(n_1570),
.B1(n_1585),
.B2(n_1578),
.C(n_1571),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1632),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1614),
.A2(n_1600),
.B(n_1582),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1643),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1633),
.B(n_1577),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1621),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1601),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1639),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1618),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1620),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1638),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1620),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1638),
.B(n_1598),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1616),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1641),
.B(n_1550),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1621),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1616),
.B(n_1579),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1536),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1621),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1531),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1622),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1463),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1623),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1615),
.B(n_1575),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1625),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1625),
.Y(n_1674)
);

NAND2x1_ASAP7_75t_L g1675 ( 
.A(n_1616),
.B(n_1560),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1629),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1628),
.A2(n_1566),
.B1(n_1576),
.B2(n_1594),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1617),
.B(n_1531),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1627),
.B(n_1588),
.C(n_1565),
.Y(n_1680)
);

NAND2x1_ASAP7_75t_SL g1681 ( 
.A(n_1644),
.B(n_1616),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1648),
.B(n_1651),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1661),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1670),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1654),
.B(n_1631),
.Y(n_1685)
);

NOR5xp2_ASAP7_75t_L g1686 ( 
.A(n_1676),
.B(n_1603),
.C(n_1592),
.D(n_1631),
.E(n_1634),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1617),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1649),
.B(n_1615),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1668),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1645),
.B(n_1634),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1661),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1656),
.B(n_1636),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1650),
.B(n_1636),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1652),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1612),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1646),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1646),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1612),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1637),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1661),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1647),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1653),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1665),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1647),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1663),
.B(n_1637),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1666),
.B(n_1619),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1650),
.B(n_1629),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1659),
.B(n_1612),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1679),
.B(n_1624),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1655),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1679),
.B(n_1624),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1653),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1653),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1644),
.A2(n_1628),
.B1(n_1624),
.B2(n_1627),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1655),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1657),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1668),
.B(n_1463),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1657),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1658),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1644),
.B(n_1635),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1678),
.A2(n_1635),
.B1(n_1606),
.B2(n_1596),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1698),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1704),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1699),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1689),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1704),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1724),
.A2(n_1678),
.B1(n_1680),
.B2(n_1659),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1709),
.B(n_1666),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1704),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1694),
.B(n_1659),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1708),
.B(n_1660),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1715),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1683),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1660),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_1720),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1694),
.B(n_1659),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1682),
.A2(n_1665),
.B1(n_1662),
.B2(n_1675),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1673),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1699),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1685),
.B(n_1687),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1703),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1715),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1690),
.B(n_1673),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1681),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1674),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1681),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1701),
.B(n_1674),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1706),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1706),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1707),
.B(n_1677),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1716),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1707),
.B(n_1692),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1662),
.C(n_1675),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1731),
.A2(n_1717),
.B1(n_1705),
.B2(n_1723),
.C(n_1683),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1753),
.B(n_1695),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1725),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1729),
.B(n_1695),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1725),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1751),
.A2(n_1717),
.B1(n_1683),
.B2(n_1697),
.C(n_1702),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_L g1768 ( 
.A1(n_1753),
.A2(n_1697),
.B(n_1691),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1728),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1760),
.A2(n_1711),
.B1(n_1684),
.B2(n_1686),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1743),
.A2(n_1691),
.B(n_1697),
.C(n_1702),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1745),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1734),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1746),
.A2(n_1711),
.B1(n_1702),
.B2(n_1691),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1745),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1735),
.A2(n_1732),
.B1(n_1730),
.B2(n_1726),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1740),
.B(n_1711),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1747),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1734),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1759),
.B(n_1700),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1726),
.A2(n_1716),
.B(n_1667),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1735),
.Y(n_1783)
);

AOI332xp33_ASAP7_75t_L g1784 ( 
.A1(n_1747),
.A2(n_1711),
.A3(n_1721),
.B1(n_1719),
.B2(n_1718),
.B3(n_1722),
.C1(n_1713),
.C2(n_1700),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1755),
.B(n_1713),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1744),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1781),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1776),
.B(n_1759),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_1732),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1766),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1766),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1763),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1762),
.Y(n_1793)
);

NOR3x1_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1750),
.C(n_1748),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1762),
.Y(n_1795)
);

NAND2x1_ASAP7_75t_L g1796 ( 
.A(n_1762),
.B(n_1741),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1776),
.B(n_1785),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1777),
.B(n_1741),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1736),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1765),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1786),
.B(n_1736),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1773),
.B(n_1688),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1780),
.B(n_1739),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1773),
.B(n_1739),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1772),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1797),
.A2(n_1770),
.B1(n_1767),
.B2(n_1774),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1795),
.B(n_1779),
.Y(n_1808)
);

OAI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1797),
.A2(n_1784),
.B(n_1771),
.C(n_1764),
.Y(n_1809)
);

AOI222xp33_ASAP7_75t_L g1810 ( 
.A1(n_1788),
.A2(n_1775),
.B1(n_1778),
.B2(n_1733),
.C1(n_1730),
.C2(n_1737),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1789),
.A2(n_1768),
.B1(n_1755),
.B2(n_1756),
.C(n_1758),
.Y(n_1811)
);

OAI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1798),
.A2(n_1779),
.B(n_1727),
.Y(n_1812)
);

NAND4xp25_ASAP7_75t_L g1813 ( 
.A(n_1794),
.B(n_1756),
.C(n_1710),
.D(n_1757),
.Y(n_1813)
);

O2A1O1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1787),
.A2(n_1752),
.B(n_1754),
.C(n_1757),
.Y(n_1814)
);

AND5x1_ASAP7_75t_L g1815 ( 
.A(n_1801),
.B(n_1593),
.C(n_1782),
.D(n_1737),
.E(n_1749),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1796),
.A2(n_1782),
.B(n_1754),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1793),
.B(n_1752),
.C(n_1742),
.Y(n_1817)
);

OAI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1795),
.A2(n_1710),
.B(n_1714),
.C(n_1712),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1805),
.A2(n_1782),
.B1(n_1758),
.B2(n_1749),
.C(n_1742),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1809),
.A2(n_1793),
.B1(n_1804),
.B2(n_1799),
.Y(n_1820)
);

NAND4xp75_ASAP7_75t_SL g1821 ( 
.A(n_1807),
.B(n_1802),
.C(n_1688),
.D(n_1696),
.Y(n_1821)
);

AO22x2_ASAP7_75t_L g1822 ( 
.A1(n_1817),
.A2(n_1806),
.B1(n_1803),
.B2(n_1800),
.Y(n_1822)
);

NOR4xp75_ASAP7_75t_L g1823 ( 
.A(n_1808),
.B(n_1793),
.C(n_1792),
.D(n_1791),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1810),
.B(n_1812),
.Y(n_1824)
);

NOR3xp33_ASAP7_75t_L g1825 ( 
.A(n_1819),
.B(n_1790),
.C(n_1733),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1814),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_L g1827 ( 
.A(n_1811),
.B(n_1816),
.C(n_1813),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1818),
.A2(n_1716),
.B1(n_1669),
.B2(n_1664),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1815),
.B(n_1719),
.C(n_1718),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1826),
.B(n_1336),
.Y(n_1830)
);

AOI211xp5_ASAP7_75t_L g1831 ( 
.A1(n_1827),
.A2(n_1824),
.B(n_1820),
.C(n_1825),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_1721),
.Y(n_1832)
);

OAI21xp33_ASAP7_75t_L g1833 ( 
.A1(n_1822),
.A2(n_1722),
.B(n_1587),
.Y(n_1833)
);

NAND4xp25_ASAP7_75t_SL g1834 ( 
.A(n_1821),
.B(n_1696),
.C(n_1516),
.D(n_1640),
.Y(n_1834)
);

NOR3xp33_ASAP7_75t_L g1835 ( 
.A(n_1828),
.B(n_1823),
.C(n_1667),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1830),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1832),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1834),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1835),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1833),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1831),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1830),
.A2(n_1664),
.B1(n_1667),
.B2(n_1669),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1841),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1840),
.B(n_1360),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1837),
.B(n_1672),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1838),
.B(n_1672),
.Y(n_1846)
);

OAI21xp33_ASAP7_75t_L g1847 ( 
.A1(n_1836),
.A2(n_1677),
.B(n_1669),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1839),
.B(n_1842),
.Y(n_1848)
);

AND3x1_ASAP7_75t_L g1849 ( 
.A(n_1844),
.B(n_1358),
.C(n_1412),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1845),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1846),
.B(n_1596),
.Y(n_1851)
);

NAND4xp75_ASAP7_75t_L g1852 ( 
.A(n_1849),
.B(n_1843),
.C(n_1848),
.D(n_1847),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1852),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1853),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1853),
.A2(n_1850),
.B(n_1851),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1855),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1855),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1857),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1856),
.A2(n_1854),
.B1(n_1855),
.B2(n_1851),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1858),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1859),
.B1(n_1358),
.B2(n_1664),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_R g1862 ( 
.A1(n_1861),
.A2(n_1358),
.B1(n_1337),
.B2(n_1548),
.C(n_1640),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1622),
.B(n_1626),
.C(n_1337),
.Y(n_1863)
);


endmodule