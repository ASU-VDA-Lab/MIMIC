module fake_jpeg_24503_n_39 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_6),
.B(n_2),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_5),
.A2(n_3),
.B1(n_6),
.B2(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_8),
.A2(n_0),
.B1(n_4),
.B2(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_4),
.B2(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_0),
.B1(n_13),
.B2(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_25),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_19),
.B(n_24),
.C(n_23),
.D(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_36),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_37),
.C(n_35),
.Y(n_39)
);


endmodule