module fake_netlist_1_7399_n_746 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_746);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_746;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_395;
wire n_132;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_15), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_54), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_19), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_78), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_34), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_53), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_58), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_80), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_27), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_16), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_17), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_36), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_38), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_69), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_29), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_4), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_76), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_33), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_48), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_57), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_23), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_44), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_41), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_72), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_14), .Y(n_124) );
CKINVDCx14_ASAP7_75t_R g125 ( .A(n_24), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_16), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_45), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_65), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_42), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_1), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_111), .Y(n_131) );
BUFx8_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_111), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_130), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_90), .Y(n_145) );
BUFx8_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_109), .B(n_0), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_96), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_98), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_116), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_88), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_93), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_89), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_83), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_81), .B(n_32), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_92), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_94), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_99), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_92), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_103), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
XNOR2xp5_ASAP7_75t_L g171 ( .A(n_117), .B(n_0), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_103), .B(n_2), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_99), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_102), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_107), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_152), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_155), .B(n_87), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_138), .B(n_95), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_172), .Y(n_182) );
OAI221xp5_ASAP7_75t_L g183 ( .A1(n_158), .A2(n_124), .B1(n_121), .B2(n_104), .C(n_126), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_124), .B1(n_121), .B2(n_104), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_168), .B(n_113), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_168), .B(n_113), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_146), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_158), .B(n_126), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_139), .B(n_115), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_139), .B(n_115), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_145), .B(n_95), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_140), .B(n_118), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_172), .B(n_112), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_147), .B(n_112), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_142), .B(n_110), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
AND2x4_ASAP7_75t_SL g214 ( .A(n_147), .B(n_110), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_136), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_140), .B(n_127), .Y(n_217) );
AND2x6_ASAP7_75t_L g218 ( .A(n_147), .B(n_114), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_163), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_141), .B(n_108), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_141), .B(n_108), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_143), .B(n_114), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_143), .B(n_119), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_163), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_132), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
AND2x6_ASAP7_75t_L g232 ( .A(n_149), .B(n_119), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_134), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_133), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_149), .B(n_128), .Y(n_236) );
INVx6_ASAP7_75t_L g237 ( .A(n_132), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_154), .B(n_128), .Y(n_238) );
INVxp33_ASAP7_75t_L g239 ( .A(n_142), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_160), .B(n_85), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_134), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_136), .A2(n_169), .B1(n_164), .B2(n_144), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_160), .B(n_106), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_187), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_190), .B(n_154), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_210), .A2(n_159), .B1(n_167), .B2(n_166), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g247 ( .A(n_201), .B(n_148), .C(n_150), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_211), .B(n_159), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
OR2x2_ASAP7_75t_SL g251 ( .A(n_177), .B(n_153), .Y(n_251) );
OR2x2_ASAP7_75t_SL g252 ( .A(n_237), .B(n_242), .Y(n_252) );
BUFx12f_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
CKINVDCx8_ASAP7_75t_R g254 ( .A(n_198), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_211), .B(n_167), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_211), .B(n_193), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_222), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_241), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_237), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_237), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_230), .Y(n_264) );
XNOR2x2_ASAP7_75t_SL g265 ( .A(n_184), .B(n_171), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_230), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_190), .A2(n_162), .B(n_157), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_231), .Y(n_268) );
NOR2xp33_ASAP7_75t_R g269 ( .A(n_187), .B(n_131), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_193), .B(n_157), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_205), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_239), .B(n_135), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_216), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_196), .B(n_166), .Y(n_275) );
INVx3_ASAP7_75t_SL g276 ( .A(n_221), .Y(n_276) );
INVx4_ASAP7_75t_L g277 ( .A(n_192), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_196), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_235), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_181), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_222), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_196), .B(n_165), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_192), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_202), .B(n_165), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_183), .B(n_174), .C(n_156), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_205), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_235), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_202), .B(n_123), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_243), .B(n_171), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_182), .B(n_100), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_186), .B(n_133), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_203), .B(n_133), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_240), .B(n_133), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_206), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_186), .B(n_137), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_234), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_234), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_217), .B(n_137), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_186), .Y(n_301) );
AOI22xp5_ASAP7_75t_SL g302 ( .A1(n_207), .A2(n_129), .B1(n_122), .B2(n_123), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_189), .B(n_105), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_189), .B(n_105), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_205), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_210), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_234), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_189), .B(n_101), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_205), .Y(n_309) );
BUFx6f_ASAP7_75t_SL g310 ( .A(n_210), .Y(n_310) );
OAI22xp5_ASAP7_75t_SL g311 ( .A1(n_180), .A2(n_100), .B1(n_101), .B2(n_6), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_234), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_205), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_214), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_227), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_214), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_315), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_315), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_258), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_248), .B(n_210), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_308), .A2(n_218), .B1(n_210), .B2(n_205), .Y(n_322) );
BUFx12f_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_305), .B(n_182), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_248), .B(n_210), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_248), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_305), .B(n_195), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_283), .B(n_240), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_278), .A2(n_218), .B1(n_243), .B2(n_195), .Y(n_330) );
BUFx2_ASAP7_75t_R g331 ( .A(n_254), .Y(n_331) );
BUFx4f_ASAP7_75t_SL g332 ( .A(n_276), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_313), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_308), .A2(n_256), .B1(n_246), .B2(n_255), .Y(n_335) );
OR2x6_ASAP7_75t_L g336 ( .A(n_308), .B(n_204), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_263), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_244), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_268), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_218), .B1(n_204), .B2(n_232), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_291), .B(n_206), .Y(n_341) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_313), .B(n_204), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_244), .Y(n_343) );
INVx2_ASAP7_75t_R g344 ( .A(n_271), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_279), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_245), .A2(n_194), .B(n_236), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_276), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_283), .B(n_206), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_275), .B(n_218), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_271), .B(n_194), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_250), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_250), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_273), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_310), .A2(n_194), .B1(n_238), .B2(n_225), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_267), .A2(n_224), .B(n_223), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_284), .B(n_220), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_306), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_280), .A2(n_218), .B1(n_232), .B2(n_226), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_272), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_304), .A2(n_213), .B(n_228), .C(n_229), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_301), .B(n_218), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_259), .B(n_274), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_297), .B(n_220), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_259), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_250), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_271), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_316), .A2(n_226), .B1(n_232), .B2(n_220), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_264), .A2(n_226), .B1(n_232), .B2(n_228), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_296), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_298), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_297), .B(n_226), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_323), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_323), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_317), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_293), .B1(n_310), .B2(n_297), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_362), .A2(n_300), .B(n_294), .C(n_270), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_322), .B(n_310), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_332), .Y(n_381) );
CKINVDCx11_ASAP7_75t_R g382 ( .A(n_319), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_328), .A2(n_293), .B1(n_311), .B2(n_303), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_329), .B(n_293), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_317), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_336), .B(n_271), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_346), .A2(n_245), .B(n_284), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_328), .A2(n_266), .B1(n_264), .B2(n_226), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_336), .B(n_271), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_336), .A2(n_254), .B1(n_266), .B2(n_265), .Y(n_392) );
AOI221x1_ASAP7_75t_SL g393 ( .A1(n_320), .A2(n_252), .B1(n_247), .B2(n_251), .C(n_208), .Y(n_393) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_290), .B(n_302), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_333), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_329), .B(n_349), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_333), .A2(n_286), .B(n_292), .C(n_229), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_327), .A2(n_226), .B1(n_232), .B2(n_292), .Y(n_398) );
NAND3xp33_ASAP7_75t_SL g399 ( .A(n_361), .B(n_269), .C(n_295), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_349), .B(n_232), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_340), .B(n_259), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_354), .B(n_290), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_318), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_336), .B(n_260), .Y(n_405) );
NAND2xp33_ASAP7_75t_SL g406 ( .A(n_324), .B(n_269), .Y(n_406) );
AOI221x1_ASAP7_75t_L g407 ( .A1(n_335), .A2(n_176), .B1(n_200), .B2(n_197), .C(n_188), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_374), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_379), .B(n_337), .Y(n_411) );
OAI322xp33_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_341), .A3(n_330), .B1(n_339), .B2(n_345), .C1(n_348), .C2(n_233), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_383), .A2(n_327), .B1(n_363), .B2(n_347), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_393), .A2(n_341), .B1(n_345), .B2(n_348), .C(n_339), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_394), .A2(n_347), .B1(n_355), .B2(n_321), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
OAI22xp33_ASAP7_75t_SL g419 ( .A1(n_403), .A2(n_364), .B1(n_331), .B2(n_360), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_388), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
BUFx4f_ASAP7_75t_SL g422 ( .A(n_386), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_365), .B1(n_350), .B2(n_326), .C(n_185), .Y(n_423) );
OA21x2_ASAP7_75t_L g424 ( .A1(n_407), .A2(n_357), .B(n_378), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_408), .B(n_371), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_388), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_394), .A2(n_365), .B1(n_359), .B2(n_352), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
OAI21x1_ASAP7_75t_L g429 ( .A1(n_407), .A2(n_357), .B(n_372), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_370), .B1(n_364), .B2(n_359), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_380), .A2(n_352), .B1(n_367), .B2(n_371), .Y(n_432) );
CKINVDCx11_ASAP7_75t_R g433 ( .A(n_382), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_376), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_387), .B(n_185), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_396), .B(n_353), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_402), .A2(n_352), .B1(n_367), .B2(n_369), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_405), .A2(n_364), .B1(n_373), .B2(n_343), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_412), .A2(n_402), .B1(n_406), .B2(n_405), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_410), .B(n_384), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_414), .B(n_386), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_418), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_412), .A2(n_397), .B1(n_403), .B2(n_375), .C(n_381), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_418), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_418), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_415), .B(n_234), .C(n_191), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_422), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_411), .A2(n_405), .B1(n_386), .B2(n_364), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_414), .B(n_405), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_427), .A2(n_405), .B1(n_402), .B2(n_390), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_429), .A2(n_389), .B(n_401), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_438), .B(n_388), .Y(n_452) );
OAI33xp33_ASAP7_75t_L g453 ( .A1(n_419), .A2(n_219), .A3(n_191), .B1(n_212), .B2(n_199), .B3(n_208), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_411), .A2(n_400), .B1(n_401), .B2(n_404), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_430), .B(n_387), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_415), .B(n_215), .C(n_199), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_430), .B(n_387), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_433), .Y(n_459) );
OAI21x1_ASAP7_75t_L g460 ( .A1(n_429), .A2(n_404), .B(n_401), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_434), .B(n_404), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_409), .A2(n_413), .B1(n_416), .B2(n_437), .Y(n_462) );
OAI21x1_ASAP7_75t_L g463 ( .A1(n_429), .A2(n_372), .B(n_368), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_435), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
OAI33xp33_ASAP7_75t_L g466 ( .A1(n_419), .A2(n_212), .A3(n_215), .B1(n_219), .B2(n_233), .B3(n_227), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_438), .B(n_388), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_423), .A2(n_377), .B1(n_353), .B2(n_367), .C(n_391), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_423), .A2(n_391), .B1(n_338), .B2(n_343), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_436), .B(n_398), .C(n_209), .D(n_179), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_420), .B(n_391), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_434), .B(n_391), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
NAND2xp33_ASAP7_75t_R g475 ( .A(n_426), .B(n_3), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_461), .Y(n_476) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_475), .B(n_420), .Y(n_477) );
AOI33xp33_ASAP7_75t_L g478 ( .A1(n_469), .A2(n_428), .A3(n_421), .B1(n_431), .B2(n_432), .B3(n_209), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_455), .B(n_421), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_461), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_464), .B(n_428), .Y(n_482) );
AND3x2_ASAP7_75t_L g483 ( .A(n_441), .B(n_425), .C(n_5), .Y(n_483) );
OAI31xp33_ASAP7_75t_L g484 ( .A1(n_448), .A2(n_425), .A3(n_426), .B(n_338), .Y(n_484) );
AND3x1_ASAP7_75t_L g485 ( .A(n_443), .B(n_426), .C(n_5), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_457), .Y(n_486) );
OAI31xp33_ASAP7_75t_L g487 ( .A1(n_450), .A2(n_426), .A3(n_285), .B(n_262), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_470), .B(n_424), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g489 ( .A1(n_462), .A2(n_3), .B1(n_6), .B2(n_7), .C1(n_8), .C2(n_9), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_455), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_458), .B(n_424), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_446), .B(n_449), .C(n_439), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_470), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_452), .B(n_424), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_473), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_465), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_452), .A2(n_424), .B1(n_366), .B2(n_358), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_460), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
AOI33xp33_ASAP7_75t_L g500 ( .A1(n_447), .A2(n_178), .A3(n_179), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_458), .B(n_7), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_452), .B(n_8), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_459), .B(n_11), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_453), .A2(n_176), .B1(n_188), .B2(n_197), .C(n_200), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_12), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_474), .B(n_12), .Y(n_512) );
AOI33xp33_ASAP7_75t_L g513 ( .A1(n_468), .A2(n_178), .A3(n_14), .B1(n_18), .B2(n_19), .B3(n_20), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_474), .B(n_13), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_467), .A2(n_366), .B1(n_262), .B2(n_277), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_451), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_467), .B(n_18), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_456), .A2(n_285), .B(n_342), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_467), .B(n_20), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_467), .B(n_77), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_440), .B(n_21), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_451), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_473), .B(n_22), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_472), .B(n_22), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_463), .Y(n_526) );
INVx4_ASAP7_75t_L g527 ( .A(n_472), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_476), .B(n_472), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_490), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_496), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_491), .B(n_472), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_496), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_476), .B(n_454), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_491), .B(n_25), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_506), .B(n_55), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_508), .B(n_459), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_480), .B(n_479), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_480), .B(n_25), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_481), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_479), .B(n_26), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_506), .B(n_61), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_481), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_486), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_501), .B(n_26), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_486), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_493), .B(n_197), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_504), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_493), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_197), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_482), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_482), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_501), .B(n_471), .Y(n_554) );
NAND4xp75_ASAP7_75t_L g555 ( .A(n_485), .B(n_466), .C(n_342), .D(n_37), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_520), .B(n_324), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_505), .Y(n_559) );
NAND3xp33_ASAP7_75t_SL g560 ( .A(n_489), .B(n_351), .C(n_277), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_488), .B(n_188), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_495), .B(n_188), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_488), .B(n_188), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
INVxp33_ASAP7_75t_L g565 ( .A(n_520), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_525), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_495), .B(n_197), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_502), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_512), .B(n_176), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_512), .B(n_176), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_489), .B(n_277), .C(n_324), .D(n_249), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_485), .A2(n_334), .B1(n_299), .B2(n_307), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_527), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_514), .B(n_200), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
OAI31xp33_ASAP7_75t_L g577 ( .A1(n_477), .A2(n_351), .A3(n_368), .B(n_334), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_527), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_519), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_494), .B(n_200), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_514), .B(n_200), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_520), .B(n_325), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_519), .Y(n_585) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_484), .A2(n_325), .B(n_287), .C(n_309), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_516), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_525), .B(n_176), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_494), .B(n_28), .Y(n_589) );
NOR2xp33_ASAP7_75t_R g590 ( .A(n_483), .B(n_30), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_560), .A2(n_522), .B(n_524), .C(n_487), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_582), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_553), .B(n_510), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_531), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_565), .A2(n_520), .B1(n_527), .B2(n_492), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_533), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_530), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_555), .A2(n_484), .B(n_500), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_557), .A2(n_487), .B(n_492), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_530), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_552), .B(n_510), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_538), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_573), .A2(n_497), .B1(n_527), .B2(n_515), .C(n_518), .Y(n_603) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_557), .A2(n_515), .B(n_507), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_540), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_532), .B(n_521), .Y(n_606) );
OR4x1_ASAP7_75t_L g607 ( .A(n_558), .B(n_521), .C(n_502), .D(n_503), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_556), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_535), .B(n_503), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_566), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_532), .B(n_523), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_569), .B(n_507), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_535), .B(n_478), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_564), .B(n_513), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_544), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_582), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_590), .B(n_516), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_547), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_576), .B(n_523), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_539), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_565), .A2(n_509), .B1(n_526), .B2(n_523), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_550), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_572), .A2(n_518), .B1(n_526), .B2(n_528), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_559), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_568), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_546), .A2(n_528), .B(n_499), .Y(n_627) );
OAI32xp33_ASAP7_75t_L g628 ( .A1(n_557), .A2(n_528), .A3(n_499), .B1(n_498), .B2(n_351), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_542), .A2(n_499), .B1(n_498), .B2(n_299), .C1(n_298), .C2(n_312), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_578), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_580), .B(n_498), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_585), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_554), .B(n_39), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_529), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_584), .A2(n_368), .B(n_287), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_555), .A2(n_309), .B(n_287), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_SL g637 ( .A1(n_537), .A2(n_334), .B(n_288), .C(n_282), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_577), .B(n_312), .C(n_298), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_529), .B(n_40), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_584), .A2(n_287), .B(n_309), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_586), .A2(n_287), .B(n_309), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_534), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_574), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_618), .A2(n_536), .B(n_543), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_605), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_624), .A2(n_574), .B1(n_579), .B2(n_589), .C(n_588), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_615), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_618), .B(n_543), .Y(n_650) );
XNOR2xp5_ASAP7_75t_L g651 ( .A(n_610), .B(n_589), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_600), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g653 ( .A1(n_641), .A2(n_536), .B(n_543), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_592), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_643), .B(n_587), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_597), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_602), .B(n_587), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_591), .A2(n_536), .B(n_579), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_613), .A2(n_549), .B1(n_541), .B2(n_581), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_638), .B(n_567), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_619), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_630), .B(n_556), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_644), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_611), .B(n_549), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_611), .B(n_541), .Y(n_666) );
NOR3xp33_ASAP7_75t_SL g667 ( .A(n_598), .B(n_583), .C(n_570), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_632), .B(n_548), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g669 ( .A1(n_595), .A2(n_581), .A3(n_541), .B(n_567), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_625), .B(n_563), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_623), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_599), .B(n_562), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_594), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_592), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_626), .B(n_563), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_621), .B(n_575), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g678 ( .A(n_606), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_634), .B(n_561), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_606), .B(n_561), .Y(n_680) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_603), .B(n_571), .C(n_46), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_593), .B(n_551), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_620), .B(n_551), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_604), .B(n_309), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_661), .A2(n_624), .B(n_622), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_659), .A2(n_614), .B1(n_645), .B2(n_627), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_678), .B(n_620), .Y(n_687) );
AND4x1_ASAP7_75t_L g688 ( .A(n_681), .B(n_629), .C(n_633), .D(n_636), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_647), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_678), .A2(n_609), .B1(n_612), .B2(n_608), .Y(n_690) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_657), .A2(n_622), .A3(n_608), .B1(n_601), .B2(n_631), .C1(n_639), .C2(n_616), .Y(n_691) );
NOR2x1p5_ASAP7_75t_SL g692 ( .A(n_655), .B(n_612), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_652), .B(n_616), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g694 ( .A1(n_648), .A2(n_628), .B(n_637), .C(n_607), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_646), .A2(n_637), .B(n_635), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_653), .A2(n_607), .B(n_640), .C(n_642), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_658), .B(n_43), .Y(n_697) );
NAND4xp75_ASAP7_75t_L g698 ( .A(n_669), .B(n_47), .C(n_49), .D(n_50), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_684), .A2(n_298), .B(n_312), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_650), .A2(n_344), .B(n_312), .C(n_307), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_655), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_664), .A2(n_307), .B1(n_299), .B2(n_344), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g703 ( .A(n_651), .B(n_344), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_647), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_672), .B(n_288), .C(n_282), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_649), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_660), .B(n_52), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_651), .B(n_62), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_689), .Y(n_709) );
NOR2x1p5_ASAP7_75t_L g710 ( .A(n_698), .B(n_682), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_687), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_704), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_685), .B(n_677), .C(n_663), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_686), .B(n_671), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_696), .A2(n_667), .B(n_649), .C(n_654), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_703), .A2(n_656), .B(n_683), .Y(n_716) );
NAND4xp75_ASAP7_75t_L g717 ( .A(n_692), .B(n_670), .C(n_680), .D(n_666), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_691), .B(n_671), .C(n_662), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_690), .A2(n_673), .B1(n_662), .B2(n_654), .C(n_674), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_694), .A2(n_676), .B(n_668), .C(n_674), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_695), .B(n_673), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_708), .B(n_675), .Y(n_722) );
AOI211xp5_ASAP7_75t_L g723 ( .A1(n_700), .A2(n_680), .B(n_666), .C(n_665), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_693), .A2(n_665), .B1(n_679), .B2(n_675), .C(n_307), .Y(n_724) );
NOR4xp25_ASAP7_75t_L g725 ( .A(n_700), .B(n_281), .C(n_257), .D(n_249), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_705), .A2(n_299), .B1(n_281), .B2(n_257), .Y(n_726) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_706), .A2(n_63), .B1(n_64), .B2(n_66), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_701), .B(n_67), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_707), .A2(n_71), .B1(n_74), .B2(n_75), .Y(n_729) );
BUFx2_ASAP7_75t_L g730 ( .A(n_701), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_701), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_705), .Y(n_732) );
OAI322xp33_ASAP7_75t_L g733 ( .A1(n_715), .A2(n_714), .A3(n_722), .B1(n_718), .B2(n_711), .C1(n_716), .C2(n_732), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_730), .Y(n_734) );
AOI211xp5_ASAP7_75t_L g735 ( .A1(n_720), .A2(n_721), .B(n_719), .C(n_724), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_721), .A2(n_713), .B1(n_717), .B2(n_710), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g737 ( .A1(n_719), .A2(n_712), .B1(n_709), .B2(n_731), .C1(n_728), .C2(n_723), .Y(n_737) );
AND3x1_ASAP7_75t_L g738 ( .A(n_736), .B(n_725), .C(n_699), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_737), .A2(n_727), .B1(n_729), .B2(n_702), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_735), .B(n_688), .C(n_697), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_740), .Y(n_741) );
OR3x1_ASAP7_75t_L g742 ( .A(n_738), .B(n_733), .C(n_734), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_741), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_742), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_744), .A2(n_739), .B1(n_699), .B2(n_726), .Y(n_745) );
AO21x1_ASAP7_75t_L g746 ( .A1(n_745), .A2(n_743), .B(n_79), .Y(n_746) );
endmodule