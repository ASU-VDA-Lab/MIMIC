module fake_ariane_2126_n_30 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_30);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_30;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_27;
wire n_29;
wire n_17;
wire n_18;
wire n_28;
wire n_11;
wire n_26;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_1),
.Y(n_18)
);

NAND2x1p5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

OAI33xp33_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_14),
.A3(n_12),
.B1(n_11),
.B2(n_10),
.B3(n_15),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_19),
.B1(n_12),
.B2(n_17),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_13),
.C(n_3),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_13),
.B(n_3),
.C(n_4),
.Y(n_26)
);

OAI311xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.C1(n_6),
.Y(n_27)
);

NOR4xp25_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_13),
.C(n_23),
.D(n_6),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_27),
.B(n_28),
.Y(n_30)
);


endmodule