module fake_jpeg_379_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_52),
.C(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_75),
.B1(n_1),
.B2(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_48),
.B1(n_41),
.B2(n_39),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_80),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_48),
.B1(n_41),
.B2(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_78),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_57),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_6),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_19),
.C(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_10),
.B1(n_15),
.B2(n_24),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_107),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_7),
.B(n_8),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_106),
.B1(n_100),
.B2(n_113),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_27),
.B(n_32),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_25),
.A3(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_111),
.Y(n_117)
);

XOR2x1_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_37),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_87),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_30),
.B1(n_31),
.B2(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_94),
.B1(n_84),
.B2(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_111),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_102),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_121),
.B(n_110),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_128),
.B1(n_127),
.B2(n_121),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_126),
.B(n_120),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_117),
.Y(n_134)
);

INVxp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_109),
.C(n_124),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_136),
.Y(n_137)
);


endmodule