module fake_jpeg_27323_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_33),
.Y(n_49)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_55),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_19),
.Y(n_70)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_23),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_39),
.B1(n_45),
.B2(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_55),
.B1(n_54),
.B2(n_47),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_51),
.B1(n_48),
.B2(n_56),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_43),
.Y(n_86)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_27),
.B(n_26),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_29),
.B(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_46),
.B1(n_15),
.B2(n_23),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_47),
.B1(n_21),
.B2(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_26),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_72),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_67),
.C(n_66),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_105),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_103),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_72),
.B1(n_69),
.B2(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_102),
.B1(n_80),
.B2(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_73),
.B(n_20),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_20),
.C(n_22),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_72),
.Y(n_101)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_57),
.B1(n_64),
.B2(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_118),
.C(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_111),
.B1(n_102),
.B2(n_92),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_18),
.A3(n_17),
.B1(n_24),
.B2(n_29),
.C(n_5),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_95),
.B1(n_57),
.B2(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_129),
.B1(n_119),
.B2(n_118),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_96),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_132),
.Y(n_142)
);

OAI322xp33_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_97),
.A3(n_99),
.B1(n_18),
.B2(n_17),
.C1(n_11),
.C2(n_10),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_8),
.C(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_8),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_109),
.B1(n_107),
.B2(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_117),
.C(n_43),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_144),
.C(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_37),
.C(n_53),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_37),
.C(n_53),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_124),
.B(n_128),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_151),
.B(n_156),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_123),
.B(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_157),
.B1(n_0),
.B2(n_1),
.Y(n_161)
);

FAx1_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_133),
.CI(n_18),
.CON(n_156),
.SN(n_156)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_17),
.B(n_1),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_143),
.C(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_151),
.B(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_17),
.C(n_42),
.Y(n_164)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.C(n_165),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_156),
.B(n_153),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_170),
.Y(n_172)
);

AOI21x1_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_0),
.B(n_3),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_158),
.B(n_6),
.C(n_7),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_173),
.B(n_174),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_4),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_172),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_4),
.B(n_6),
.Y(n_178)
);


endmodule