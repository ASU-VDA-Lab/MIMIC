module fake_jpeg_11683_n_221 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_221);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_55),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_61),
.Y(n_67)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_18),
.B1(n_28),
.B2(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_31),
.B1(n_34),
.B2(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_37),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_86),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_115),
.B1(n_125),
.B2(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_99),
.Y(n_136)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_103),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_71),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_46),
.B1(n_40),
.B2(n_52),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_53),
.B1(n_54),
.B2(n_19),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_93),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_25),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_25),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_121),
.B(n_127),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_25),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_95),
.C(n_96),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_10),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_11),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_10),
.B1(n_11),
.B2(n_83),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_80),
.B1(n_74),
.B2(n_96),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_11),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_75),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_144),
.C(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_106),
.B1(n_107),
.B2(n_120),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_71),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_71),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_162),
.C(n_165),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_160),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_102),
.Y(n_160)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_119),
.B1(n_127),
.B2(n_109),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_163),
.B(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_147),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_101),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_119),
.B(n_121),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_134),
.B(n_138),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_118),
.CON(n_168),
.SN(n_168)
);

AOI322xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_131),
.A3(n_146),
.B1(n_128),
.B2(n_118),
.C1(n_150),
.C2(n_113),
.Y(n_174)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_178),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_167),
.A2(n_134),
.B(n_136),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_183),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_141),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_123),
.B(n_103),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_129),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_154),
.C(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_155),
.C(n_157),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_169),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_169),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_164),
.B1(n_156),
.B2(n_112),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_184),
.B1(n_180),
.B2(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_129),
.C(n_116),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_182),
.B1(n_183),
.B2(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_184),
.B1(n_178),
.B2(n_182),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_198),
.B(n_190),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_191),
.CI(n_198),
.CON(n_210),
.SN(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_212),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_203),
.C(n_201),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_211),
.A3(n_209),
.B1(n_210),
.B2(n_213),
.C1(n_149),
.C2(n_80),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_210),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_218),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_219),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_217),
.C(n_89),
.Y(n_221)
);


endmodule