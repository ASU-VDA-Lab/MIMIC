module fake_jpeg_26478_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_68),
.Y(n_92)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_20),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_81),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_26),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_89),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_35),
.B1(n_48),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_51),
.B1(n_61),
.B2(n_60),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_85),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_32),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_96),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_49),
.C(n_45),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_61),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_126),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_35),
.B1(n_50),
.B2(n_57),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_108),
.B1(n_109),
.B2(n_129),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_57),
.B1(n_50),
.B2(n_66),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_50),
.B1(n_57),
.B2(n_62),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_91),
.B(n_43),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_125),
.B1(n_90),
.B2(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_122),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_123)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_62),
.B1(n_55),
.B2(n_25),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_23),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_55),
.B1(n_25),
.B2(n_28),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_146),
.B1(n_142),
.B2(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_154),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_25),
.C(n_30),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_149),
.C(n_65),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_142),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_90),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_29),
.B(n_22),
.C(n_34),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_144),
.B(n_132),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_29),
.B(n_22),
.C(n_34),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_99),
.A3(n_95),
.B1(n_87),
.B2(n_70),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_42),
.C(n_43),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_86),
.B1(n_83),
.B2(n_81),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_71),
.B1(n_128),
.B2(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_155),
.Y(n_188)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_127),
.B(n_100),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_125),
.B(n_116),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_161),
.B(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_179),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_154),
.B1(n_80),
.B2(n_120),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_117),
.C(n_102),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_114),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_114),
.B(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_176),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_115),
.B1(n_128),
.B2(n_104),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_173),
.B1(n_186),
.B2(n_176),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_126),
.B1(n_115),
.B2(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_174),
.B(n_30),
.Y(n_212)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_115),
.B(n_100),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_130),
.B1(n_149),
.B2(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_183),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_184),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_70),
.B1(n_120),
.B2(n_80),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_0),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_171),
.B1(n_167),
.B2(n_158),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_208),
.C(n_159),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_197),
.Y(n_236)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_198),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_196),
.A2(n_199),
.B(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_137),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2x1p5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_134),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_212),
.Y(n_242)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_143),
.B1(n_144),
.B2(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_205),
.B(n_207),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_45),
.C(n_42),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_217),
.B1(n_183),
.B2(n_160),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_104),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_25),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_181),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_166),
.B(n_30),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_28),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_28),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_161),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_219),
.B1(n_216),
.B2(n_217),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_235),
.C(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_233),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_238),
.B1(n_244),
.B2(n_178),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_165),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_185),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_239),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_196),
.B1(n_195),
.B2(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_166),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_173),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_174),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_201),
.B1(n_196),
.B2(n_200),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_264),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_219),
.B1(n_216),
.B2(n_199),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_203),
.C(n_211),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_256),
.C(n_261),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_211),
.C(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_204),
.C(n_206),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_204),
.C(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_238),
.C(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_193),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_239),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_193),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_245),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B1(n_233),
.B2(n_242),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_245),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_271),
.B1(n_283),
.B2(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_232),
.B1(n_221),
.B2(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_237),
.C(n_227),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_273),
.C(n_275),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_260),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_229),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_286),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_241),
.B1(n_230),
.B2(n_234),
.Y(n_283)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_222),
.B1(n_4),
.B2(n_5),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_261),
.B1(n_250),
.B2(n_248),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_224),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_289),
.B(n_274),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_251),
.B(n_249),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_267),
.B1(n_268),
.B2(n_228),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_256),
.C(n_266),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.C(n_278),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_266),
.C(n_252),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_265),
.B(n_264),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_302),
.B1(n_269),
.B2(n_272),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_10),
.C(n_16),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_306),
.Y(n_317)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_270),
.C(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_291),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_270),
.B1(n_276),
.B2(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_315),
.B1(n_296),
.B2(n_302),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_276),
.C(n_19),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_9),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_19),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_293),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_12),
.B(n_15),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_310),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_322),
.B(n_12),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_307),
.C(n_309),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_294),
.B(n_295),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_303),
.B(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_327),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_304),
.C(n_312),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_308),
.C(n_313),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_330),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_331),
.B(n_15),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_316),
.A2(n_16),
.B(n_13),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_320),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_332),
.A2(n_335),
.B(n_319),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_337),
.A3(n_333),
.B1(n_4),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_6),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.C(n_7),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_6),
.C(n_7),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);


endmodule