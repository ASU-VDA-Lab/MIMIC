module real_jpeg_23984_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_131)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_77),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_42),
.B(n_87),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_99),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_5),
.A2(n_102),
.B1(n_188),
.B2(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_5),
.A2(n_37),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_25),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_27),
.B1(n_37),
.B2(n_70),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_70),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_27),
.B1(n_37),
.B2(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_82),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_82),
.Y(n_180)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_27),
.B1(n_37),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_64),
.B1(n_71),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_94),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_13),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_27),
.B1(n_37),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_67),
.Y(n_128)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_19),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_100),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_20),
.A2(n_21),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_22),
.B(n_54),
.C(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_23),
.A2(n_38),
.B1(n_39),
.B2(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_23),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_71),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_25),
.A2(n_33),
.B(n_35),
.Y(n_96)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_27),
.A2(n_37),
.B1(n_57),
.B2(n_61),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_27),
.B(n_35),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_35),
.A2(n_59),
.B(n_89),
.C(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_35),
.B(n_90),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_35),
.B(n_196),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_37),
.A2(n_57),
.A3(n_59),
.B1(n_208),
.B2(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_40),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_40),
.A2(n_105),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_41),
.A2(n_42),
.B1(n_87),
.B2(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_41),
.B(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_45),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_45),
.A2(n_47),
.B(n_126),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_49),
.B(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_50),
.A2(n_102),
.B1(n_180),
.B2(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_63),
.B(n_65),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_63),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_55),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_55),
.A2(n_98),
.B1(n_99),
.B2(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_56),
.A2(n_120),
.B1(n_146),
.B2(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_59),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_58),
.B(n_61),
.Y(n_215)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_66),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_73),
.B1(n_77),
.B2(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_83),
.B(n_100),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.C(n_97),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_97),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_85),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_85),
.A2(n_163),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_85),
.A2(n_171),
.B1(n_172),
.B2(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_108),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_90),
.A2(n_130),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_90),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_91),
.B(n_171),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_107),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_102),
.A2(n_127),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_102),
.A2(n_104),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_111),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_124),
.CI(n_132),
.CON(n_111),
.SN(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_130),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_153),
.B(n_243),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_150),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_137),
.B(n_150),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_138),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_140),
.A2(n_142),
.B1(n_143),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_148),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_144),
.B(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_147),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_237),
.B(n_242),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_221),
.B(n_236),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_201),
.B(n_220),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_176),
.B(n_200),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_158),
.B(n_166),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_173),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_173),
.C(n_174),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_184),
.B(n_199),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_182),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_198),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_212),
.C(n_218),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_231),
.C(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule