module fake_jpeg_30216_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_69),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_91),
.Y(n_160)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_19),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_79),
.Y(n_134)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_13),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_34),
.B(n_13),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_11),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_33),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_125),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_26),
.B(n_20),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g170 ( 
.A(n_119),
.B(n_30),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_122),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_53),
.B(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_28),
.B1(n_42),
.B2(n_38),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_131),
.A2(n_70),
.B1(n_71),
.B2(n_81),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_145),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_79),
.A2(n_19),
.B1(n_37),
.B2(n_32),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_141),
.A2(n_30),
.B1(n_84),
.B2(n_78),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_55),
.B(n_33),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx4f_ASAP7_75t_SL g148 ( 
.A(n_61),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_59),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_157),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_52),
.B(n_48),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_85),
.B(n_22),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_77),
.B(n_22),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_167),
.B(n_191),
.Y(n_259)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g251 ( 
.A(n_170),
.B(n_187),
.Y(n_251)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_65),
.C(n_75),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_172),
.B(n_196),
.C(n_112),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_173),
.B(n_202),
.Y(n_246)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_101),
.B1(n_59),
.B2(n_82),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_182),
.A2(n_118),
.B1(n_166),
.B2(n_155),
.Y(n_255)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_36),
.B(n_26),
.C(n_30),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_36),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_136),
.B(n_116),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_132),
.A2(n_102),
.B1(n_99),
.B2(n_95),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_212),
.B1(n_213),
.B2(n_223),
.Y(n_237)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_107),
.B(n_45),
.Y(n_202)
);

CKINVDCx12_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_110),
.B(n_113),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_208),
.A2(n_209),
.B1(n_227),
.B2(n_42),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_110),
.A2(n_28),
.B1(n_38),
.B2(n_21),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_163),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_215),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_144),
.Y(n_211)
);

BUFx4f_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_93),
.B1(n_76),
.B2(n_46),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_118),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_113),
.B(n_28),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_219),
.Y(n_273)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_143),
.A2(n_30),
.B(n_11),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_218),
.B(n_0),
.Y(n_257)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_143),
.B(n_21),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_105),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_222),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_127),
.A2(n_46),
.B1(n_29),
.B2(n_37),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_226),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_141),
.A2(n_38),
.B1(n_21),
.B2(n_42),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_139),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_245),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_142),
.B1(n_156),
.B2(n_137),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_243),
.A2(n_153),
.B1(n_82),
.B2(n_221),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_174),
.B(n_162),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_196),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_263),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_176),
.B(n_45),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_266),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_272),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_172),
.B(n_161),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_196),
.B(n_152),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_185),
.B(n_45),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_170),
.B(n_46),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_179),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_269),
.B(n_1),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_121),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_154),
.C(n_115),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_228),
.C(n_188),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_190),
.B1(n_214),
.B2(n_200),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_278),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_229),
.B1(n_251),
.B2(n_245),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_283),
.B(n_292),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_237),
.A2(n_224),
.B1(n_213),
.B2(n_204),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_284),
.A2(n_287),
.B1(n_297),
.B2(n_315),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_246),
.B(n_188),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_285),
.B(n_286),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_237),
.A2(n_194),
.B1(n_199),
.B2(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_251),
.A2(n_228),
.B(n_182),
.C(n_148),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_291),
.A2(n_271),
.B(n_242),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_177),
.C(n_180),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_282),
.C(n_280),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_184),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_295),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_225),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_296),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_178),
.B1(n_37),
.B2(n_32),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_300),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_45),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_301),
.A2(n_318),
.B1(n_323),
.B2(n_317),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_232),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_45),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_311),
.Y(n_351)
);

AOI22x1_ASAP7_75t_SL g305 ( 
.A1(n_234),
.A2(n_168),
.B1(n_153),
.B2(n_180),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_305),
.A2(n_326),
.B(n_234),
.Y(n_328)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_306),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_234),
.B1(n_240),
.B2(n_275),
.Y(n_327)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_0),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_232),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_312),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_168),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_214),
.B1(n_200),
.B2(n_217),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_181),
.B(n_31),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_316),
.A2(n_233),
.B(n_265),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_277),
.A2(n_159),
.B1(n_31),
.B2(n_3),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_231),
.Y(n_321)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_322),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_323)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_324),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_1),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_233),
.Y(n_352)
);

INVx13_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

INVx13_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_329),
.A2(n_367),
.B(n_294),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_342),
.C(n_344),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_281),
.A2(n_254),
.B(n_266),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_340),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_284),
.B1(n_286),
.B2(n_288),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_352),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_308),
.A2(n_245),
.B(n_229),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_257),
.C(n_238),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_L g348 ( 
.A1(n_298),
.A2(n_236),
.B(n_264),
.Y(n_348)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_SL g354 ( 
.A(n_299),
.B(n_260),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_320),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_265),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_363),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_239),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_283),
.C(n_299),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_305),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_317),
.A2(n_267),
.B1(n_258),
.B2(n_231),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_290),
.B(n_261),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_364),
.B(n_300),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_297),
.B1(n_325),
.B2(n_316),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_271),
.B(n_242),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_292),
.Y(n_374)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_400),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_335),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_346),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_379),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_361),
.B(n_311),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_384),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_386),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

INVx13_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_329),
.A2(n_291),
.B1(n_318),
.B2(n_315),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_357),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_389),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_351),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_391),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_304),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_309),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_392),
.B(n_396),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_366),
.A2(n_294),
.B1(n_299),
.B2(n_321),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_393),
.A2(n_398),
.B1(n_343),
.B2(n_334),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_350),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_401),
.B(n_367),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_337),
.B(n_351),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_334),
.A2(n_310),
.B1(n_303),
.B2(n_307),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_365),
.B(n_289),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_350),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_360),
.A2(n_319),
.B(n_314),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_360),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_SL g439 ( 
.A(n_403),
.B(n_386),
.C(n_387),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_360),
.B(n_362),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_410),
.A2(n_402),
.B(n_363),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_412),
.A2(n_416),
.B(n_383),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_397),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_414),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_395),
.A2(n_340),
.B(n_365),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_417),
.B(n_369),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_427),
.Y(n_435)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_359),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_430),
.Y(n_434)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_425),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_344),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_372),
.A2(n_343),
.B1(n_342),
.B2(n_354),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_381),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_404),
.A2(n_372),
.B1(n_386),
.B2(n_390),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_448),
.B1(n_427),
.B2(n_418),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_438),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_406),
.B(n_400),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_454),
.B(n_455),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_408),
.A2(n_393),
.B1(n_398),
.B2(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_379),
.Y(n_441)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_368),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_449),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_426),
.B(n_409),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_452),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_404),
.A2(n_380),
.B1(n_382),
.B2(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_411),
.A2(n_373),
.B1(n_382),
.B2(n_401),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_378),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_391),
.Y(n_450)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_374),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_456),
.C(n_459),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_364),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_389),
.C(n_388),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_474),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_439),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_463),
.B(n_469),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_475),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_481),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_412),
.C(n_416),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_445),
.B(n_411),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_470),
.Y(n_489)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_415),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_415),
.C(n_418),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_480),
.Y(n_485)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_394),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_418),
.C(n_410),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_451),
.C(n_442),
.Y(n_481)
);

OAI31xp33_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_455),
.A3(n_436),
.B(n_454),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_487),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_468),
.A2(n_403),
.B(n_448),
.Y(n_487)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_407),
.B1(n_405),
.B2(n_432),
.Y(n_490)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_424),
.B1(n_447),
.B2(n_376),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_492),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_464),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_475),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_494),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_413),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_456),
.B(n_449),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_495),
.A2(n_480),
.B(n_477),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_402),
.B(n_375),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_496),
.B(n_402),
.Y(n_510)
);

AO221x1_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_353),
.B1(n_420),
.B2(n_414),
.C(n_385),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_478),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_489),
.A2(n_461),
.B1(n_469),
.B2(n_462),
.Y(n_499)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_488),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_502),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_510),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_483),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_481),
.C(n_466),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_507),
.B(n_509),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_489),
.B(n_466),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_472),
.C(n_460),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_485),
.C(n_495),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_512),
.A2(n_492),
.B1(n_487),
.B2(n_493),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_514),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_485),
.C(n_484),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_520),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_498),
.C(n_472),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_498),
.C(n_494),
.Y(n_528)
);

XOR2x1_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_486),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_496),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_516),
.A2(n_518),
.B(n_514),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_523),
.B(n_525),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_519),
.A2(n_503),
.B1(n_501),
.B2(n_500),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_506),
.B(n_505),
.Y(n_526)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_526),
.A2(n_521),
.A3(n_515),
.B1(n_336),
.B2(n_338),
.C1(n_326),
.C2(n_324),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_529),
.A3(n_336),
.B1(n_338),
.B2(n_306),
.C1(n_460),
.C2(n_438),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_521),
.B1(n_420),
.B2(n_413),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_530),
.A2(n_528),
.B1(n_527),
.B2(n_524),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_533),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_532),
.B1(n_261),
.B2(n_256),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_536),
.A2(n_537),
.B(n_535),
.Y(n_538)
);

AOI322xp5_ASAP7_75t_L g537 ( 
.A1(n_534),
.A2(n_256),
.A3(n_247),
.B1(n_241),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_537)
);

AOI322xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_247),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_539)
);

AO221x1_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_7),
.C(n_8),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_9),
.C(n_10),
.Y(n_542)
);


endmodule