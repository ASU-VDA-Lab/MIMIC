module fake_ibex_1559_n_2703 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_482, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2703);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2703;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_2230;
wire n_1782;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_2176;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2263;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2669;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_2433;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1385;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_704;
wire n_2357;
wire n_2104;
wire n_2618;
wire n_2653;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2453;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g496 ( 
.A(n_418),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_43),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_56),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_358),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_140),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_114),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_193),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_379),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_296),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_99),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_237),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_223),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_315),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_97),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_35),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_234),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_261),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_265),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_226),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_298),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_443),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_285),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_248),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_280),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_316),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_140),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_178),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_19),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_19),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_455),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_99),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_409),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_153),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_350),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_202),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_43),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_313),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_484),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_145),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_459),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_413),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_111),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_339),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_70),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_71),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_161),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_289),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_159),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_367),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_402),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_204),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_363),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_197),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_251),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_184),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_401),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_122),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_211),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_35),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_411),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_36),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_295),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_150),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_365),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_147),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_477),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_377),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_467),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_303),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_219),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_63),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_174),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_52),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_420),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_371),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_188),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_299),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_142),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_148),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_432),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_352),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_329),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_3),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_36),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_230),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_272),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_267),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_240),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_155),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_376),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_364),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_186),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_74),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_300),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_132),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_90),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_160),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_143),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_121),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_453),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_270),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_341),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_209),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_146),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_215),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_190),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_58),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_274),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_8),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_220),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_104),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_104),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_254),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_198),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_210),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_347),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_419),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_86),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_325),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_205),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_129),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_206),
.Y(n_621)
);

BUFx8_ASAP7_75t_SL g622 ( 
.A(n_12),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_157),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_429),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_9),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_410),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_149),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_102),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_85),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_318),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_67),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_45),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_472),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_218),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_264),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_286),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_408),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_112),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_336),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_475),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_331),
.Y(n_641)
);

CKINVDCx14_ASAP7_75t_R g642 ( 
.A(n_126),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_427),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_129),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_74),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_241),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_242),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_111),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_422),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_245),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_6),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_1),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_123),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_155),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_214),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_108),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_257),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_482),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_330),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_76),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_259),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_271),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_378),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_133),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_192),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_142),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_164),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_118),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_87),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_333),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_124),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_292),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_273),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_22),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_47),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_115),
.Y(n_676)
);

CKINVDCx14_ASAP7_75t_R g677 ( 
.A(n_182),
.Y(n_677)
);

BUFx8_ASAP7_75t_SL g678 ( 
.A(n_243),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_229),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_460),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_462),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_384),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_394),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_119),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_461),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_20),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_400),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_175),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_278),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_433),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_312),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_451),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_101),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_110),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_95),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_253),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_79),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_372),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_290),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_49),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_486),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_407),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_133),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_82),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_233),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_145),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_32),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_470),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_366),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_11),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_362),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_353),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_335),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_480),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_162),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_398),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_212),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_423),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_391),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_93),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_165),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_392),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_416),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_326),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_2),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_28),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_332),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_176),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_115),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_144),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_415),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_277),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_93),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_247),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_493),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_199),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_66),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_321),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_108),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_27),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_385),
.Y(n_741)
);

BUFx8_ASAP7_75t_SL g742 ( 
.A(n_45),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_67),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_386),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_51),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_73),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_236),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_291),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_343),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_12),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_88),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_334),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_436),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_469),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_293),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_130),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_360),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_301),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_121),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_27),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_239),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_275),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_40),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_22),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_88),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_232),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_113),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_110),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_345),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_490),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_124),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_268),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_485),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_344),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_123),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_96),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_76),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_464),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_150),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_180),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_61),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_34),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_11),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_314),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_39),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_20),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_97),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_167),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_355),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_308),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_483),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_387),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_458),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_369),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_389),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_0),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_488),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_317),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_302),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_109),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_23),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_135),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_255),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_474),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_258),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_307),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_395),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_166),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_425),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_441),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_15),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_128),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_262),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_130),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_147),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_381),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_119),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_3),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_228),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_473),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_139),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_494),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_309),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_456),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_297),
.Y(n_825)
);

BUFx12f_ASAP7_75t_L g826 ( 
.A(n_777),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_678),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_616),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_616),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_499),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_559),
.B(n_0),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_804),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_800),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_770),
.B(n_1),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_805),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_800),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_559),
.B(n_2),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_664),
.Y(n_839)
);

BUFx8_ASAP7_75t_SL g840 ( 
.A(n_622),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_616),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_664),
.B(n_4),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_695),
.B(n_4),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_616),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_698),
.Y(n_845)
);

INVx5_ASAP7_75t_L g846 ( 
.A(n_499),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_695),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_775),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_777),
.Y(n_849)
);

INVx5_ASAP7_75t_L g850 ( 
.A(n_499),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_698),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_775),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_581),
.B(n_5),
.Y(n_853)
);

BUFx8_ASAP7_75t_SL g854 ( 
.A(n_742),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_497),
.B(n_5),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_681),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_777),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_516),
.B(n_6),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_783),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_783),
.B(n_7),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_516),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_681),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_563),
.B(n_7),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_681),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_642),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_698),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_576),
.B(n_8),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_576),
.B(n_9),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_563),
.B(n_10),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_10),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_644),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_524),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_731),
.B(n_13),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_666),
.B(n_13),
.Y(n_874)
);

BUFx8_ASAP7_75t_SL g875 ( 
.A(n_591),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_666),
.B(n_14),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_523),
.B(n_492),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_555),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_644),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_731),
.B(n_14),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_769),
.B(n_15),
.Y(n_881)
);

AND2x6_ASAP7_75t_L g882 ( 
.A(n_512),
.B(n_156),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_644),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_629),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_512),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_769),
.B(n_16),
.Y(n_886)
);

BUFx12f_ASAP7_75t_L g887 ( 
.A(n_524),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_656),
.B(n_16),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_644),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_569),
.B(n_502),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_698),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_568),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_527),
.B(n_17),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_502),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_812),
.B(n_17),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_568),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_538),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_599),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_599),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_540),
.B(n_18),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_624),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_574),
.B(n_18),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_525),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_547),
.B(n_21),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_547),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_609),
.B(n_636),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_587),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_597),
.B(n_21),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_625),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_624),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_638),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_673),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_609),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_525),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_529),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_508),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_645),
.Y(n_917)
);

BUFx8_ASAP7_75t_SL g918 ( 
.A(n_591),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_652),
.B(n_23),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_654),
.B(n_24),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_660),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_673),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_674),
.B(n_24),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_809),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_636),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_675),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_720),
.B(n_25),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_730),
.B(n_25),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_662),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_809),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_739),
.B(n_743),
.Y(n_931)
);

BUFx8_ASAP7_75t_L g932 ( 
.A(n_496),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_662),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_778),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_529),
.B(n_26),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_745),
.B(n_26),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_532),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_746),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_778),
.B(n_28),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_29),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_807),
.B(n_29),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_807),
.Y(n_942)
);

AND2x6_ASAP7_75t_L g943 ( 
.A(n_506),
.B(n_489),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_523),
.B(n_158),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_507),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_764),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_677),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_820),
.Y(n_948)
);

BUFx8_ASAP7_75t_SL g949 ( 
.A(n_631),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_518),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_631),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_532),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_535),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_503),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_826),
.B(n_776),
.Y(n_955)
);

OAI22xp33_ASAP7_75t_R g956 ( 
.A1(n_884),
.A2(n_668),
.B1(n_763),
.B2(n_617),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_878),
.A2(n_541),
.B1(n_802),
.B2(n_535),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_878),
.A2(n_802),
.B1(n_541),
.B2(n_519),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_865),
.B(n_526),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_832),
.Y(n_960)
);

OAI22xp33_ASAP7_75t_L g961 ( 
.A1(n_951),
.A2(n_693),
.B1(n_725),
.B2(n_648),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_903),
.A2(n_500),
.B1(n_501),
.B2(n_498),
.Y(n_962)
);

OAI22xp33_ASAP7_75t_L g963 ( 
.A1(n_903),
.A2(n_693),
.B1(n_725),
.B2(n_648),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_832),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_857),
.B(n_831),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_896),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_865),
.B(n_526),
.Y(n_967)
);

OAI22xp33_ASAP7_75t_L g968 ( 
.A1(n_915),
.A2(n_767),
.B1(n_815),
.B2(n_737),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_953),
.B(n_528),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_896),
.Y(n_970)
);

OAI22xp33_ASAP7_75t_SL g971 ( 
.A1(n_915),
.A2(n_505),
.B1(n_510),
.B2(n_509),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_838),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_831),
.B(n_781),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_828),
.A2(n_508),
.B1(n_536),
.B2(n_519),
.Y(n_974)
);

AND2x2_ASAP7_75t_SL g975 ( 
.A(n_867),
.B(n_785),
.Y(n_975)
);

AOI22x1_ASAP7_75t_L g976 ( 
.A1(n_834),
.A2(n_533),
.B1(n_539),
.B2(n_521),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_840),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_SL g978 ( 
.A1(n_842),
.A2(n_553),
.B1(n_557),
.B2(n_522),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_833),
.A2(n_579),
.B1(n_588),
.B2(n_536),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_896),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_838),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_853),
.A2(n_588),
.B1(n_657),
.B2(n_579),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_898),
.Y(n_983)
);

CKINVDCx6p67_ASAP7_75t_R g984 ( 
.A(n_872),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_898),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_857),
.B(n_528),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_867),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_888),
.A2(n_688),
.B1(n_723),
.B2(n_657),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_887),
.A2(n_767),
.B1(n_815),
.B2(n_737),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_856),
.B(n_530),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_831),
.B(n_530),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_914),
.B(n_786),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_868),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_937),
.A2(n_723),
.B1(n_744),
.B2(n_688),
.Y(n_994)
);

AO22x2_ASAP7_75t_L g995 ( 
.A1(n_855),
.A2(n_796),
.B1(n_801),
.B2(n_787),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_952),
.B(n_817),
.Y(n_996)
);

OAI22xp33_ASAP7_75t_L g997 ( 
.A1(n_836),
.A2(n_755),
.B1(n_757),
.B2(n_744),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_831),
.B(n_531),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_846),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_868),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_849),
.A2(n_757),
.B1(n_798),
.B2(n_755),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_846),
.B(n_545),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_898),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_874),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_846),
.B(n_821),
.Y(n_1005)
);

AO22x2_ASAP7_75t_L g1006 ( 
.A1(n_870),
.A2(n_551),
.B1(n_562),
.B2(n_552),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_893),
.A2(n_575),
.B1(n_582),
.B2(n_571),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_846),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_874),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_935),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_876),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_850),
.B(n_531),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_895),
.A2(n_798),
.B1(n_567),
.B2(n_580),
.Y(n_1013)
);

OAI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_902),
.A2(n_593),
.B1(n_594),
.B2(n_561),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_893),
.A2(n_603),
.B1(n_606),
.B2(n_596),
.Y(n_1015)
);

AO22x2_ASAP7_75t_L g1016 ( 
.A1(n_900),
.A2(n_908),
.B1(n_928),
.B2(n_923),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_900),
.A2(n_610),
.B1(n_611),
.B2(n_608),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_850),
.B(n_534),
.Y(n_1018)
);

OA22x2_ASAP7_75t_L g1019 ( 
.A1(n_827),
.A2(n_627),
.B1(n_628),
.B2(n_620),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_922),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_876),
.Y(n_1021)
);

AO22x2_ASAP7_75t_L g1022 ( 
.A1(n_908),
.A2(n_584),
.B1(n_585),
.B2(n_583),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_916),
.Y(n_1023)
);

AO22x2_ASAP7_75t_L g1024 ( 
.A1(n_923),
.A2(n_590),
.B1(n_598),
.B2(n_589),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_850),
.B(n_534),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_922),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_928),
.A2(n_651),
.B1(n_653),
.B2(n_632),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_SL g1028 ( 
.A1(n_875),
.A2(n_671),
.B1(n_676),
.B2(n_669),
.Y(n_1028)
);

OAI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_902),
.A2(n_920),
.B1(n_927),
.B2(n_919),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_875),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_922),
.Y(n_1031)
);

OAI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_919),
.A2(n_686),
.B1(n_694),
.B2(n_684),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_924),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_850),
.B(n_537),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_842),
.A2(n_700),
.B1(n_703),
.B2(n_697),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_924),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_862),
.B(n_537),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_SL g1038 ( 
.A1(n_918),
.A2(n_949),
.B1(n_704),
.B2(n_707),
.Y(n_1038)
);

OAI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_920),
.A2(n_706),
.B1(n_726),
.B2(n_710),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_909),
.B(n_729),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_885),
.Y(n_1041)
);

OAI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_927),
.A2(n_733),
.B1(n_750),
.B2(n_740),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_862),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_835),
.A2(n_751),
.B1(n_760),
.B2(n_759),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_938),
.B(n_765),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_862),
.B(n_542),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_950),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_918),
.A2(n_768),
.B1(n_779),
.B2(n_771),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_873),
.B(n_880),
.Y(n_1049)
);

INVx8_ASAP7_75t_L g1050 ( 
.A(n_862),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_864),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_835),
.A2(n_782),
.B1(n_814),
.B2(n_811),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_890),
.A2(n_795),
.B1(n_797),
.B2(n_542),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_890),
.A2(n_797),
.B1(n_799),
.B2(n_795),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_931),
.A2(n_602),
.B1(n_612),
.B2(n_601),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_864),
.B(n_799),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_924),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_931),
.A2(n_803),
.B1(n_634),
.B2(n_635),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_864),
.B(n_803),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_864),
.B(n_504),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_SL g1061 ( 
.A1(n_946),
.A2(n_637),
.B1(n_643),
.B2(n_613),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_858),
.A2(n_649),
.B1(n_661),
.B2(n_646),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_847),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_840),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_936),
.A2(n_692),
.B1(n_699),
.B2(n_691),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_848),
.B(n_511),
.Y(n_1066)
);

OA22x2_ASAP7_75t_L g1067 ( 
.A1(n_907),
.A2(n_709),
.B1(n_715),
.B2(n_708),
.Y(n_1067)
);

OAI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_936),
.A2(n_718),
.B1(n_719),
.B2(n_716),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_897),
.A2(n_732),
.B1(n_734),
.B2(n_724),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_839),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_852),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_859),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_854),
.Y(n_1073)
);

AO22x2_ASAP7_75t_L g1074 ( 
.A1(n_843),
.A2(n_860),
.B1(n_880),
.B2(n_873),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_843),
.A2(n_738),
.B1(n_741),
.B2(n_736),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_897),
.B(n_911),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_945),
.B(n_748),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_858),
.A2(n_761),
.B1(n_766),
.B2(n_758),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_860),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_861),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_911),
.B(n_513),
.Y(n_1081)
);

AO22x2_ASAP7_75t_L g1082 ( 
.A1(n_881),
.A2(n_792),
.B1(n_793),
.B2(n_780),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_917),
.B(n_514),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_947),
.B(n_794),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_881),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_837),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_899),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_917),
.B(n_921),
.Y(n_1088)
);

OAI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_877),
.A2(n_813),
.B1(n_822),
.B2(n_808),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_863),
.Y(n_1090)
);

AO22x2_ASAP7_75t_L g1091 ( 
.A1(n_940),
.A2(n_570),
.B1(n_825),
.B2(n_543),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_921),
.B(n_515),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_930),
.Y(n_1093)
);

AO22x2_ASAP7_75t_L g1094 ( 
.A1(n_940),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_863),
.A2(n_520),
.B1(n_544),
.B2(n_517),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_950),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_926),
.B(n_30),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_869),
.A2(n_548),
.B1(n_549),
.B2(n_546),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_926),
.B(n_550),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_854),
.B(n_31),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_894),
.B(n_33),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_869),
.A2(n_886),
.B1(n_939),
.B2(n_904),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_886),
.A2(n_824),
.B1(n_556),
.B2(n_558),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_950),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_934),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_904),
.A2(n_560),
.B1(n_564),
.B2(n_554),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_934),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_877),
.A2(n_566),
.B1(n_572),
.B2(n_565),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_939),
.A2(n_577),
.B1(n_578),
.B2(n_573),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_905),
.A2(n_37),
.B1(n_33),
.B2(n_34),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_947),
.B(n_586),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_947),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_947),
.B(n_592),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_944),
.A2(n_600),
.B1(n_604),
.B2(n_595),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_948),
.B(n_605),
.Y(n_1115)
);

OAI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_944),
.A2(n_614),
.B1(n_615),
.B2(n_607),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_934),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_948),
.B(n_618),
.Y(n_1118)
);

OA22x2_ASAP7_75t_L g1119 ( 
.A1(n_913),
.A2(n_621),
.B1(n_623),
.B2(n_619),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_925),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_929),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_941),
.A2(n_630),
.B1(n_633),
.B2(n_626),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_933),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_R g1124 ( 
.A1(n_941),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1124)
);

AOI22x1_ASAP7_75t_SL g1125 ( 
.A1(n_932),
.A2(n_640),
.B1(n_641),
.B2(n_639),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_932),
.A2(n_650),
.B1(n_655),
.B2(n_647),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_861),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_942),
.B(n_658),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_SL g1129 ( 
.A1(n_906),
.A2(n_663),
.B1(n_665),
.B2(n_659),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_948),
.B(n_667),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_948),
.B(n_670),
.Y(n_1131)
);

OAI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_906),
.A2(n_679),
.B1(n_680),
.B2(n_672),
.Y(n_1132)
);

AND2x2_ASAP7_75t_SL g1133 ( 
.A(n_882),
.B(n_682),
.Y(n_1133)
);

AO22x2_ASAP7_75t_L g1134 ( 
.A1(n_871),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_892),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_879),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_892),
.A2(n_910),
.B1(n_912),
.B2(n_901),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_954),
.B(n_683),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_892),
.Y(n_1139)
);

AO22x2_ASAP7_75t_L g1140 ( 
.A1(n_883),
.A2(n_889),
.B1(n_943),
.B2(n_882),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_892),
.A2(n_687),
.B1(n_689),
.B2(n_685),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_943),
.A2(n_823),
.B1(n_696),
.B2(n_701),
.Y(n_1142)
);

AO22x2_ASAP7_75t_L g1143 ( 
.A1(n_943),
.A2(n_44),
.B1(n_41),
.B2(n_42),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_901),
.B(n_690),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_943),
.A2(n_882),
.B1(n_705),
.B2(n_711),
.Y(n_1145)
);

OAI22xp33_ASAP7_75t_R g1146 ( 
.A1(n_901),
.A2(n_46),
.B1(n_42),
.B2(n_44),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_901),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_910),
.B(n_702),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_882),
.A2(n_819),
.B1(n_713),
.B2(n_714),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_910),
.B(n_712),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_910),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_912),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_SL g1153 ( 
.A1(n_912),
.A2(n_816),
.B1(n_721),
.B2(n_722),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_954),
.A2(n_727),
.B1(n_728),
.B2(n_717),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_912),
.B(n_46),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_SL g1156 ( 
.A1(n_954),
.A2(n_747),
.B1(n_749),
.B2(n_735),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_954),
.A2(n_810),
.B1(n_753),
.B2(n_754),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_829),
.A2(n_762),
.B1(n_773),
.B2(n_752),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_829),
.Y(n_1159)
);

AO22x2_ASAP7_75t_L g1160 ( 
.A1(n_829),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_830),
.B(n_774),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_891),
.B(n_784),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_830),
.A2(n_789),
.B1(n_790),
.B2(n_788),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_841),
.A2(n_806),
.B1(n_791),
.B2(n_51),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_841),
.A2(n_52),
.B1(n_48),
.B2(n_50),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_841),
.A2(n_54),
.B1(n_50),
.B2(n_53),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_844),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_844),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1085),
.A2(n_851),
.B(n_845),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1079),
.B(n_845),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1120),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1121),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1029),
.A2(n_851),
.B(n_845),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1076),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_1001),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_1145),
.B(n_851),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1010),
.B(n_55),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1088),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1070),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1071),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1072),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1063),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1097),
.Y(n_1183)
);

XNOR2xp5_ASAP7_75t_L g1184 ( 
.A(n_982),
.B(n_56),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1010),
.B(n_57),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_964),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1074),
.B(n_866),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1040),
.B(n_163),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1047),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_964),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_987),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1049),
.A2(n_1074),
.B(n_1140),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_987),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_969),
.B(n_57),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_959),
.B(n_58),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_988),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1004),
.Y(n_1197)
);

XNOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_974),
.B(n_59),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1004),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1023),
.B(n_963),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_958),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1101),
.Y(n_1202)
);

AND2x2_ASAP7_75t_SL g1203 ( 
.A(n_979),
.B(n_59),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1047),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1102),
.B(n_866),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_960),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1096),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_986),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_984),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_972),
.Y(n_1210)
);

XOR2x2_ASAP7_75t_L g1211 ( 
.A(n_1038),
.B(n_60),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1080),
.B(n_60),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_981),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1016),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1081),
.B(n_866),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_967),
.B(n_61),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1127),
.B(n_62),
.Y(n_1217)
);

INVxp33_ASAP7_75t_L g1218 ( 
.A(n_1028),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1016),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1048),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1123),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1123),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1086),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_957),
.B(n_62),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1096),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_990),
.B(n_63),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_965),
.B(n_1128),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1013),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_993),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1000),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1009),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1045),
.B(n_168),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1011),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1105),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1066),
.B(n_169),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_975),
.B(n_64),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1107),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1128),
.B(n_1083),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1021),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1117),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1133),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1092),
.B(n_891),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1082),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1082),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_955),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1069),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1149),
.B(n_891),
.Y(n_1247)
);

XOR2xp5_ASAP7_75t_L g1248 ( 
.A(n_961),
.B(n_64),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1087),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1093),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_966),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1067),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1099),
.B(n_965),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1160),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1005),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_970),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1005),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1155),
.Y(n_1258)
);

XOR2xp5_ASAP7_75t_L g1259 ( 
.A(n_994),
.B(n_65),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_995),
.B(n_65),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1143),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1007),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1007),
.Y(n_1263)
);

XNOR2x2_ASAP7_75t_L g1264 ( 
.A(n_1160),
.B(n_66),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1022),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1022),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1024),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1024),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_995),
.B(n_68),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1055),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1100),
.B(n_68),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1055),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_980),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1053),
.B(n_69),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1043),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1090),
.B(n_170),
.Y(n_1276)
);

INVxp33_ASAP7_75t_L g1277 ( 
.A(n_1054),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_983),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1140),
.A2(n_172),
.B(n_171),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1108),
.B(n_173),
.Y(n_1281)
);

XOR2xp5_ASAP7_75t_L g1282 ( 
.A(n_1125),
.B(n_69),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_985),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1110),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_955),
.B(n_70),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1090),
.B(n_177),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1006),
.B(n_71),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1110),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1041),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_973),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_R g1291 ( 
.A(n_977),
.B(n_72),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1151),
.A2(n_181),
.B(n_179),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1114),
.B(n_183),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1050),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1050),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_992),
.B(n_72),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_991),
.B(n_185),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1003),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1062),
.A2(n_487),
.B(n_189),
.Y(n_1299)
);

INVxp33_ASAP7_75t_L g1300 ( 
.A(n_1061),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1006),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_999),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1008),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_976),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1094),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_998),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_992),
.B(n_73),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1046),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_996),
.B(n_1044),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1094),
.Y(n_1310)
);

CKINVDCx14_ASAP7_75t_R g1311 ( 
.A(n_1064),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1095),
.B(n_187),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1134),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1020),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_968),
.B(n_75),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1030),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1026),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1018),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1034),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1134),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1098),
.B(n_191),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1103),
.B(n_194),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1037),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1058),
.B(n_195),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1056),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1106),
.B(n_1078),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1162),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1119),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1132),
.B(n_196),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_997),
.B(n_75),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1031),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1051),
.Y(n_1332)
);

XOR2x2_ASAP7_75t_L g1333 ( 
.A(n_1019),
.B(n_77),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1075),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1129),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1077),
.Y(n_1336)
);

INVx4_ASAP7_75t_SL g1337 ( 
.A(n_996),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1015),
.B(n_200),
.Y(n_1338)
);

XOR2xp5_ASAP7_75t_L g1339 ( 
.A(n_989),
.B(n_77),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1065),
.A2(n_203),
.B(n_201),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1002),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1104),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1012),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1025),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1091),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_R g1346 ( 
.A(n_1100),
.B(n_78),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1033),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1068),
.A2(n_208),
.B(n_207),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1142),
.A2(n_216),
.B(n_213),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1060),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1164),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1017),
.B(n_217),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1036),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1052),
.B(n_78),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1057),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1091),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1084),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1135),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1027),
.B(n_79),
.Y(n_1359)
);

INVxp33_ASAP7_75t_SL g1360 ( 
.A(n_1109),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1126),
.B(n_80),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1139),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1116),
.B(n_221),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1014),
.A2(n_224),
.B(n_222),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1147),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1154),
.B(n_80),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1059),
.B(n_225),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1152),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1032),
.B(n_227),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1165),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1113),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1136),
.Y(n_1372)
);

XNOR2x2_ASAP7_75t_L g1373 ( 
.A(n_956),
.B(n_81),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1166),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1168),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_978),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1035),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1144),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1157),
.B(n_81),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1148),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1150),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1115),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1073),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1118),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1130),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1089),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1158),
.B(n_1163),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1159),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1039),
.Y(n_1389)
);

XOR2xp5_ASAP7_75t_L g1390 ( 
.A(n_1122),
.B(n_82),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1042),
.B(n_231),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1112),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_962),
.Y(n_1393)
);

INVxp33_ASAP7_75t_L g1394 ( 
.A(n_956),
.Y(n_1394)
);

XNOR2xp5_ASAP7_75t_L g1395 ( 
.A(n_971),
.B(n_83),
.Y(n_1395)
);

XOR2xp5_ASAP7_75t_L g1396 ( 
.A(n_1156),
.B(n_83),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1131),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1141),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1153),
.B(n_1138),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1161),
.B(n_84),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1137),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1111),
.Y(n_1402)
);

XNOR2xp5_ASAP7_75t_L g1403 ( 
.A(n_1124),
.B(n_84),
.Y(n_1403)
);

XNOR2xp5_ASAP7_75t_L g1404 ( 
.A(n_1124),
.B(n_85),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1146),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1146),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1167),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1079),
.B(n_235),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1079),
.B(n_238),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1076),
.Y(n_1410)
);

XOR2xp5_ASAP7_75t_L g1411 ( 
.A(n_1001),
.B(n_86),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1080),
.B(n_87),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1076),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1080),
.B(n_89),
.Y(n_1414)
);

XNOR2x2_ASAP7_75t_L g1415 ( 
.A(n_1160),
.B(n_89),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1079),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1076),
.Y(n_1417)
);

XNOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1160),
.B(n_90),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1076),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_969),
.Y(n_1420)
);

XOR2x2_ASAP7_75t_SL g1421 ( 
.A(n_1001),
.B(n_91),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1076),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1076),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1079),
.B(n_91),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1076),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1076),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1076),
.Y(n_1427)
);

XOR2xp5_ASAP7_75t_L g1428 ( 
.A(n_1001),
.B(n_92),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1079),
.B(n_92),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1085),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1076),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1076),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1149),
.B(n_244),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1076),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1079),
.B(n_94),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1080),
.B(n_94),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1076),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1076),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1430),
.B(n_95),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1170),
.Y(n_1440)
);

OR2x2_ASAP7_75t_SL g1441 ( 
.A(n_1405),
.B(n_96),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1170),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1416),
.B(n_98),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1416),
.B(n_98),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1420),
.B(n_100),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1186),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1171),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1389),
.B(n_100),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1172),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1190),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1420),
.B(n_101),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1200),
.B(n_102),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1296),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1359),
.B(n_103),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1302),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1279),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1337),
.B(n_103),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1173),
.A2(n_249),
.B(n_246),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1206),
.B(n_105),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1359),
.B(n_105),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1271),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1296),
.B(n_1214),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1271),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1191),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1210),
.B(n_106),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1187),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1271),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1213),
.B(n_106),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1337),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1183),
.B(n_107),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1290),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1294),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1336),
.B(n_107),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1209),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1229),
.B(n_109),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1372),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1219),
.B(n_112),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1187),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1424),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1201),
.B(n_113),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1203),
.B(n_114),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1236),
.B(n_116),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1202),
.B(n_116),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1212),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1212),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1173),
.A2(n_348),
.B(n_479),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1217),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1192),
.A2(n_346),
.B(n_478),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1177),
.B(n_117),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1292),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1217),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1230),
.B(n_117),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1193),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1303),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1231),
.B(n_118),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1233),
.B(n_120),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1185),
.B(n_120),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1197),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1199),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1182),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1239),
.B(n_122),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1429),
.B(n_125),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1254),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1435),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1245),
.B(n_125),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1241),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1295),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1205),
.A2(n_351),
.B(n_476),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1406),
.B(n_126),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1323),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1261),
.B(n_127),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1258),
.B(n_127),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1325),
.Y(n_1515)
);

AND2x2_ASAP7_75t_SL g1516 ( 
.A(n_1261),
.B(n_1280),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1254),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1241),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1316),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1412),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1412),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1311),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1246),
.B(n_128),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1277),
.B(n_131),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1358),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1326),
.B(n_131),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1249),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1383),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1334),
.B(n_132),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1362),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1205),
.A2(n_357),
.B(n_471),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1208),
.B(n_134),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1414),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1414),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1241),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1382),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1224),
.B(n_134),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1365),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1227),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1436),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1238),
.B(n_135),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1192),
.A2(n_361),
.B(n_468),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1436),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1384),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1300),
.B(n_136),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1226),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1309),
.B(n_136),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1385),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1250),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1326),
.B(n_137),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1332),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1368),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1378),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1175),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1226),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1350),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1376),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1174),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1227),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1394),
.B(n_138),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1398),
.B(n_141),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1176),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1264),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1215),
.Y(n_1564)
);

AND2x2_ASAP7_75t_SL g1565 ( 
.A(n_1305),
.B(n_141),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1253),
.B(n_143),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1215),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1242),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1318),
.B(n_144),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1195),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1354),
.B(n_146),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1315),
.B(n_148),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1380),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1178),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1318),
.B(n_149),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1410),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1301),
.B(n_151),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1242),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1413),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1274),
.B(n_151),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1417),
.B(n_152),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1270),
.B(n_152),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1377),
.B(n_153),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1260),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1251),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1381),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_SL g1587 ( 
.A(n_1285),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1419),
.B(n_154),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1422),
.B(n_154),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1423),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1319),
.B(n_250),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1421),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1289),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1400),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1425),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1343),
.A2(n_1344),
.B(n_1341),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1319),
.B(n_481),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1426),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1427),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1431),
.B(n_252),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1216),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1432),
.B(n_466),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1434),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1371),
.B(n_256),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1437),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1176),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1438),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1327),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1256),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1272),
.B(n_260),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1273),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1176),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1330),
.B(n_263),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1176),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1179),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1346),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1180),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1181),
.B(n_465),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1269),
.B(n_266),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1386),
.B(n_1306),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1223),
.B(n_463),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1392),
.B(n_269),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1287),
.B(n_457),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1194),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1278),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1252),
.B(n_276),
.Y(n_1626)
);

AND2x2_ASAP7_75t_SL g1627 ( 
.A(n_1310),
.B(n_1284),
.Y(n_1627)
);

BUFx5_ASAP7_75t_L g1628 ( 
.A(n_1247),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1255),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1283),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1243),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1257),
.B(n_454),
.Y(n_1632)
);

INVx4_ASAP7_75t_L g1633 ( 
.A(n_1247),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1298),
.Y(n_1634)
);

AND2x6_ASAP7_75t_L g1635 ( 
.A(n_1244),
.B(n_1313),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1317),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1393),
.B(n_279),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1411),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1307),
.B(n_452),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1357),
.A2(n_1409),
.B(n_1408),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1345),
.B(n_281),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1275),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1262),
.B(n_282),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1400),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1345),
.B(n_283),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1388),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1308),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1402),
.A2(n_284),
.B(n_287),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1349),
.B(n_450),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1263),
.B(n_288),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1184),
.B(n_449),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1355),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1428),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1328),
.B(n_294),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1265),
.B(n_448),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1266),
.B(n_304),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1288),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1267),
.B(n_1268),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1247),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1401),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1361),
.B(n_447),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1198),
.B(n_305),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1169),
.A2(n_306),
.B(n_310),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1415),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1218),
.B(n_446),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1366),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1221),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1228),
.B(n_311),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1370),
.B(n_445),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1247),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1248),
.B(n_319),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1320),
.B(n_320),
.Y(n_1672)
);

NOR2xp67_ASAP7_75t_L g1673 ( 
.A(n_1356),
.B(n_322),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1314),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1418),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1169),
.A2(n_323),
.B(n_324),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1222),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1196),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1374),
.B(n_444),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1351),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1349),
.B(n_327),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1314),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1379),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1369),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1387),
.B(n_1399),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1339),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1342),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1375),
.B(n_328),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1324),
.B(n_1188),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1360),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1403),
.B(n_337),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1397),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1369),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1304),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1391),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1297),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1297),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1407),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1232),
.B(n_442),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1235),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1404),
.B(n_1259),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1333),
.B(n_338),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1338),
.B(n_340),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1329),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1352),
.B(n_1312),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1321),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1276),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1395),
.B(n_1335),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1363),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1340),
.B(n_342),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1322),
.B(n_349),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1390),
.B(n_354),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1286),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1396),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1331),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1211),
.B(n_440),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1220),
.B(n_356),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1331),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1433),
.B(n_439),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1364),
.A2(n_368),
.B(n_370),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1340),
.B(n_373),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1433),
.B(n_438),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1282),
.B(n_1364),
.Y(n_1723)
);

AND2x2_ASAP7_75t_SL g1724 ( 
.A(n_1281),
.B(n_374),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1507),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1502),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1443),
.B(n_1299),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1615),
.Y(n_1728)
);

AND2x6_ASAP7_75t_L g1729 ( 
.A(n_1610),
.B(n_1367),
.Y(n_1729)
);

BUFx2_ASAP7_75t_SL g1730 ( 
.A(n_1610),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1519),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1666),
.B(n_1373),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1443),
.B(n_1299),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1526),
.B(n_1348),
.Y(n_1734)
);

INVx6_ASAP7_75t_L g1735 ( 
.A(n_1507),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1584),
.B(n_1281),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1674),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1642),
.B(n_1348),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_SL g1739 ( 
.A(n_1513),
.B(n_1353),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1642),
.B(n_1189),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1462),
.B(n_1293),
.Y(n_1741)
);

BUFx4f_ASAP7_75t_L g1742 ( 
.A(n_1513),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1594),
.B(n_1204),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1564),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1507),
.B(n_1291),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1477),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1513),
.B(n_1207),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1508),
.Y(n_1748)
);

BUFx8_ASAP7_75t_SL g1749 ( 
.A(n_1475),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1526),
.B(n_1293),
.Y(n_1750)
);

CKINVDCx16_ASAP7_75t_R g1751 ( 
.A(n_1464),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1454),
.B(n_1225),
.Y(n_1752)
);

INVx6_ASAP7_75t_SL g1753 ( 
.A(n_1458),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1477),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1564),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1567),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1594),
.B(n_1240),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1567),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1472),
.Y(n_1759)
);

BUFx4f_ASAP7_75t_L g1760 ( 
.A(n_1458),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1517),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1568),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1528),
.B(n_1353),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1528),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1470),
.B(n_1478),
.Y(n_1765)
);

NAND2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1458),
.B(n_1353),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1685),
.B(n_1237),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1472),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1724),
.B(n_1347),
.Y(n_1769)
);

OR2x6_ASAP7_75t_L g1770 ( 
.A(n_1464),
.B(n_1347),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1568),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1617),
.Y(n_1772)
);

AND2x6_ASAP7_75t_L g1773 ( 
.A(n_1610),
.B(n_1347),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1674),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1444),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1674),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1508),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1724),
.B(n_1234),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1470),
.B(n_437),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1578),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1478),
.B(n_375),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1546),
.B(n_380),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1454),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1445),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1522),
.Y(n_1785)
);

NAND2xp33_ASAP7_75t_L g1786 ( 
.A(n_1628),
.B(n_382),
.Y(n_1786)
);

AND2x6_ASAP7_75t_L g1787 ( 
.A(n_1643),
.B(n_383),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1581),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1468),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1578),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1546),
.B(n_388),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1631),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1674),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1546),
.B(n_390),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1685),
.B(n_1704),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1695),
.B(n_393),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1550),
.B(n_396),
.Y(n_1797)
);

INVx4_ASAP7_75t_L g1798 ( 
.A(n_1508),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1588),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1584),
.B(n_397),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1589),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1440),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1555),
.B(n_435),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1508),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1658),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1440),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1442),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1683),
.B(n_399),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1485),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1518),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1518),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1455),
.B(n_403),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1554),
.B(n_404),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1555),
.B(n_434),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1638),
.B(n_405),
.Y(n_1815)
);

NAND2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1555),
.B(n_406),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1518),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1518),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1631),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1468),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1551),
.B(n_412),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1551),
.B(n_431),
.Y(n_1822)
);

NAND2x1p5_ASAP7_75t_L g1823 ( 
.A(n_1534),
.B(n_414),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1442),
.Y(n_1824)
);

OR2x6_ASAP7_75t_L g1825 ( 
.A(n_1463),
.B(n_417),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1461),
.B(n_421),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1522),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1608),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1687),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1592),
.B(n_424),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1558),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1561),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1692),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1506),
.B(n_428),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_SL g1835 ( 
.A(n_1616),
.B(n_430),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1534),
.B(n_1473),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1706),
.B(n_1660),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1616),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1687),
.Y(n_1839)
);

AND2x2_ASAP7_75t_SL g1840 ( 
.A(n_1643),
.B(n_1650),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1574),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1692),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1596),
.B(n_1481),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1463),
.Y(n_1844)
);

INVx6_ASAP7_75t_L g1845 ( 
.A(n_1473),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1643),
.B(n_1650),
.Y(n_1846)
);

AND2x6_ASAP7_75t_L g1847 ( 
.A(n_1650),
.B(n_1672),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1517),
.Y(n_1848)
);

NAND2x1p5_ASAP7_75t_L g1849 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1849)
);

BUFx4f_ASAP7_75t_L g1850 ( 
.A(n_1523),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1481),
.B(n_1660),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1723),
.B(n_1547),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1483),
.B(n_1482),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1509),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1553),
.B(n_1573),
.Y(n_1855)
);

NAND2x1p5_ASAP7_75t_L g1856 ( 
.A(n_1523),
.B(n_1535),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1448),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1647),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1698),
.Y(n_1859)
);

INVx4_ASAP7_75t_L g1860 ( 
.A(n_1535),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1651),
.B(n_1572),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1662),
.B(n_1671),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1448),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1690),
.B(n_1565),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1553),
.B(n_1573),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1638),
.B(n_1678),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1570),
.B(n_1601),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1576),
.B(n_1579),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1450),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1590),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1657),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1698),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1595),
.B(n_1598),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1875)
);

BUFx12f_ASAP7_75t_L g1876 ( 
.A(n_1690),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1605),
.B(n_1607),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1450),
.Y(n_1878)
);

NAND2x1p5_ASAP7_75t_L g1879 ( 
.A(n_1523),
.B(n_1535),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1525),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1624),
.B(n_1705),
.Y(n_1881)
);

BUFx12f_ASAP7_75t_L g1882 ( 
.A(n_1441),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1586),
.B(n_1593),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1715),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1715),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1587),
.B(n_1624),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1672),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1525),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1586),
.B(n_1593),
.Y(n_1889)
);

AND2x2_ASAP7_75t_SL g1890 ( 
.A(n_1561),
.B(n_1565),
.Y(n_1890)
);

INVx5_ASAP7_75t_L g1891 ( 
.A(n_1561),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1521),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1530),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1587),
.B(n_1539),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1530),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1539),
.B(n_1559),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1686),
.B(n_1653),
.Y(n_1897)
);

BUFx12f_ASAP7_75t_L g1898 ( 
.A(n_1582),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1686),
.B(n_1653),
.Y(n_1899)
);

BUFx4f_ASAP7_75t_L g1900 ( 
.A(n_1582),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1538),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1446),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1536),
.B(n_1544),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1538),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1479),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1668),
.B(n_1712),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1559),
.B(n_1644),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1552),
.Y(n_1908)
);

INVx4_ASAP7_75t_L g1909 ( 
.A(n_1582),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1552),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1479),
.B(n_1489),
.Y(n_1911)
);

CKINVDCx8_ASAP7_75t_R g1912 ( 
.A(n_1479),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1493),
.B(n_1521),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1672),
.B(n_1520),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1540),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1520),
.B(n_1533),
.Y(n_1916)
);

INVx4_ASAP7_75t_L g1917 ( 
.A(n_1633),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1548),
.B(n_1556),
.Y(n_1918)
);

INVx5_ASAP7_75t_L g1919 ( 
.A(n_1562),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1613),
.B(n_1566),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1680),
.B(n_1512),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1629),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1515),
.B(n_1620),
.Y(n_1923)
);

AND2x6_ASAP7_75t_L g1924 ( 
.A(n_1659),
.B(n_1670),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1471),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1580),
.B(n_1453),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1675),
.B(n_1533),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1701),
.B(n_1714),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_SL g1929 ( 
.A(n_1633),
.B(n_1563),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1452),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1527),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1545),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1540),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1456),
.B(n_1496),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1702),
.B(n_1571),
.Y(n_1935)
);

CKINVDCx8_ASAP7_75t_R g1936 ( 
.A(n_1635),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1456),
.B(n_1496),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1532),
.B(n_1639),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1537),
.B(n_1691),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1484),
.B(n_1716),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1560),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1543),
.B(n_1516),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1543),
.B(n_1516),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1439),
.Y(n_1944)
);

NAND2x1_ASAP7_75t_L g1945 ( 
.A(n_1635),
.B(n_1682),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1467),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1527),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1447),
.B(n_1451),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1708),
.B(n_1511),
.Y(n_1949)
);

INVx5_ASAP7_75t_L g1950 ( 
.A(n_1562),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1717),
.B(n_1675),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1514),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1524),
.B(n_1491),
.Y(n_1953)
);

OR2x6_ASAP7_75t_SL g1954 ( 
.A(n_1654),
.B(n_1569),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1689),
.B(n_1524),
.Y(n_1955)
);

INVx6_ASAP7_75t_SL g1956 ( 
.A(n_1563),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1467),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1467),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1499),
.B(n_1529),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_SL g1960 ( 
.A(n_1633),
.B(n_1664),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1577),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1467),
.Y(n_1962)
);

NAND2x1_ASAP7_75t_L g1963 ( 
.A(n_1635),
.B(n_1682),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1465),
.B(n_1495),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1693),
.B(n_1583),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1541),
.B(n_1474),
.Y(n_1966)
);

BUFx12f_ASAP7_75t_L g1967 ( 
.A(n_1635),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1583),
.B(n_1661),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1664),
.B(n_1627),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1627),
.B(n_1684),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1505),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1667),
.B(n_1707),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1575),
.B(n_1449),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1659),
.B(n_1670),
.Y(n_1975)
);

OR2x6_ASAP7_75t_L g1976 ( 
.A(n_1665),
.B(n_1562),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1646),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1684),
.B(n_1619),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1623),
.B(n_1504),
.Y(n_1979)
);

AO21x2_ASAP7_75t_L g1980 ( 
.A1(n_1649),
.A2(n_1681),
.B(n_1710),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1635),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1480),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1557),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1646),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1505),
.B(n_1628),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1707),
.B(n_1713),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1480),
.Y(n_1987)
);

NAND2x1_ASAP7_75t_SL g1988 ( 
.A(n_1721),
.B(n_1703),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1549),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1677),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1549),
.B(n_1460),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1641),
.B(n_1645),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1677),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1480),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1466),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1480),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1606),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1606),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1713),
.B(n_1700),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1469),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1637),
.B(n_1606),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1476),
.B(n_1494),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1585),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1585),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1609),
.Y(n_2005)
);

INVx4_ASAP7_75t_L g2006 ( 
.A(n_1612),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1497),
.B(n_1503),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1498),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1696),
.B(n_1697),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1609),
.B(n_1611),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1626),
.B(n_1688),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1688),
.B(n_1703),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1711),
.B(n_1656),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1711),
.B(n_1655),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1611),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1600),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1602),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1625),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1604),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1604),
.B(n_1697),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1612),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1625),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1669),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1696),
.B(n_1709),
.Y(n_2024)
);

OR2x6_ASAP7_75t_L g2025 ( 
.A(n_1612),
.B(n_1614),
.Y(n_2025)
);

OR2x6_ASAP7_75t_L g2026 ( 
.A(n_1614),
.B(n_1490),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1630),
.B(n_1636),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1630),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1709),
.B(n_1640),
.Y(n_2029)
);

BUFx12f_ASAP7_75t_L g2030 ( 
.A(n_1785),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1753),
.Y(n_2031)
);

CKINVDCx20_ASAP7_75t_R g2032 ( 
.A(n_1749),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1840),
.Y(n_2033)
);

BUFx4f_ASAP7_75t_SL g2034 ( 
.A(n_1876),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1833),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1847),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2010),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2027),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1839),
.Y(n_2039)
);

BUFx12f_ASAP7_75t_L g2040 ( 
.A(n_1827),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1795),
.B(n_1694),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_1847),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1928),
.B(n_1636),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1936),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1882),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1839),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1847),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1859),
.Y(n_2048)
);

INVx3_ASAP7_75t_L g2049 ( 
.A(n_1847),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_1900),
.Y(n_2050)
);

BUFx2_ASAP7_75t_SL g2051 ( 
.A(n_1912),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1890),
.A2(n_1710),
.B1(n_1614),
.B2(n_1628),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1753),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_1730),
.Y(n_2054)
);

BUFx2_ASAP7_75t_R g2055 ( 
.A(n_1838),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_1730),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_SL g2057 ( 
.A(n_1745),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1972),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_1967),
.Y(n_2059)
);

INVx6_ASAP7_75t_L g2060 ( 
.A(n_1873),
.Y(n_2060)
);

BUFx4f_ASAP7_75t_SL g2061 ( 
.A(n_1956),
.Y(n_2061)
);

AO21x2_ASAP7_75t_L g2062 ( 
.A1(n_1750),
.A2(n_1681),
.B(n_1459),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_1868),
.Y(n_2063)
);

BUFx2_ASAP7_75t_SL g2064 ( 
.A(n_1891),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1742),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1888),
.Y(n_2066)
);

BUFx12f_ASAP7_75t_L g2067 ( 
.A(n_1842),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1888),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_1858),
.Y(n_2069)
);

INVx8_ASAP7_75t_L g2070 ( 
.A(n_1745),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1895),
.Y(n_2071)
);

INVxp33_ASAP7_75t_L g2072 ( 
.A(n_1764),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1895),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1900),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1742),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_1760),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1910),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1737),
.Y(n_2078)
);

NAND2x1p5_ASAP7_75t_L g2079 ( 
.A(n_1760),
.B(n_1682),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_1845),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1910),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1850),
.B(n_1614),
.Y(n_2082)
);

INVx6_ASAP7_75t_L g2083 ( 
.A(n_1845),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1917),
.Y(n_2084)
);

INVx3_ASAP7_75t_SL g2085 ( 
.A(n_1735),
.Y(n_2085)
);

INVx6_ASAP7_75t_SL g2086 ( 
.A(n_1825),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1843),
.B(n_1679),
.Y(n_2087)
);

BUFx12f_ASAP7_75t_L g2088 ( 
.A(n_1731),
.Y(n_2088)
);

INVx6_ASAP7_75t_SL g2089 ( 
.A(n_1825),
.Y(n_2089)
);

INVx5_ASAP7_75t_L g2090 ( 
.A(n_1747),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1725),
.Y(n_2091)
);

BUFx8_ASAP7_75t_L g2092 ( 
.A(n_1898),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1737),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1744),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1744),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1747),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1756),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1756),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1790),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1759),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1848),
.Y(n_2101)
);

INVxp67_ASAP7_75t_SL g2102 ( 
.A(n_1850),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1768),
.Y(n_2103)
);

NAND2x1p5_ASAP7_75t_L g2104 ( 
.A(n_1891),
.B(n_1490),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1790),
.Y(n_2105)
);

INVx4_ASAP7_75t_L g2106 ( 
.A(n_1891),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_SL g2107 ( 
.A(n_1927),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1854),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1735),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1909),
.B(n_1597),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1844),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1917),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1983),
.B(n_1935),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_1909),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1765),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1945),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1765),
.Y(n_2117)
);

HB1xp67_ASAP7_75t_L g2118 ( 
.A(n_2005),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_1907),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1802),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1836),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2028),
.Y(n_2122)
);

INVx5_ASAP7_75t_L g2123 ( 
.A(n_1787),
.Y(n_2123)
);

BUFx12f_ASAP7_75t_L g2124 ( 
.A(n_1867),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1806),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_1865),
.A2(n_1955),
.B1(n_1940),
.B2(n_1861),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1807),
.Y(n_2127)
);

BUFx12f_ASAP7_75t_L g2128 ( 
.A(n_1897),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1824),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1755),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1758),
.Y(n_2131)
);

CKINVDCx6p67_ASAP7_75t_R g2132 ( 
.A(n_1751),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1762),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1771),
.Y(n_2134)
);

INVxp67_ASAP7_75t_SL g2135 ( 
.A(n_1846),
.Y(n_2135)
);

INVx8_ASAP7_75t_L g2136 ( 
.A(n_1787),
.Y(n_2136)
);

CKINVDCx20_ASAP7_75t_R g2137 ( 
.A(n_1789),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1843),
.B(n_1591),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1780),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_1761),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_1773),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1829),
.Y(n_2142)
);

BUFx2_ASAP7_75t_SL g2143 ( 
.A(n_1787),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1880),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1852),
.B(n_1652),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1849),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_1939),
.A2(n_1628),
.B1(n_1632),
.B2(n_1488),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_1951),
.A2(n_1628),
.B1(n_1622),
.B2(n_1510),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_1956),
.Y(n_2149)
);

INVx4_ASAP7_75t_L g2150 ( 
.A(n_1787),
.Y(n_2150)
);

INVx6_ASAP7_75t_L g2151 ( 
.A(n_1907),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1774),
.Y(n_2152)
);

CKINVDCx20_ASAP7_75t_R g2153 ( 
.A(n_1820),
.Y(n_2153)
);

BUFx2_ASAP7_75t_SL g2154 ( 
.A(n_1779),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1883),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1893),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1881),
.B(n_1634),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1945),
.Y(n_2158)
);

BUFx4f_ASAP7_75t_L g2159 ( 
.A(n_1773),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1901),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1904),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1908),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_1773),
.Y(n_2163)
);

NAND2x1p5_ASAP7_75t_L g2164 ( 
.A(n_1919),
.B(n_1542),
.Y(n_2164)
);

BUFx2_ASAP7_75t_L g2165 ( 
.A(n_1927),
.Y(n_2165)
);

INVx5_ASAP7_75t_L g2166 ( 
.A(n_1773),
.Y(n_2166)
);

BUFx2_ASAP7_75t_SL g2167 ( 
.A(n_1779),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_1781),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1774),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_1883),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1853),
.B(n_1923),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1774),
.Y(n_2172)
);

CKINVDCx20_ASAP7_75t_R g2173 ( 
.A(n_1899),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1886),
.Y(n_2174)
);

INVx4_ASAP7_75t_L g2175 ( 
.A(n_1919),
.Y(n_2175)
);

INVx4_ASAP7_75t_L g2176 ( 
.A(n_1919),
.Y(n_2176)
);

INVx2_ASAP7_75t_R g2177 ( 
.A(n_1950),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1746),
.Y(n_2178)
);

INVx5_ASAP7_75t_L g2179 ( 
.A(n_1810),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1754),
.Y(n_2180)
);

NAND2x1p5_ASAP7_75t_L g2181 ( 
.A(n_1950),
.B(n_1542),
.Y(n_2181)
);

BUFx12f_ASAP7_75t_L g2182 ( 
.A(n_1815),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1776),
.Y(n_2183)
);

INVx3_ASAP7_75t_SL g2184 ( 
.A(n_1889),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1872),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1872),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1857),
.Y(n_2187)
);

INVx8_ASAP7_75t_L g2188 ( 
.A(n_1889),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_1781),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1863),
.Y(n_2190)
);

NAND2x1p5_ASAP7_75t_L g2191 ( 
.A(n_1950),
.B(n_1634),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1862),
.B(n_1732),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1906),
.B(n_1618),
.Y(n_2193)
);

INVx6_ASAP7_75t_SL g2194 ( 
.A(n_1803),
.Y(n_2194)
);

BUFx10_ASAP7_75t_L g2195 ( 
.A(n_1803),
.Y(n_2195)
);

CKINVDCx11_ASAP7_75t_R g2196 ( 
.A(n_1954),
.Y(n_2196)
);

CKINVDCx6p67_ASAP7_75t_R g2197 ( 
.A(n_1941),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_1855),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_1934),
.B(n_1673),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1932),
.Y(n_2200)
);

BUFx3_ASAP7_75t_L g2201 ( 
.A(n_1977),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1776),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1776),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1793),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1870),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_1989),
.Y(n_2206)
);

INVx1_ASAP7_75t_SL g2207 ( 
.A(n_1994),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1934),
.B(n_1621),
.Y(n_2208)
);

CKINVDCx5p33_ASAP7_75t_R g2209 ( 
.A(n_1949),
.Y(n_2209)
);

BUFx4_ASAP7_75t_SL g2210 ( 
.A(n_1770),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1878),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_1855),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_1866),
.Y(n_2213)
);

BUFx2_ASAP7_75t_SL g2214 ( 
.A(n_1814),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1986),
.B(n_1719),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1851),
.B(n_1652),
.Y(n_2216)
);

BUFx4f_ASAP7_75t_L g2217 ( 
.A(n_1856),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1866),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_1937),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2018),
.Y(n_2220)
);

INVx5_ASAP7_75t_L g2221 ( 
.A(n_1810),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1937),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1726),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1728),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_1948),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1772),
.Y(n_2226)
);

INVx5_ASAP7_75t_L g2227 ( 
.A(n_1810),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_1896),
.Y(n_2228)
);

BUFx12f_ASAP7_75t_L g2229 ( 
.A(n_1814),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_1896),
.Y(n_2230)
);

INVx5_ASAP7_75t_L g2231 ( 
.A(n_1817),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1793),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1805),
.B(n_1628),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1792),
.Y(n_2234)
);

BUFx2_ASAP7_75t_SL g2235 ( 
.A(n_1834),
.Y(n_2235)
);

BUFx3_ASAP7_75t_L g2236 ( 
.A(n_1996),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_1963),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1851),
.B(n_1720),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_1948),
.Y(n_2239)
);

NAND2x1p5_ASAP7_75t_L g2240 ( 
.A(n_1963),
.B(n_1720),
.Y(n_2240)
);

INVx4_ASAP7_75t_L g2241 ( 
.A(n_1887),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_1879),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_1757),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1792),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2003),
.Y(n_2245)
);

BUFx12f_ASAP7_75t_L g2246 ( 
.A(n_1813),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1975),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1959),
.B(n_1828),
.Y(n_2248)
);

NAND2x1p5_ASAP7_75t_L g2249 ( 
.A(n_1887),
.B(n_1718),
.Y(n_2249)
);

OR2x6_ASAP7_75t_L g2250 ( 
.A(n_1911),
.B(n_1531),
.Y(n_2250)
);

BUFx2_ASAP7_75t_SL g2251 ( 
.A(n_1834),
.Y(n_2251)
);

INVx3_ASAP7_75t_SL g2252 ( 
.A(n_1770),
.Y(n_2252)
);

CKINVDCx11_ASAP7_75t_R g2253 ( 
.A(n_2025),
.Y(n_2253)
);

CKINVDCx20_ASAP7_75t_R g2254 ( 
.A(n_2032),
.Y(n_2254)
);

CKINVDCx11_ASAP7_75t_R g2255 ( 
.A(n_2030),
.Y(n_2255)
);

BUFx2_ASAP7_75t_SL g2256 ( 
.A(n_2057),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2039),
.Y(n_2257)
);

OAI21xp33_ASAP7_75t_SL g2258 ( 
.A1(n_2150),
.A2(n_1914),
.B(n_1988),
.Y(n_2258)
);

CKINVDCx11_ASAP7_75t_R g2259 ( 
.A(n_2040),
.Y(n_2259)
);

INVx6_ASAP7_75t_L g2260 ( 
.A(n_2092),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2223),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_2092),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2188),
.Y(n_2263)
);

INVx4_ASAP7_75t_L g2264 ( 
.A(n_2136),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2094),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2039),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2086),
.A2(n_1778),
.B1(n_1769),
.B2(n_1887),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2086),
.A2(n_1832),
.B1(n_1905),
.B2(n_1835),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2171),
.B(n_1831),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_2034),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2063),
.B(n_1841),
.Y(n_2271)
);

CKINVDCx6p67_ASAP7_75t_R g2272 ( 
.A(n_2132),
.Y(n_2272)
);

BUFx3_ASAP7_75t_L g2273 ( 
.A(n_2048),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2113),
.A2(n_1999),
.B1(n_1920),
.B2(n_1942),
.Y(n_2274)
);

OAI21xp33_ASAP7_75t_SL g2275 ( 
.A1(n_2150),
.A2(n_1988),
.B(n_1741),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2154),
.A2(n_2014),
.B1(n_2013),
.B2(n_2012),
.Y(n_2276)
);

BUFx2_ASAP7_75t_SL g2277 ( 
.A(n_2057),
.Y(n_2277)
);

BUFx3_ASAP7_75t_L g2278 ( 
.A(n_2103),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2095),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_2089),
.Y(n_2280)
);

INVx5_ASAP7_75t_L g2281 ( 
.A(n_2136),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2099),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2223),
.Y(n_2283)
);

OAI21xp5_ASAP7_75t_SL g2284 ( 
.A1(n_2168),
.A2(n_1830),
.B(n_1736),
.Y(n_2284)
);

AOI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2196),
.A2(n_2089),
.B1(n_2126),
.B2(n_2192),
.Y(n_2285)
);

BUFx8_ASAP7_75t_L g2286 ( 
.A(n_2067),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_2167),
.A2(n_1968),
.B1(n_2011),
.B2(n_1965),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2224),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_2188),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2078),
.Y(n_2290)
);

BUFx12f_ASAP7_75t_L g2291 ( 
.A(n_2045),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_2194),
.Y(n_2292)
);

CKINVDCx6p67_ASAP7_75t_R g2293 ( 
.A(n_2085),
.Y(n_2293)
);

NAND2x1p5_ASAP7_75t_L g2294 ( 
.A(n_2166),
.B(n_1821),
.Y(n_2294)
);

INVx6_ASAP7_75t_L g2295 ( 
.A(n_2060),
.Y(n_2295)
);

OAI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_2189),
.A2(n_1905),
.B1(n_1978),
.B2(n_1960),
.Y(n_2296)
);

INVx6_ASAP7_75t_L g2297 ( 
.A(n_2060),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2128),
.A2(n_1953),
.B1(n_1969),
.B2(n_1729),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2070),
.A2(n_1729),
.B1(n_1944),
.B2(n_2009),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2063),
.B(n_1871),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_2194),
.Y(n_2301)
);

BUFx4f_ASAP7_75t_SL g2302 ( 
.A(n_2088),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2105),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2070),
.A2(n_1729),
.B1(n_1995),
.B2(n_2008),
.Y(n_2304)
);

INVx6_ASAP7_75t_L g2305 ( 
.A(n_2035),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2229),
.A2(n_2136),
.B1(n_2058),
.B2(n_2209),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_SL g2307 ( 
.A(n_2055),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_2083),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2066),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2081),
.Y(n_2310)
);

BUFx12f_ASAP7_75t_L g2311 ( 
.A(n_2253),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_L g2312 ( 
.A(n_2078),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2037),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2078),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2173),
.A2(n_1729),
.B1(n_1995),
.B2(n_2008),
.Y(n_2315)
);

CKINVDCx11_ASAP7_75t_R g2316 ( 
.A(n_2124),
.Y(n_2316)
);

INVx8_ASAP7_75t_L g2317 ( 
.A(n_2090),
.Y(n_2317)
);

BUFx10_ASAP7_75t_L g2318 ( 
.A(n_2107),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2038),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_2166),
.Y(n_2320)
);

BUFx2_ASAP7_75t_SL g2321 ( 
.A(n_2107),
.Y(n_2321)
);

BUFx2_ASAP7_75t_L g2322 ( 
.A(n_2137),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2235),
.A2(n_2000),
.B1(n_1992),
.B2(n_1938),
.Y(n_2323)
);

AOI22xp33_ASAP7_75t_L g2324 ( 
.A1(n_2251),
.A2(n_2000),
.B1(n_1992),
.B2(n_1938),
.Y(n_2324)
);

BUFx4f_ASAP7_75t_L g2325 ( 
.A(n_2036),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2224),
.Y(n_2326)
);

BUFx12f_ASAP7_75t_L g2327 ( 
.A(n_2200),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2215),
.A2(n_1952),
.B1(n_1925),
.B2(n_1943),
.Y(n_2328)
);

BUFx12f_ASAP7_75t_L g2329 ( 
.A(n_2065),
.Y(n_2329)
);

CKINVDCx11_ASAP7_75t_R g2330 ( 
.A(n_2153),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_2093),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2033),
.A2(n_1926),
.B1(n_1966),
.B2(n_1979),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2226),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2214),
.A2(n_1822),
.B1(n_1821),
.B2(n_2019),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2248),
.B(n_1869),
.Y(n_2335)
);

CKINVDCx20_ASAP7_75t_R g2336 ( 
.A(n_2197),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2033),
.A2(n_2193),
.B1(n_2182),
.B2(n_2246),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2143),
.A2(n_1822),
.B1(n_1902),
.B2(n_1733),
.Y(n_2338)
);

AOI22xp33_ASAP7_75t_SL g2339 ( 
.A1(n_2123),
.A2(n_1739),
.B1(n_1929),
.B2(n_1985),
.Y(n_2339)
);

INVx8_ASAP7_75t_L g2340 ( 
.A(n_2090),
.Y(n_2340)
);

CKINVDCx11_ASAP7_75t_R g2341 ( 
.A(n_2184),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2123),
.B(n_1739),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2046),
.Y(n_2343)
);

CKINVDCx20_ASAP7_75t_R g2344 ( 
.A(n_2061),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2041),
.B(n_1874),
.Y(n_2345)
);

AOI21x1_ASAP7_75t_L g2346 ( 
.A1(n_2250),
.A2(n_2026),
.B(n_1734),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2043),
.B(n_1964),
.Y(n_2347)
);

BUFx2_ASAP7_75t_SL g2348 ( 
.A(n_2123),
.Y(n_2348)
);

INVx4_ASAP7_75t_L g2349 ( 
.A(n_2166),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_2033),
.A2(n_1974),
.B1(n_1973),
.B2(n_1738),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2097),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_SL g2352 ( 
.A1(n_2051),
.A2(n_1800),
.B1(n_1894),
.B2(n_1924),
.Y(n_2352)
);

INVx6_ASAP7_75t_L g2353 ( 
.A(n_2083),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2145),
.B(n_1875),
.Y(n_2354)
);

OAI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2058),
.A2(n_1970),
.B1(n_1763),
.B2(n_1727),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2087),
.A2(n_1738),
.B1(n_2007),
.B2(n_2002),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2174),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2046),
.Y(n_2358)
);

OAI21xp5_ASAP7_75t_SL g2359 ( 
.A1(n_2042),
.A2(n_2049),
.B(n_2047),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2068),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_2069),
.A2(n_2023),
.B1(n_2029),
.B2(n_2020),
.Y(n_2361)
);

CKINVDCx6p67_ASAP7_75t_R g2362 ( 
.A(n_2090),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2108),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2234),
.B(n_1877),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2234),
.B(n_1903),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2225),
.A2(n_1784),
.B1(n_1775),
.B2(n_1783),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2093),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2093),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2239),
.A2(n_1930),
.B1(n_1913),
.B2(n_1837),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2097),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2210),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2111),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2226),
.Y(n_2373)
);

BUFx10_ASAP7_75t_L g2374 ( 
.A(n_2075),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2159),
.A2(n_1766),
.B1(n_1991),
.B2(n_1794),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2185),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2185),
.Y(n_2377)
);

OAI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2140),
.A2(n_1915),
.B1(n_1933),
.B2(n_1767),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2098),
.Y(n_2379)
);

BUFx12f_ASAP7_75t_L g2380 ( 
.A(n_2149),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2165),
.A2(n_2017),
.B1(n_2016),
.B2(n_1808),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_L g2382 ( 
.A1(n_2276),
.A2(n_2101),
.B1(n_2138),
.B2(n_2216),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2285),
.A2(n_2195),
.B1(n_2049),
.B2(n_2186),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2261),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2322),
.B(n_2072),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2283),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2288),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2347),
.B(n_2134),
.Y(n_2388)
);

AOI22xp33_ASAP7_75t_SL g2389 ( 
.A1(n_2334),
.A2(n_2195),
.B1(n_2042),
.B2(n_2047),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_2332),
.A2(n_2186),
.B1(n_2244),
.B2(n_2047),
.Y(n_2390)
);

AOI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2328),
.A2(n_2244),
.B1(n_2036),
.B2(n_2096),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2326),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2356),
.A2(n_2287),
.B1(n_2378),
.B2(n_2315),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2306),
.B(n_2036),
.Y(n_2394)
);

OAI21xp33_ASAP7_75t_L g2395 ( 
.A1(n_2274),
.A2(n_2091),
.B(n_2135),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2284),
.A2(n_2159),
.B1(n_2056),
.B2(n_2054),
.Y(n_2396)
);

AOI22xp33_ASAP7_75t_SL g2397 ( 
.A1(n_2352),
.A2(n_2064),
.B1(n_2054),
.B2(n_2056),
.Y(n_2397)
);

OAI222xp33_ASAP7_75t_L g2398 ( 
.A1(n_2264),
.A2(n_2206),
.B1(n_2250),
.B2(n_2207),
.C1(n_2071),
.C2(n_2073),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2330),
.B(n_2329),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2336),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2265),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2279),
.Y(n_2402)
);

AOI22xp5_ASAP7_75t_SL g2403 ( 
.A1(n_2344),
.A2(n_2059),
.B1(n_2074),
.B2(n_2050),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2341),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2313),
.B(n_2098),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2357),
.B(n_2100),
.Y(n_2406)
);

OAI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2350),
.A2(n_2206),
.B1(n_2122),
.B2(n_2115),
.Y(n_2407)
);

OAI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2381),
.A2(n_2122),
.B1(n_2117),
.B2(n_2052),
.Y(n_2408)
);

NAND3xp33_ASAP7_75t_L g2409 ( 
.A(n_2361),
.B(n_1809),
.C(n_2118),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2333),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_SL g2411 ( 
.A1(n_2264),
.A2(n_2102),
.B1(n_2076),
.B2(n_2151),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2282),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2257),
.Y(n_2413)
);

NAND3xp33_ASAP7_75t_L g2414 ( 
.A(n_2337),
.B(n_1799),
.C(n_1788),
.Y(n_2414)
);

OAI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2281),
.A2(n_2073),
.B1(n_2071),
.B2(n_2077),
.Y(n_2415)
);

OAI222xp33_ASAP7_75t_L g2416 ( 
.A1(n_2338),
.A2(n_2207),
.B1(n_2068),
.B2(n_2077),
.C1(n_2141),
.C2(n_2163),
.Y(n_2416)
);

AOI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_2298),
.A2(n_1819),
.B1(n_1961),
.B2(n_2238),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2319),
.B(n_2236),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2345),
.A2(n_1819),
.B1(n_2119),
.B2(n_2151),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2373),
.Y(n_2420)
);

AOI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_2256),
.A2(n_2024),
.B1(n_2157),
.B2(n_2220),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2299),
.A2(n_2217),
.B1(n_2076),
.B2(n_2148),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2257),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2335),
.B(n_2243),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2269),
.B(n_2220),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2266),
.Y(n_2426)
);

BUFx2_ASAP7_75t_L g2427 ( 
.A(n_2372),
.Y(n_2427)
);

NAND3xp33_ASAP7_75t_L g2428 ( 
.A(n_2366),
.B(n_1801),
.C(n_1921),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_2305),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2281),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2277),
.A2(n_2233),
.B1(n_1971),
.B2(n_1964),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2354),
.B(n_2120),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2321),
.A2(n_2268),
.B1(n_2304),
.B2(n_2323),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_SL g2434 ( 
.A(n_2262),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2324),
.A2(n_2199),
.B1(n_1826),
.B2(n_1812),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2376),
.B(n_2120),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2294),
.A2(n_2217),
.B1(n_2106),
.B2(n_2112),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2266),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_SL g2439 ( 
.A1(n_2339),
.A2(n_2059),
.B(n_2044),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2296),
.A2(n_2281),
.B1(n_2280),
.B2(n_2343),
.Y(n_2440)
);

AOI222xp33_ASAP7_75t_L g2441 ( 
.A1(n_2260),
.A2(n_1918),
.B1(n_1971),
.B2(n_1922),
.C1(n_2053),
.C2(n_2031),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2343),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2369),
.A2(n_2106),
.B1(n_2084),
.B2(n_2112),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2362),
.A2(n_2364),
.B1(n_2365),
.B2(n_2307),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2303),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2358),
.A2(n_2199),
.B1(n_2208),
.B2(n_2110),
.Y(n_2446)
);

AOI22xp33_ASAP7_75t_SL g2447 ( 
.A1(n_2317),
.A2(n_2141),
.B1(n_2163),
.B2(n_2114),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2273),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2358),
.A2(n_2208),
.B1(n_2110),
.B2(n_2044),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2375),
.A2(n_2271),
.B1(n_2300),
.B2(n_2348),
.Y(n_2450)
);

AOI22xp33_ASAP7_75t_L g2451 ( 
.A1(n_2360),
.A2(n_2247),
.B1(n_1976),
.B2(n_1892),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2309),
.Y(n_2452)
);

OAI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2317),
.A2(n_2340),
.B1(n_2342),
.B2(n_2360),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2340),
.A2(n_2084),
.B1(n_2252),
.B2(n_2114),
.Y(n_2454)
);

INVx5_ASAP7_75t_SL g2455 ( 
.A(n_2272),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2377),
.Y(n_2456)
);

AOI22xp33_ASAP7_75t_L g2457 ( 
.A1(n_2311),
.A2(n_2247),
.B1(n_2230),
.B2(n_2228),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2310),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2351),
.Y(n_2459)
);

AOI222xp33_ASAP7_75t_L g2460 ( 
.A1(n_2260),
.A2(n_1864),
.B1(n_2109),
.B2(n_2121),
.C1(n_2146),
.C2(n_2162),
.Y(n_2460)
);

INVx1_ASAP7_75t_SL g2461 ( 
.A(n_2305),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2370),
.A2(n_2155),
.B1(n_2170),
.B2(n_2162),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_2263),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2349),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2379),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2270),
.Y(n_2466)
);

BUFx4f_ASAP7_75t_SL g2467 ( 
.A(n_2286),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2292),
.A2(n_2161),
.B1(n_2156),
.B2(n_2160),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2301),
.A2(n_2161),
.B1(n_2156),
.B2(n_2160),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2393),
.A2(n_2355),
.B1(n_2342),
.B2(n_2380),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2423),
.B(n_2346),
.Y(n_2471)
);

AOI22xp33_ASAP7_75t_SL g2472 ( 
.A1(n_2444),
.A2(n_2396),
.B1(n_2450),
.B2(n_2453),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2382),
.A2(n_2349),
.B1(n_2267),
.B2(n_2359),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2393),
.A2(n_1976),
.B1(n_2001),
.B2(n_2320),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2413),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2441),
.A2(n_2001),
.B1(n_2320),
.B2(n_2241),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_SL g2477 ( 
.A1(n_2443),
.A2(n_2275),
.B1(n_2258),
.B2(n_2302),
.Y(n_2477)
);

NAND3xp33_ASAP7_75t_L g2478 ( 
.A(n_2414),
.B(n_1796),
.C(n_2080),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2409),
.A2(n_1797),
.B(n_1791),
.Y(n_2479)
);

AOI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2382),
.A2(n_2241),
.B1(n_2218),
.B2(n_2219),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2421),
.A2(n_2325),
.B1(n_2371),
.B2(n_2293),
.Y(n_2481)
);

AOI22xp33_ASAP7_75t_L g2482 ( 
.A1(n_2433),
.A2(n_2212),
.B1(n_2242),
.B2(n_2198),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2433),
.A2(n_2242),
.B1(n_2213),
.B2(n_2318),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2397),
.B(n_2290),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2432),
.B(n_2125),
.Y(n_2485)
);

OAI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2421),
.A2(n_2325),
.B1(n_1782),
.B2(n_1816),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2428),
.A2(n_1823),
.B(n_2147),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2395),
.A2(n_2318),
.B1(n_2222),
.B2(n_2363),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2384),
.B(n_2125),
.Y(n_2489)
);

AOI22xp33_ASAP7_75t_L g2490 ( 
.A1(n_2417),
.A2(n_2222),
.B1(n_2278),
.B2(n_1981),
.Y(n_2490)
);

OAI222xp33_ASAP7_75t_L g2491 ( 
.A1(n_2389),
.A2(n_2391),
.B1(n_2394),
.B2(n_2415),
.C1(n_2383),
.C2(n_2468),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2413),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2426),
.B(n_2240),
.Y(n_2493)
);

AOI22xp33_ASAP7_75t_L g2494 ( 
.A1(n_2417),
.A2(n_1981),
.B1(n_2176),
.B2(n_2175),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_2464),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2438),
.B(n_2290),
.Y(n_2496)
);

OAI221xp5_ASAP7_75t_SL g2497 ( 
.A1(n_2383),
.A2(n_1984),
.B1(n_2308),
.B2(n_2026),
.C(n_2201),
.Y(n_2497)
);

OAI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2391),
.A2(n_2104),
.B1(n_2263),
.B2(n_2289),
.Y(n_2498)
);

AOI22xp33_ASAP7_75t_L g2499 ( 
.A1(n_2424),
.A2(n_2175),
.B1(n_2176),
.B2(n_1931),
.Y(n_2499)
);

AOI21xp33_ASAP7_75t_SL g2500 ( 
.A1(n_2460),
.A2(n_2316),
.B(n_2286),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2435),
.A2(n_2390),
.B1(n_2385),
.B2(n_2422),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2442),
.B(n_2290),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2419),
.A2(n_2263),
.B1(n_2289),
.B2(n_2297),
.Y(n_2503)
);

AOI22xp33_ASAP7_75t_L g2504 ( 
.A1(n_2390),
.A2(n_1947),
.B1(n_1931),
.B2(n_2116),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2386),
.B(n_2127),
.Y(n_2505)
);

AOI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_2408),
.A2(n_1947),
.B1(n_2116),
.B2(n_2158),
.Y(n_2506)
);

AOI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_2419),
.A2(n_2289),
.B1(n_2295),
.B2(n_2297),
.Y(n_2507)
);

OAI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2468),
.A2(n_2129),
.B1(n_2139),
.B2(n_2131),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2456),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2387),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2392),
.B(n_2127),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2440),
.A2(n_2158),
.B1(n_2237),
.B2(n_2139),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2410),
.Y(n_2513)
);

NAND2xp33_ASAP7_75t_SL g2514 ( 
.A(n_2434),
.B(n_2254),
.Y(n_2514)
);

OAI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2469),
.A2(n_2133),
.B1(n_2131),
.B2(n_2130),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2449),
.A2(n_2237),
.B1(n_2133),
.B2(n_2129),
.Y(n_2516)
);

NOR3xp33_ASAP7_75t_L g2517 ( 
.A(n_2439),
.B(n_2255),
.C(n_2259),
.Y(n_2517)
);

OAI221xp5_ASAP7_75t_SL g2518 ( 
.A1(n_2431),
.A2(n_2130),
.B1(n_1722),
.B2(n_1752),
.C(n_2142),
.Y(n_2518)
);

OAI222xp33_ASAP7_75t_L g2519 ( 
.A1(n_2415),
.A2(n_2164),
.B1(n_2181),
.B2(n_2079),
.C1(n_2082),
.C2(n_2191),
.Y(n_2519)
);

AOI222xp33_ASAP7_75t_L g2520 ( 
.A1(n_2467),
.A2(n_2327),
.B1(n_2374),
.B2(n_2291),
.C1(n_2295),
.C2(n_2144),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2420),
.B(n_2178),
.Y(n_2521)
);

OAI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2469),
.A2(n_2179),
.B1(n_2231),
.B2(n_2227),
.Y(n_2522)
);

AOI22xp33_ASAP7_75t_L g2523 ( 
.A1(n_2388),
.A2(n_1993),
.B1(n_1990),
.B2(n_1975),
.Y(n_2523)
);

OAI221xp5_ASAP7_75t_L g2524 ( 
.A1(n_2431),
.A2(n_2353),
.B1(n_1916),
.B2(n_1648),
.C(n_1663),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2446),
.A2(n_1990),
.B1(n_1993),
.B2(n_1924),
.Y(n_2525)
);

NAND3xp33_ASAP7_75t_L g2526 ( 
.A(n_2472),
.B(n_2427),
.C(n_2462),
.Y(n_2526)
);

OAI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_2483),
.A2(n_2462),
.B1(n_2447),
.B2(n_2411),
.Y(n_2527)
);

HB1xp67_ASAP7_75t_L g2528 ( 
.A(n_2495),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2509),
.B(n_2510),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_2478),
.B(n_2403),
.C(n_2407),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2500),
.B(n_2464),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2509),
.B(n_2513),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2514),
.B(n_2467),
.Y(n_2533)
);

AND2x2_ASAP7_75t_SL g2534 ( 
.A(n_2517),
.B(n_2430),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2485),
.B(n_2459),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2475),
.Y(n_2536)
);

AOI221xp5_ASAP7_75t_L g2537 ( 
.A1(n_2491),
.A2(n_2425),
.B1(n_2398),
.B2(n_2418),
.C(n_2416),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2475),
.B(n_2465),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2481),
.B(n_2429),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_L g2540 ( 
.A(n_2470),
.B(n_2457),
.C(n_2451),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2496),
.B(n_2461),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2496),
.B(n_2448),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2495),
.B(n_2401),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2492),
.B(n_2402),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2477),
.B(n_2412),
.Y(n_2545)
);

NAND3xp33_ASAP7_75t_L g2546 ( 
.A(n_2514),
.B(n_2457),
.C(n_2445),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2501),
.A2(n_2434),
.B1(n_2404),
.B2(n_2405),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2476),
.A2(n_2482),
.B1(n_2518),
.B2(n_2490),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2497),
.A2(n_2455),
.B1(n_2430),
.B2(n_2454),
.Y(n_2549)
);

OAI221xp5_ASAP7_75t_L g2550 ( 
.A1(n_2488),
.A2(n_2399),
.B1(n_2463),
.B2(n_2400),
.C(n_2406),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2484),
.B(n_2452),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2502),
.B(n_2458),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2503),
.A2(n_2455),
.B1(n_2437),
.B2(n_2436),
.Y(n_2553)
);

OAI21xp5_ASAP7_75t_SL g2554 ( 
.A1(n_2520),
.A2(n_2455),
.B(n_1676),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_2484),
.B(n_2374),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2502),
.B(n_2312),
.Y(n_2556)
);

INVxp67_ASAP7_75t_L g2557 ( 
.A(n_2528),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2526),
.A2(n_2474),
.B1(n_2473),
.B2(n_2523),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2536),
.B(n_2492),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2541),
.B(n_2542),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2529),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2552),
.B(n_2471),
.Y(n_2562)
);

NOR3xp33_ASAP7_75t_L g2563 ( 
.A(n_2533),
.B(n_2524),
.C(n_2479),
.Y(n_2563)
);

OR2x2_ASAP7_75t_SL g2564 ( 
.A(n_2530),
.B(n_2489),
.Y(n_2564)
);

AO21x2_ASAP7_75t_L g2565 ( 
.A1(n_2551),
.A2(n_2487),
.B(n_2505),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2556),
.B(n_2471),
.Y(n_2566)
);

OR2x2_ASAP7_75t_L g2567 ( 
.A(n_2532),
.B(n_2493),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2544),
.B(n_2493),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2538),
.B(n_2535),
.Y(n_2569)
);

AOI221xp5_ASAP7_75t_L g2570 ( 
.A1(n_2537),
.A2(n_2515),
.B1(n_2508),
.B2(n_2498),
.C(n_2511),
.Y(n_2570)
);

AOI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2548),
.A2(n_2521),
.B1(n_2486),
.B2(n_2506),
.C(n_2519),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2539),
.B(n_2543),
.Y(n_2572)
);

OA211x2_ASAP7_75t_L g2573 ( 
.A1(n_2545),
.A2(n_2494),
.B(n_2504),
.C(n_2516),
.Y(n_2573)
);

NAND3xp33_ASAP7_75t_L g2574 ( 
.A(n_2545),
.B(n_2507),
.C(n_2512),
.Y(n_2574)
);

NAND3xp33_ASAP7_75t_L g2575 ( 
.A(n_2547),
.B(n_2480),
.C(n_2499),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2543),
.Y(n_2576)
);

AOI22xp33_ASAP7_75t_L g2577 ( 
.A1(n_2534),
.A2(n_2525),
.B1(n_2522),
.B2(n_2211),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_R g2578 ( 
.A(n_2534),
.B(n_2466),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2547),
.B(n_1786),
.C(n_2368),
.Y(n_2579)
);

NOR3xp33_ASAP7_75t_L g2580 ( 
.A(n_2554),
.B(n_2540),
.C(n_2531),
.Y(n_2580)
);

NOR2x1_ASAP7_75t_L g2581 ( 
.A(n_2555),
.B(n_2549),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2539),
.B(n_2312),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2560),
.Y(n_2583)
);

XOR2x2_ASAP7_75t_L g2584 ( 
.A(n_2580),
.B(n_2550),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2561),
.B(n_2551),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2569),
.B(n_2546),
.Y(n_2586)
);

XOR2x2_ASAP7_75t_L g2587 ( 
.A(n_2580),
.B(n_2553),
.Y(n_2587)
);

INVx2_ASAP7_75t_SL g2588 ( 
.A(n_2562),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2559),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2557),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2576),
.B(n_2527),
.Y(n_2591)
);

NAND4xp75_ASAP7_75t_L g2592 ( 
.A(n_2573),
.B(n_1946),
.C(n_1987),
.D(n_1957),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2566),
.B(n_2312),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2572),
.B(n_2557),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2567),
.Y(n_2595)
);

NAND4xp75_ASAP7_75t_L g2596 ( 
.A(n_2581),
.B(n_1962),
.C(n_1982),
.D(n_1958),
.Y(n_2596)
);

NOR3xp33_ASAP7_75t_L g2597 ( 
.A(n_2571),
.B(n_2006),
.C(n_2021),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2565),
.B(n_2062),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2568),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2582),
.Y(n_2600)
);

XNOR2xp5_ASAP7_75t_L g2601 ( 
.A(n_2564),
.B(n_1757),
.Y(n_2601)
);

XNOR2xp5_ASAP7_75t_L g2602 ( 
.A(n_2575),
.B(n_1743),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2565),
.B(n_2062),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2574),
.Y(n_2604)
);

INVx4_ASAP7_75t_L g2605 ( 
.A(n_2578),
.Y(n_2605)
);

NAND4xp75_ASAP7_75t_L g2606 ( 
.A(n_2570),
.B(n_2205),
.C(n_2190),
.D(n_2187),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2585),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2594),
.B(n_2578),
.Y(n_2608)
);

XOR2x2_ASAP7_75t_L g2609 ( 
.A(n_2584),
.B(n_2563),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2590),
.Y(n_2610)
);

XNOR2x2_ASAP7_75t_L g2611 ( 
.A(n_2587),
.B(n_2596),
.Y(n_2611)
);

XOR2x2_ASAP7_75t_L g2612 ( 
.A(n_2605),
.B(n_2563),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2583),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2585),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2605),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2589),
.Y(n_2616)
);

AO22x2_ASAP7_75t_L g2617 ( 
.A1(n_2604),
.A2(n_2579),
.B1(n_2577),
.B2(n_2558),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2599),
.Y(n_2618)
);

BUFx2_ASAP7_75t_L g2619 ( 
.A(n_2588),
.Y(n_2619)
);

AOI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2612),
.A2(n_2597),
.B1(n_2591),
.B2(n_2592),
.Y(n_2620)
);

INVxp67_ASAP7_75t_L g2621 ( 
.A(n_2612),
.Y(n_2621)
);

OA22x2_ASAP7_75t_L g2622 ( 
.A1(n_2615),
.A2(n_2591),
.B1(n_2601),
.B2(n_2602),
.Y(n_2622)
);

CKINVDCx14_ASAP7_75t_R g2623 ( 
.A(n_2609),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2619),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2616),
.Y(n_2625)
);

OAI22x1_ASAP7_75t_L g2626 ( 
.A1(n_2608),
.A2(n_2611),
.B1(n_2613),
.B2(n_2609),
.Y(n_2626)
);

OA22x2_ASAP7_75t_L g2627 ( 
.A1(n_2611),
.A2(n_2595),
.B1(n_2600),
.B2(n_2593),
.Y(n_2627)
);

XOR2x2_ASAP7_75t_L g2628 ( 
.A(n_2618),
.B(n_2606),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2613),
.Y(n_2629)
);

AOI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2617),
.A2(n_2597),
.B1(n_2607),
.B2(n_2614),
.Y(n_2630)
);

NOR2x1_ASAP7_75t_L g2631 ( 
.A(n_2610),
.B(n_2586),
.Y(n_2631)
);

XOR2x2_ASAP7_75t_L g2632 ( 
.A(n_2617),
.B(n_2558),
.Y(n_2632)
);

OA22x2_ASAP7_75t_L g2633 ( 
.A1(n_2617),
.A2(n_2603),
.B1(n_2598),
.B2(n_2577),
.Y(n_2633)
);

OAI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2610),
.A2(n_2603),
.B1(n_2598),
.B2(n_2353),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_SL g2635 ( 
.A1(n_2615),
.A2(n_2231),
.B1(n_2221),
.B2(n_2227),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2625),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_SL g2637 ( 
.A(n_2626),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2632),
.A2(n_1998),
.B1(n_2368),
.B2(n_2331),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2625),
.Y(n_2639)
);

OAI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2627),
.A2(n_2368),
.B1(n_2367),
.B2(n_2331),
.Y(n_2640)
);

AOI22x1_ASAP7_75t_L g2641 ( 
.A1(n_2621),
.A2(n_1860),
.B1(n_1804),
.B2(n_1798),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2624),
.Y(n_2642)
);

INVx2_ASAP7_75t_SL g2643 ( 
.A(n_2629),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2631),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2635),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2630),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2620),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2623),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_L g2649 ( 
.A(n_2634),
.B(n_2179),
.Y(n_2649)
);

INVxp67_ASAP7_75t_L g2650 ( 
.A(n_2648),
.Y(n_2650)
);

AOI32xp33_ASAP7_75t_L g2651 ( 
.A1(n_2647),
.A2(n_2645),
.A3(n_2646),
.B1(n_2648),
.B2(n_2644),
.Y(n_2651)
);

OA22x2_ASAP7_75t_L g2652 ( 
.A1(n_2637),
.A2(n_2622),
.B1(n_2633),
.B2(n_2628),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2642),
.Y(n_2653)
);

OAI221xp5_ASAP7_75t_L g2654 ( 
.A1(n_2638),
.A2(n_2025),
.B1(n_2227),
.B2(n_2231),
.C(n_2221),
.Y(n_2654)
);

AOI22x1_ASAP7_75t_L g2655 ( 
.A1(n_2637),
.A2(n_1997),
.B1(n_2021),
.B2(n_2006),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2643),
.A2(n_1924),
.B1(n_2331),
.B2(n_2314),
.Y(n_2656)
);

AOI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2640),
.A2(n_1924),
.B1(n_2314),
.B2(n_2367),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2636),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2649),
.A2(n_2367),
.B1(n_2314),
.B2(n_2179),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2639),
.A2(n_1997),
.B1(n_2245),
.B2(n_2180),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2641),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2637),
.A2(n_1798),
.B1(n_1804),
.B2(n_1860),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2650),
.Y(n_2663)
);

INVxp67_ASAP7_75t_SL g2664 ( 
.A(n_2661),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2653),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2658),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2660),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2652),
.A2(n_1743),
.B1(n_1740),
.B2(n_2221),
.Y(n_2668)
);

OAI22x1_ASAP7_75t_L g2669 ( 
.A1(n_2655),
.A2(n_2651),
.B1(n_2657),
.B2(n_2656),
.Y(n_2669)
);

AOI221xp5_ASAP7_75t_L g2670 ( 
.A1(n_2654),
.A2(n_1740),
.B1(n_2022),
.B2(n_2015),
.C(n_2004),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2662),
.A2(n_1980),
.B1(n_1885),
.B2(n_1884),
.Y(n_2671)
);

AOI221xp5_ASAP7_75t_L g2672 ( 
.A1(n_2659),
.A2(n_1492),
.B1(n_1457),
.B2(n_1885),
.C(n_1884),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2650),
.Y(n_2673)
);

AOI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2652),
.A2(n_1885),
.B1(n_1884),
.B2(n_1818),
.Y(n_2674)
);

OAI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2652),
.A2(n_2249),
.B1(n_2232),
.B2(n_2204),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2650),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2673),
.A2(n_2232),
.B1(n_2204),
.B2(n_2203),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2676),
.Y(n_2678)
);

NOR2x1_ASAP7_75t_L g2679 ( 
.A(n_2663),
.B(n_1777),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2664),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2667),
.A2(n_2177),
.B1(n_2172),
.B2(n_2204),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2675),
.B(n_2152),
.Y(n_2682)
);

NOR3xp33_ASAP7_75t_L g2683 ( 
.A(n_2675),
.B(n_1818),
.C(n_1777),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2666),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2684),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2678),
.A2(n_2669),
.B1(n_2668),
.B2(n_2674),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2680),
.A2(n_2665),
.B1(n_2671),
.B2(n_2672),
.Y(n_2687)
);

BUFx3_ASAP7_75t_L g2688 ( 
.A(n_2677),
.Y(n_2688)
);

AOI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2681),
.A2(n_2670),
.B1(n_2232),
.B2(n_2203),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2685),
.Y(n_2690)
);

BUFx2_ASAP7_75t_L g2691 ( 
.A(n_2688),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2691),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2690),
.A2(n_2686),
.B1(n_2687),
.B2(n_2679),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2692),
.Y(n_2694)
);

OA22x2_ASAP7_75t_L g2695 ( 
.A1(n_2693),
.A2(n_2689),
.B1(n_2682),
.B2(n_2683),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2694),
.Y(n_2696)
);

INVxp67_ASAP7_75t_SL g2697 ( 
.A(n_2695),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2697),
.A2(n_2203),
.B1(n_2202),
.B2(n_2183),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2698),
.Y(n_2699)
);

OAI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2699),
.A2(n_2696),
.B1(n_2202),
.B2(n_2183),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2700),
.Y(n_2701)
);

AOI221xp5_ASAP7_75t_L g2702 ( 
.A1(n_2701),
.A2(n_1811),
.B1(n_1748),
.B2(n_2172),
.C(n_2169),
.Y(n_2702)
);

AOI211xp5_ASAP7_75t_L g2703 ( 
.A1(n_2702),
.A2(n_1699),
.B(n_2202),
.C(n_2183),
.Y(n_2703)
);


endmodule