module fake_netlist_1_7032_n_260 (n_20, n_2, n_38, n_44, n_36, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_29, n_43, n_7, n_40, n_27, n_39, n_260);
input n_20;
input n_2;
input n_38;
input n_44;
input n_36;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_260;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_57;
wire n_88;
wire n_52;
wire n_244;
wire n_50;
wire n_102;
wire n_73;
wire n_49;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_80;
wire n_167;
wire n_107;
wire n_158;
wire n_60;
wire n_114;
wire n_121;
wire n_94;
wire n_65;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_87;
wire n_180;
wire n_104;
wire n_160;
wire n_98;
wire n_74;
wire n_206;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_45;
wire n_85;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_47;
wire n_215;
wire n_116;
wire n_91;
wire n_108;
wire n_155;
wire n_209;
wire n_217;
wire n_139;
wire n_229;
wire n_230;
wire n_198;
wire n_169;
wire n_193;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_95;
wire n_124;
wire n_156;
wire n_238;
wire n_128;
wire n_120;
wire n_129;
wire n_70;
wire n_90;
wire n_71;
wire n_63;
wire n_56;
wire n_135;
wire n_188;
wire n_78;
wire n_247;
wire n_197;
wire n_201;
wire n_242;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_79;
wire n_210;
wire n_202;
wire n_64;
wire n_142;
wire n_184;
wire n_245;
wire n_191;
wire n_232;
wire n_200;
wire n_46;
wire n_208;
wire n_211;
wire n_58;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_84;
wire n_131;
wire n_112;
wire n_55;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_166;
wire n_162;
wire n_186;
wire n_75;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_231;
wire n_72;
wire n_136;
wire n_76;
wire n_89;
wire n_176;
wire n_68;
wire n_144;
wire n_53;
wire n_183;
wire n_256;
wire n_67;
wire n_77;
wire n_216;
wire n_147;
wire n_199;
wire n_54;
wire n_148;
wire n_123;
wire n_83;
wire n_172;
wire n_48;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_59;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_66;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_82;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_246;
wire n_153;
wire n_61;
wire n_259;
wire n_99;
wire n_109;
wire n_93;
wire n_132;
wire n_151;
wire n_51;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_96;
wire n_225;
INVx1_ASAP7_75t_L g45 ( .A(n_17), .Y(n_45) );
XOR2xp5_ASAP7_75t_L g46 ( .A(n_41), .B(n_31), .Y(n_46) );
INVxp33_ASAP7_75t_L g47 ( .A(n_4), .Y(n_47) );
INVx1_ASAP7_75t_L g48 ( .A(n_37), .Y(n_48) );
INVx1_ASAP7_75t_L g49 ( .A(n_33), .Y(n_49) );
INVx1_ASAP7_75t_L g50 ( .A(n_24), .Y(n_50) );
CKINVDCx5p33_ASAP7_75t_R g51 ( .A(n_28), .Y(n_51) );
CKINVDCx5p33_ASAP7_75t_R g52 ( .A(n_16), .Y(n_52) );
INVx1_ASAP7_75t_L g53 ( .A(n_30), .Y(n_53) );
INVx1_ASAP7_75t_L g54 ( .A(n_34), .Y(n_54) );
INVx1_ASAP7_75t_L g55 ( .A(n_21), .Y(n_55) );
INVx1_ASAP7_75t_L g56 ( .A(n_36), .Y(n_56) );
INVx1_ASAP7_75t_L g57 ( .A(n_11), .Y(n_57) );
INVx2_ASAP7_75t_L g58 ( .A(n_27), .Y(n_58) );
INVx1_ASAP7_75t_L g59 ( .A(n_29), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_22), .Y(n_60) );
BUFx3_ASAP7_75t_L g61 ( .A(n_23), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_6), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_13), .Y(n_63) );
INVx3_ASAP7_75t_L g64 ( .A(n_10), .Y(n_64) );
BUFx3_ASAP7_75t_L g65 ( .A(n_15), .Y(n_65) );
BUFx2_ASAP7_75t_SL g66 ( .A(n_26), .Y(n_66) );
BUFx6f_ASAP7_75t_L g67 ( .A(n_32), .Y(n_67) );
CKINVDCx5p33_ASAP7_75t_R g68 ( .A(n_25), .Y(n_68) );
BUFx6f_ASAP7_75t_L g69 ( .A(n_43), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_7), .Y(n_70) );
INVx2_ASAP7_75t_L g71 ( .A(n_40), .Y(n_71) );
BUFx3_ASAP7_75t_L g72 ( .A(n_14), .Y(n_72) );
INVxp33_ASAP7_75t_L g73 ( .A(n_5), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_9), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_8), .Y(n_75) );
HB1xp67_ASAP7_75t_L g76 ( .A(n_42), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_35), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_64), .Y(n_82) );
AND2x2_ASAP7_75t_SL g83 ( .A(n_76), .B(n_44), .Y(n_83) );
BUFx8_ASAP7_75t_L g84 ( .A(n_67), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_48), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_48), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_67), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_45), .B(n_0), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_49), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx6_ASAP7_75t_L g93 ( .A(n_61), .Y(n_93) );
AND2x2_ASAP7_75t_L g94 ( .A(n_47), .B(n_1), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_50), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_45), .B(n_2), .Y(n_96) );
AND2x2_ASAP7_75t_L g97 ( .A(n_73), .B(n_3), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_50), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_79), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_86), .B(n_58), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_84), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_79), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_81), .B(n_51), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_87), .B(n_71), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_80), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_79), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_82), .B(n_72), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_90), .B(n_77), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
AO22x2_ASAP7_75t_L g112 ( .A1(n_83), .A2(n_46), .B1(n_54), .B2(n_53), .Y(n_112) );
AO22x2_ASAP7_75t_L g113 ( .A1(n_83), .A2(n_46), .B1(n_55), .B2(n_54), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_94), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_85), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_88), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_94), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_97), .B(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_95), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_102), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_115), .A2(n_97), .B1(n_99), .B2(n_98), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_119), .A2(n_96), .B(n_89), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_104), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_116), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_116), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_118), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_118), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_121), .Y(n_132) );
OR2x6_ASAP7_75t_L g133 ( .A(n_112), .B(n_66), .Y(n_133) );
OR2x2_ASAP7_75t_L g134 ( .A(n_119), .B(n_52), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_120), .B(n_57), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_115), .B(n_70), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_106), .B(n_55), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_105), .B(n_68), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_110), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_114), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_113), .B(n_70), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_114), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_113), .B(n_75), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_132), .A2(n_59), .B(n_56), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_144), .A2(n_74), .B1(n_62), .B2(n_63), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_126), .A2(n_111), .B(n_103), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_130), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_136), .B(n_139), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
NOR2x1_ASAP7_75t_SL g167 ( .A(n_133), .B(n_60), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_144), .B1(n_147), .B2(n_146), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_162), .A2(n_124), .B1(n_123), .B2(n_138), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_172), .B(n_137), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_165), .B(n_141), .Y(n_177) );
INVx5_ASAP7_75t_L g178 ( .A(n_171), .Y(n_178) );
INVxp67_ASAP7_75t_SL g179 ( .A(n_170), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_171), .B(n_78), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_156), .A2(n_117), .B(n_100), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_159), .A2(n_91), .B(n_92), .C(n_108), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_163), .B1(n_168), .B2(n_150), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_173), .A2(n_154), .B1(n_155), .B2(n_153), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_177), .B(n_148), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_179), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_181), .A2(n_167), .B(n_151), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_185), .A2(n_169), .B1(n_166), .B2(n_160), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_185), .A2(n_169), .B1(n_166), .B2(n_160), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_175), .A2(n_158), .B1(n_152), .B2(n_151), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_174), .B(n_149), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_178), .B(n_12), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_180), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_183), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_176), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_182), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_188), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_187), .B(n_184), .Y(n_201) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_192), .A2(n_38), .B(n_39), .Y(n_202) );
AO31x2_ASAP7_75t_L g203 ( .A1(n_190), .A2(n_191), .A3(n_186), .B(n_189), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_197), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_197), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_193), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_198), .B(n_194), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_196), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_196), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_187), .B(n_199), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_211), .B(n_201), .Y(n_212) );
AND2x4_ASAP7_75t_SL g213 ( .A(n_207), .B(n_200), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_206), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_204), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_205), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_205), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_208), .B(n_210), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_209), .B(n_210), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_202), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_203), .B(n_211), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_222), .B(n_212), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_213), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_214), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_216), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_215), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_217), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_219), .B(n_220), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_224), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_225), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_223), .B(n_221), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_226), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_227), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_229), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_229), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_230), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_232), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_234), .B(n_231), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_235), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_233), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_236), .B(n_228), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_241), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_243), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_245), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_246), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_248), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_247), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_249), .Y(n_251) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_250), .B(n_242), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_251), .B(n_240), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_252), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_253), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_254), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_256), .B(n_244), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_255), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_258), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_259), .A2(n_257), .B1(n_237), .B2(n_238), .C(n_239), .Y(n_260) );
endmodule