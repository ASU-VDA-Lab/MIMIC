module fake_jpeg_18718_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_52),
.B1(n_51),
.B2(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_53),
.B1(n_54),
.B2(n_6),
.Y(n_84)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_76),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_47),
.B1(n_40),
.B2(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_71),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_56),
.B1(n_39),
.B2(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_39),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_55),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_50),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_53),
.B1(n_41),
.B2(n_46),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_7),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_100),
.B1(n_19),
.B2(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_99),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_9),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_24),
.B(n_25),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_12),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_31),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_27),
.C(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_97),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_93),
.B1(n_94),
.B2(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_109),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_92),
.A3(n_107),
.B1(n_112),
.B2(n_110),
.C1(n_100),
.C2(n_38),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_33),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_34),
.Y(n_121)
);


endmodule