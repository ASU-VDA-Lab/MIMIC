module real_jpeg_6197_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_0),
.A2(n_40),
.B1(n_200),
.B2(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_0),
.B(n_292),
.C(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_0),
.B(n_121),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_0),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_0),
.B(n_178),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_0),
.B(n_358),
.Y(n_357)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_2),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_2),
.A2(n_134),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_2),
.A2(n_58),
.B1(n_134),
.B2(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_2),
.A2(n_134),
.B1(n_182),
.B2(n_202),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_3),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_3),
.A2(n_135),
.B1(n_176),
.B2(n_223),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_3),
.A2(n_176),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_5),
.A2(n_62),
.B1(n_175),
.B2(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_7),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_7),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_73),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_12),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_12),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_12),
.A2(n_96),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_12),
.A2(n_96),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_12),
.A2(n_96),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_28),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_13),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_80),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_13),
.A2(n_80),
.B1(n_181),
.B2(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_13),
.A2(n_80),
.B1(n_302),
.B2(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_14),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_14),
.Y(n_157)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_14),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_14),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_15),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_16),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_16),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_251),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_250),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_213),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_21),
.B(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_144),
.C(n_195),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_22),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_23),
.B(n_77),
.C(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_24),
.A2(n_45),
.B1(n_46),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_24),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.A3(n_30),
.B1(n_33),
.B2(n_39),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_27),
.Y(n_360)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_32),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_39),
.A2(n_40),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_40),
.B(n_83),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_40),
.A2(n_47),
.B(n_299),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g354 ( 
.A1(n_40),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B1(n_63),
.B2(n_66),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_47),
.A2(n_187),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_47),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_48),
.A2(n_64),
.B1(n_67),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_48),
.A2(n_55),
.B1(n_64),
.B2(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_48),
.B(n_301),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_48),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_51),
.Y(n_304)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_53),
.Y(n_165)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_53),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_60),
.Y(n_247)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_61),
.Y(n_330)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_68),
.Y(n_245)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_70),
.Y(n_194)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_71),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_72),
.Y(n_191)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_75),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_106),
.B2(n_107),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_94),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_79),
.A2(n_83),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_84),
.B(n_95),
.Y(n_208)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_101),
.A2(n_205),
.B(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_101),
.Y(n_227)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_104),
.Y(n_229)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_130),
.B(n_137),
.Y(n_107)
);

AOI22x1_ASAP7_75t_L g219 ( 
.A1(n_108),
.A2(n_121),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_108),
.B(n_220),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_108),
.A2(n_137),
.B(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_109),
.A2(n_131),
.B1(n_143),
.B2(n_210),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_110)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_111),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_118),
.Y(n_370)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_135),
.A2(n_357),
.A3(n_366),
.B1(n_369),
.B2(n_371),
.Y(n_365)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_143),
.A2(n_210),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_144),
.A2(n_145),
.B1(n_195),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_185),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_146),
.B(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_171),
.B1(n_177),
.B2(n_179),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_147),
.A2(n_281),
.B(n_285),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_147),
.A2(n_177),
.B1(n_308),
.B2(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_147),
.A2(n_285),
.B(n_351),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_148),
.A2(n_178),
.B1(n_180),
.B2(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_160),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_152),
.B1(n_155),
.B2(n_158),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_159),
.Y(n_368)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_160),
.A2(n_197),
.B(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_177),
.B(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_174),
.Y(n_311)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_178),
.B(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_193),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.C(n_209),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_196),
.B(n_209),
.Y(n_256)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_203),
.A2(n_204),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_233),
.B1(n_248),
.B2(n_249),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_238),
.B(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_274),
.B(n_391),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_254),
.B(n_271),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_261),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_255),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_261),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.C(n_270),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_262),
.B(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_264),
.B(n_270),
.Y(n_382)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_385),
.B(n_390),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_374),
.B(n_384),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_345),
.B(n_373),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_314),
.B(n_344),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_294),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_294),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_280),
.A2(n_286),
.B1(n_287),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_305),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_306),
.C(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx11_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_336),
.B(n_343),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_325),
.B(n_335),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_334),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_334),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_331),
.B(n_333),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_363),
.B(n_364),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_341),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_347),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_361),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_352),
.C(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

INVx6_ASAP7_75t_SL g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_365),
.Y(n_380)
);

INVx5_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_375),
.B(n_376),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_383),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_380),
.C(n_383),
.Y(n_386)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_386),
.B(n_387),
.Y(n_390)
);


endmodule