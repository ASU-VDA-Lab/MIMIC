module real_jpeg_33632_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_0),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_1),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_82),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_82),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_448),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_2),
.B(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_46),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_6),
.A2(n_46),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_6),
.A2(n_46),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_6),
.B(n_258),
.Y(n_257)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_6),
.A2(n_282),
.A3(n_284),
.B1(n_286),
.B2(n_292),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_6),
.B(n_92),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_6),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_6),
.B(n_137),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_10),
.A2(n_106),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_10),
.A2(n_106),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

AOI22x1_ASAP7_75t_L g33 ( 
.A1(n_12),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_33)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_12),
.A2(n_41),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_12),
.A2(n_41),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_13),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_204),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_202),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_183),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_18),
.B(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.C(n_147),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_19),
.A2(n_125),
.B1(n_126),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_19),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_58),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_20),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_20),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_21),
.Y(n_219)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_22),
.B(n_212),
.C(n_215),
.Y(n_396)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g388 ( 
.A1(n_23),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_23),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B(n_42),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_24),
.B(n_182),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_24),
.A2(n_33),
.B1(n_182),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_50),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_25),
.Y(n_258)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_41),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_41),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_43),
.B(n_181),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g192 ( 
.A(n_43),
.Y(n_192)
);

OAI21x1_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_46),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_46),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_46),
.B(n_330),
.Y(n_329)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_47),
.A2(n_223),
.A3(n_227),
.B1(n_230),
.B2(n_232),
.Y(n_222)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

AOI22x1_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_54),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_90),
.B2(n_124),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_59),
.B(n_124),
.C(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_60),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_81),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_61),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_73),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_73),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_73),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_65),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_65),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_65),
.Y(n_333)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_68),
.Y(n_328)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_72),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_73),
.B(n_275),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_75),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_78),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_79),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_129),
.B1(n_135),
.B2(n_137),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_84),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_94),
.B1(n_97),
.B2(n_101),
.Y(n_93)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_88),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_103),
.B(n_110),
.Y(n_90)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_91),
.A2(n_103),
.B1(n_195),
.B2(n_201),
.Y(n_194)
);

AOI21x1_ASAP7_75t_L g390 ( 
.A1(n_91),
.A2(n_139),
.B(n_201),
.Y(n_390)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_92),
.B(n_141),
.Y(n_216)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_111),
.B(n_115),
.Y(n_217)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_121),
.Y(n_291)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_127),
.A2(n_128),
.B(n_138),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_138),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_137),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g273 ( 
.A1(n_135),
.A2(n_137),
.B1(n_213),
.B2(n_274),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_138),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_138),
.A2(n_255),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_138),
.B(n_189),
.C(n_371),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g394 ( 
.A1(n_138),
.A2(n_190),
.B1(n_191),
.B2(n_255),
.Y(n_394)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_147),
.B(n_441),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_158),
.B(n_179),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_148),
.B(n_418),
.Y(n_417)
);

AOI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_157),
.B(n_158),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_149),
.B(n_157),
.Y(n_410)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_151),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_158),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_158),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_158),
.A2(n_179),
.B1(n_180),
.B2(n_411),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_159),
.Y(n_376)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_165),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_166),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_167),
.B(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

OAI22x1_ASAP7_75t_L g375 ( 
.A1(n_168),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_375)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_238),
.B1(n_244),
.B2(n_247),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_169),
.B(n_247),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_175),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_189),
.B(n_215),
.C(n_414),
.Y(n_421)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_190),
.A2(n_191),
.B1(n_214),
.B2(n_215),
.Y(n_415)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_438),
.B(n_446),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_430),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_365),
.B(n_429),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_299),
.B(n_364),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_266),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_209),
.B(n_266),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_210),
.B(n_221),
.C(n_254),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_218),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_214),
.A2(n_215),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_214),
.B(n_352),
.C(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_219),
.B(n_405),
.C(n_406),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_219),
.B(n_405),
.C(n_406),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_254),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_237),
.B1(n_252),
.B2(n_253),
.Y(n_221)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_222),
.B(n_253),
.Y(n_371)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_237),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_237),
.B(n_345),
.Y(n_346)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx4f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_253),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_270)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_314),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_259),
.B(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_339),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.B(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_263),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_265),
.A2(n_378),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.C(n_280),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_267),
.A2(n_268),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_309),
.C(n_310),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_272),
.A2(n_280),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

OAI22x1_ASAP7_75t_L g373 ( 
.A1(n_272),
.A2(n_358),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_310),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

NAND2x1_ASAP7_75t_L g414 ( 
.A(n_273),
.B(n_375),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_298),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_281),
.B(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx4f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_355),
.B(n_363),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_311),
.B(n_354),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_308),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_315),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_385),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_305),
.B(n_385),
.Y(n_395)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_348),
.B(n_353),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_337),
.B(n_347),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_321),
.B1(n_329),
.B2(n_334),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_334),
.B(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_344),
.B(n_346),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_351),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_361),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_357),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_401),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_397),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_392),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_392),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_369),
.B(n_427),
.C(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_383),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_395),
.C(n_396),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_400),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_396),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_399),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_422),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_416),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_416),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.C(n_412),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_413),
.Y(n_425)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_444),
.C(n_445),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_421),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_426),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_437),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B(n_435),
.C(n_436),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_443),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);


endmodule