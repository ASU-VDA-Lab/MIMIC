module fake_netlist_6_2751_n_5199 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5199);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5199;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_1971;
wire n_1781;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4839;
wire n_4489;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_1003;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g701 ( 
.A(n_27),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_541),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_563),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_608),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_80),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_140),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_115),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_65),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_373),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_634),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_33),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_362),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_22),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_348),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_578),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_16),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_573),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_140),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_404),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_186),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_289),
.Y(n_722)
);

CKINVDCx16_ASAP7_75t_R g723 ( 
.A(n_346),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_179),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_239),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_169),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_157),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_525),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_561),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_4),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_173),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_617),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_340),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_49),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_159),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_417),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_604),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_439),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_641),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_575),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_41),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_210),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_65),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_43),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_499),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_482),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_558),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_346),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_453),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_66),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_106),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_227),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_26),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_116),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_594),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_488),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_478),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_669),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_697),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_183),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_255),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_273),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_360),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_264),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_305),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_658),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_404),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_79),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_29),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_288),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_155),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_8),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_524),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_425),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_420),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_373),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_352),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_623),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_362),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_278),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_304),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_338),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_437),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_639),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_110),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_598),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_405),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_306),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_311),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_614),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_385),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_477),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_116),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_252),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_512),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_75),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_228),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_391),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_456),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_67),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_301),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_361),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_424),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_124),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_27),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_470),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_16),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_323),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_53),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_663),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_588),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_466),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_587),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_341),
.Y(n_814)
);

CKINVDCx14_ASAP7_75t_R g815 ( 
.A(n_592),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_530),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_498),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_276),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_382),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_178),
.Y(n_820)
);

INVx4_ASAP7_75t_R g821 ( 
.A(n_223),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_666),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_390),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_48),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_81),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_3),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_400),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_383),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_320),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_219),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_635),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_432),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_386),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_478),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_326),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_423),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_130),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_567),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_409),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_134),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_546),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_170),
.Y(n_842)
);

BUFx5_ASAP7_75t_L g843 ( 
.A(n_609),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_158),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_314),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_191),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_675),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_273),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_531),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

CKINVDCx16_ASAP7_75t_R g851 ( 
.A(n_90),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_472),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_156),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_532),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_616),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_255),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_302),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_566),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_523),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_381),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_671),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_163),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_464),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_393),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_95),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_345),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_215),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_410),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_257),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_75),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_447),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_687),
.Y(n_872)
);

CKINVDCx16_ASAP7_75t_R g873 ( 
.A(n_347),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_501),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_677),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_279),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_418),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_96),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_252),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_653),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_204),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_586),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_427),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_522),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_694),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_228),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_295),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_337),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_552),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_275),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_196),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_263),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_52),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_515),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_309),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_170),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_37),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_434),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_417),
.Y(n_899)
);

CKINVDCx16_ASAP7_75t_R g900 ( 
.A(n_60),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_166),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_50),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_18),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_388),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_155),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_690),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_29),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_245),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_521),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_605),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_349),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_630),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_485),
.Y(n_913)
);

BUFx10_ASAP7_75t_L g914 ( 
.A(n_324),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_254),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_326),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_188),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_60),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_274),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_433),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_188),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_85),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_248),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_337),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_209),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_534),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_646),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_348),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_24),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_432),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_468),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_493),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_674),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_187),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_45),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_490),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_554),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_582),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_518),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_419),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_629),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_52),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_292),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_449),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_130),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_327),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_517),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_284),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_529),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_117),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_20),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_493),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_483),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_323),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_676),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_176),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_41),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_121),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_377),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_504),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_520),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_117),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_44),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_388),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_224),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_371),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_90),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_268),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_33),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_538),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_328),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_123),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_232),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_452),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_428),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_577),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_18),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_46),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_231),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_184),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_540),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_681),
.Y(n_982)
);

BUFx5_ASAP7_75t_L g983 ( 
.A(n_537),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_329),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_332),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_516),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_294),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_699),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_504),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_25),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_679),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_94),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_518),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_501),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_157),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_218),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_209),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_245),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_208),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_590),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_229),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_519),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_13),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_64),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_185),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_294),
.Y(n_1006)
);

BUFx5_ASAP7_75t_L g1007 ( 
.A(n_207),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_250),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_418),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_277),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_500),
.Y(n_1011)
);

BUFx10_ASAP7_75t_L g1012 ( 
.A(n_377),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_644),
.Y(n_1013)
);

BUFx2_ASAP7_75t_SL g1014 ( 
.A(n_249),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_184),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_309),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_437),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_433),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_84),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_665),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_329),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_163),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_290),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_310),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_109),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_673),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_194),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_196),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_661),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_645),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_372),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_169),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_257),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_371),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_112),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_243),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_703),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1007),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1007),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_704),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1007),
.Y(n_1041)
);

INVxp33_ASAP7_75t_L g1042 ( 
.A(n_934),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_715),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1007),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1007),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1007),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_737),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1007),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_729),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1024),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1024),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_740),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_755),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1024),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_786),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_737),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_790),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_758),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_726),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_726),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1036),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1036),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_760),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_813),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_760),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_816),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_761),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_838),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_761),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_723),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_841),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_781),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_849),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_781),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_843),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_763),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_758),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_788),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_851),
.Y(n_1079)
);

CKINVDCx14_ASAP7_75t_R g1080 ( 
.A(n_815),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_872),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_788),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_805),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_843),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_875),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_880),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_805),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_946),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_946),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_837),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_837),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_882),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_837),
.Y(n_1093)
);

BUFx5_ASAP7_75t_L g1094 ( 
.A(n_716),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_837),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_953),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_953),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_721),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_885),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_906),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_910),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_953),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_953),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_964),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_926),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_964),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_843),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_964),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_927),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_758),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_933),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_964),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_701),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_705),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_712),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_714),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_950),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_937),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_938),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_731),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_843),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_941),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_734),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_969),
.B(n_817),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_721),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_736),
.Y(n_1126)
);

BUFx5_ASAP7_75t_L g1127 ( 
.A(n_732),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_746),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_749),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_955),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_752),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1020),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1020),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_976),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_769),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_770),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_981),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_771),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1000),
.Y(n_1139)
);

BUFx2_ASAP7_75t_SL g1140 ( 
.A(n_810),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1013),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_843),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_775),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1029),
.Y(n_1144)
);

INVxp33_ASAP7_75t_SL g1145 ( 
.A(n_719),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_870),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_702),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_742),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_843),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_742),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_776),
.Y(n_1151)
);

BUFx5_ASAP7_75t_L g1152 ( 
.A(n_739),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_779),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_873),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_900),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_782),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_919),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_843),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1020),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_810),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_783),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_855),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_855),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_817),
.B(n_0),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_785),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_861),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_806),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_792),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_983),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_861),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_983),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_748),
.Y(n_1172)
);

INVxp33_ASAP7_75t_L g1173 ( 
.A(n_720),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_706),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_707),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_702),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_708),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_709),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_711),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_713),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_794),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_795),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_983),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_748),
.Y(n_1184)
);

BUFx5_ASAP7_75t_L g1185 ( 
.A(n_747),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_983),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_764),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_717),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_799),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_804),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_807),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_719),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_733),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_735),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_738),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_808),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_812),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_806),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_741),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_983),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_819),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_743),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_823),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_827),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_744),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_834),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_983),
.Y(n_1207)
);

BUFx10_ASAP7_75t_L g1208 ( 
.A(n_854),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_983),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_702),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_835),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_764),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_864),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_720),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_710),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_745),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_806),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_768),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_725),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_750),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_702),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_868),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_768),
.Y(n_1223)
);

BUFx10_ASAP7_75t_L g1224 ( 
.A(n_820),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_874),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_722),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_876),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_878),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_753),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_754),
.Y(n_1230)
);

BUFx8_ASAP7_75t_SL g1231 ( 
.A(n_856),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_848),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_881),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_756),
.Y(n_1234)
);

CKINVDCx16_ASAP7_75t_R g1235 ( 
.A(n_815),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_890),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_757),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_894),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_887),
.B(n_0),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_848),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_762),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_759),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_899),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_905),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_722),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_765),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_907),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_908),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_911),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_767),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_916),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_811),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_856),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_725),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_773),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_724),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_860),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_939),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_774),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_940),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_949),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_724),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_777),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_860),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_848),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_914),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_784),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_954),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_956),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_957),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_883),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_914),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_847),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_780),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_883),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_787),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_789),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_886),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_730),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_730),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_960),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_886),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_914),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_972),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_751),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_959),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_850),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_987),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_820),
.B(n_1),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_791),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_727),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_1001),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_793),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_959),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_811),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_1001),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_858),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_796),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_990),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_797),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_798),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_992),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_800),
.Y(n_1303)
);

INVx4_ASAP7_75t_R g1304 ( 
.A(n_718),
.Y(n_1304)
);

BUFx2_ASAP7_75t_SL g1305 ( 
.A(n_766),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_801),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_751),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_802),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_828),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_803),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_727),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_828),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_809),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1001),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_993),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_909),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1005),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1009),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1010),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1015),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_814),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1016),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_818),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_978),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_824),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1017),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1023),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_728),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1025),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1031),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_1012),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_889),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_909),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_912),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_825),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_928),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_928),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_970),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_1012),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_826),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_982),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_829),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_988),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_830),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_991),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1030),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_832),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_833),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_978),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_766),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_1012),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_971),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_778),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_836),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_839),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_778),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_840),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_822),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_822),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_842),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_844),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_845),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_728),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_971),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1003),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_846),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1003),
.Y(n_1367)
);

CKINVDCx14_ASAP7_75t_R g1368 ( 
.A(n_1026),
.Y(n_1368)
);

BUFx2_ASAP7_75t_SL g1369 ( 
.A(n_831),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_986),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_852),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1004),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_853),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1018),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1026),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_857),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_986),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_811),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1004),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1008),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1008),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_859),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1028),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1028),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_862),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_811),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_863),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1014),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_930),
.B(n_1),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_895),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_772),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_975),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1018),
.Y(n_1393)
);

BUFx10_ASAP7_75t_L g1394 ( 
.A(n_865),
.Y(n_1394)
);

BUFx8_ASAP7_75t_SL g1395 ( 
.A(n_1019),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_866),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_867),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_869),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1019),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_871),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1037),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1090),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1070),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1091),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1098),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1093),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1040),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1095),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1096),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_1375),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1097),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1102),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1103),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1043),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1104),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1049),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1052),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1053),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1106),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1055),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1108),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1057),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1064),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1369),
.B(n_1033),
.Y(n_1424)
);

CKINVDCx16_ASAP7_75t_R g1425 ( 
.A(n_1283),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1112),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1054),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1054),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1066),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1146),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1079),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1068),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1098),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1071),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1050),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1051),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1073),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1378),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1160),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1378),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1081),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1332),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1174),
.B(n_877),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_1192),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1334),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1338),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1085),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1341),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1343),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1345),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1086),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1092),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_L g1453 ( 
.A(n_1357),
.B(n_533),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1346),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1080),
.B(n_879),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1219),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1113),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1114),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1125),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1125),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1115),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1099),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1148),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1116),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1375),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1328),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1120),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1162),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1163),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1123),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1126),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1166),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1128),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1170),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1129),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1131),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1148),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1150),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1175),
.B(n_888),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1100),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1150),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1154),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1172),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1101),
.B(n_892),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1135),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1136),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1177),
.B(n_893),
.Y(n_1487)
);

INVxp33_ASAP7_75t_SL g1488 ( 
.A(n_1155),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1172),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1105),
.Y(n_1490)
);

INVxp33_ASAP7_75t_SL g1491 ( 
.A(n_1157),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1138),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1143),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_L g1494 ( 
.A(n_1109),
.B(n_535),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1151),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1184),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1111),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1047),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1153),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1156),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1161),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1165),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1140),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1118),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1119),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1168),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1181),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1184),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1182),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1189),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1122),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1190),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1191),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1130),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1178),
.B(n_897),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1196),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1187),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1197),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1201),
.Y(n_1519)
);

INVxp33_ASAP7_75t_SL g1520 ( 
.A(n_1134),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1203),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1137),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1139),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1204),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1206),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1141),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1211),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1144),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1187),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1213),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1222),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1179),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1047),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1147),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1080),
.B(n_898),
.Y(n_1535)
);

INVxp33_ASAP7_75t_SL g1536 ( 
.A(n_1180),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1188),
.B(n_901),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1225),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1193),
.Y(n_1539)
);

CKINVDCx14_ASAP7_75t_R g1540 ( 
.A(n_1368),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1374),
.Y(n_1541)
);

INVxp33_ASAP7_75t_L g1542 ( 
.A(n_1254),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1194),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1212),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1291),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1311),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1195),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1227),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1228),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1199),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1212),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1218),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1202),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1218),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1056),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1233),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1235),
.B(n_902),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1056),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1223),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1236),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1205),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1216),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1238),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1223),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1253),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1147),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1220),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1229),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1243),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1396),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1400),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1147),
.Y(n_1572)
);

NOR2xp67_ASAP7_75t_L g1573 ( 
.A(n_1230),
.B(n_536),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1234),
.B(n_1237),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1244),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1368),
.B(n_903),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1241),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1246),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1253),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1393),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1386),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1247),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1250),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1255),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1248),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1257),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1259),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1249),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1263),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1274),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1276),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1251),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1277),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1290),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1258),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1293),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1260),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1261),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1298),
.Y(n_1599)
);

INVxp33_ASAP7_75t_SL g1600 ( 
.A(n_1300),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1301),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1147),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1303),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1306),
.B(n_904),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1268),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1269),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1308),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1257),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_1292),
.Y(n_1609)
);

NOR2xp67_ASAP7_75t_L g1610 ( 
.A(n_1310),
.B(n_539),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1270),
.Y(n_1611)
);

CKINVDCx14_ASAP7_75t_R g1612 ( 
.A(n_1076),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1264),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1386),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1313),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1363),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1321),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1281),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1391),
.B(n_884),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1176),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1284),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1288),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1299),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1302),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1315),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1264),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1317),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1271),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1323),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1318),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1319),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1325),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1335),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1271),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1275),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1275),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1320),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1322),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1176),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1340),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1242),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1326),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1327),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1329),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1393),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1167),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1342),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1330),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1059),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1217),
.B(n_1265),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1344),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1370),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1347),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1348),
.Y(n_1654)
);

NOR2xp67_ASAP7_75t_L g1655 ( 
.A(n_1354),
.B(n_542),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1060),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1278),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1355),
.B(n_913),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1360),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1361),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1278),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1362),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1061),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1062),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1366),
.B(n_915),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1063),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1371),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1388),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1373),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1376),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1382),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1385),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1242),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1282),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1065),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1282),
.Y(n_1676)
);

BUFx10_ASAP7_75t_L g1677 ( 
.A(n_1387),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1397),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1067),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1069),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1176),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1286),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1398),
.Y(n_1683)
);

NOR2xp67_ASAP7_75t_L g1684 ( 
.A(n_1272),
.B(n_543),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1072),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1074),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1395),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1399),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1078),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1082),
.Y(n_1690)
);

CKINVDCx20_ASAP7_75t_R g1691 ( 
.A(n_1286),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1395),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1231),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1231),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1266),
.Y(n_1695)
);

NOR2xp67_ASAP7_75t_L g1696 ( 
.A(n_1117),
.B(n_544),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1176),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1083),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1087),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1088),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1089),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1394),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1294),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1038),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1394),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1039),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1498),
.B(n_1390),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1572),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1581),
.B(n_1314),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1534),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1619),
.A2(n_1124),
.B1(n_1289),
.B2(n_1164),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1533),
.B(n_1392),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1704),
.A2(n_1706),
.B(n_1566),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1572),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1572),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1534),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1649),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1424),
.A2(n_1389),
.B1(n_1399),
.B2(n_1145),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1566),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1646),
.Y(n_1720)
);

BUFx12f_ASAP7_75t_L g1721 ( 
.A(n_1677),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1620),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1494),
.B(n_1296),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1695),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1555),
.B(n_1215),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1620),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1650),
.B(n_891),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1572),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1614),
.B(n_1215),
.Y(n_1729)
);

CKINVDCx8_ASAP7_75t_R g1730 ( 
.A(n_1425),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1602),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1602),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1656),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1639),
.A2(n_1044),
.B(n_1041),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1558),
.B(n_1214),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1663),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1664),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1666),
.Y(n_1738)
);

CKINVDCx8_ASAP7_75t_R g1739 ( 
.A(n_1609),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1675),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1679),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1456),
.A2(n_1389),
.B1(n_1145),
.B2(n_1239),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1652),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1405),
.A2(n_1294),
.B1(n_1349),
.B2(n_1324),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1602),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1639),
.A2(n_1046),
.B(n_1045),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1680),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1602),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1641),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1438),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1681),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1641),
.B(n_1214),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1440),
.B(n_1048),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1673),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1681),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1697),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1668),
.B(n_1058),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1612),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1697),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1402),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1466),
.A2(n_896),
.B1(n_997),
.B2(n_921),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1673),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1404),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1406),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1685),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1557),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1541),
.A2(n_1042),
.B1(n_998),
.B2(n_1022),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1444),
.B(n_1540),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1686),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1573),
.B(n_1305),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1401),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1545),
.A2(n_1042),
.B1(n_1022),
.B2(n_1027),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1612),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1443),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1427),
.B(n_1094),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1428),
.B(n_1094),
.Y(n_1777)
);

OA21x2_ASAP7_75t_L g1778 ( 
.A1(n_1408),
.A2(n_1353),
.B(n_1350),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1442),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1689),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1407),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1409),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1445),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1690),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1414),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1698),
.Y(n_1786)
);

AND2x6_ASAP7_75t_L g1787 ( 
.A(n_1455),
.B(n_1075),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1411),
.A2(n_1413),
.B(n_1412),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1444),
.B(n_1540),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1435),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1415),
.A2(n_1421),
.B(n_1419),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1405),
.A2(n_1349),
.B1(n_1377),
.B2(n_1324),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1426),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1446),
.B(n_1094),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1448),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1699),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1457),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1449),
.B(n_1094),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1458),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1477),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1700),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1701),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1461),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1450),
.B(n_1094),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1454),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1436),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1464),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1542),
.B(n_1058),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1467),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1542),
.B(n_1077),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1478),
.Y(n_1811)
);

OA21x2_ASAP7_75t_L g1812 ( 
.A1(n_1484),
.A2(n_1358),
.B(n_1356),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1479),
.B(n_1077),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1470),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1410),
.B(n_1094),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1433),
.A2(n_1377),
.B1(n_1027),
.B2(n_1021),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1471),
.Y(n_1817)
);

BUFx8_ASAP7_75t_L g1818 ( 
.A(n_1580),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1535),
.A2(n_1084),
.B(n_1075),
.Y(n_1819)
);

AND2x2_ASAP7_75t_SL g1820 ( 
.A(n_1645),
.B(n_1331),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1473),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1475),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1487),
.B(n_1110),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1476),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1485),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1486),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1492),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1493),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1465),
.B(n_1495),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1499),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1500),
.B(n_1094),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1515),
.B(n_1110),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1501),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1502),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1537),
.B(n_1132),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1506),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1507),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1509),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1510),
.B(n_1226),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1512),
.B(n_1226),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1513),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1516),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1518),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1519),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1521),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1524),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1430),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1604),
.B(n_1132),
.Y(n_1848)
);

OA21x2_ASAP7_75t_L g1849 ( 
.A1(n_1525),
.A2(n_1359),
.B(n_1107),
.Y(n_1849)
);

AND2x6_ASAP7_75t_L g1850 ( 
.A(n_1574),
.B(n_1084),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1546),
.A2(n_1021),
.B1(n_1173),
.B2(n_917),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1658),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1527),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1530),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1616),
.A2(n_1173),
.B1(n_918),
.B2(n_923),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1531),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1538),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1548),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1439),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1549),
.Y(n_1860)
);

OA21x2_ASAP7_75t_L g1861 ( 
.A1(n_1556),
.A2(n_1121),
.B(n_1107),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1560),
.B(n_1127),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1563),
.B(n_1245),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1569),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1575),
.B(n_1245),
.Y(n_1865)
);

OAI22x1_ASAP7_75t_SL g1866 ( 
.A1(n_1433),
.A2(n_920),
.B1(n_924),
.B2(n_922),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1582),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1585),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1588),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1481),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1592),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1595),
.Y(n_1872)
);

BUFx12f_ASAP7_75t_L g1873 ( 
.A(n_1677),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1597),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1598),
.A2(n_1142),
.B(n_1121),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1605),
.B(n_1256),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1403),
.A2(n_925),
.B1(n_932),
.B2(n_931),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1606),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1611),
.B(n_1256),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1431),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1618),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1621),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1622),
.B(n_1623),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1624),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1625),
.B(n_1627),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1630),
.Y(n_1886)
);

CKINVDCx16_ASAP7_75t_R g1887 ( 
.A(n_1483),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1631),
.B(n_1262),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1637),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1638),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1642),
.B(n_1262),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1643),
.B(n_1644),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1503),
.A2(n_929),
.B1(n_942),
.B2(n_936),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1696),
.A2(n_935),
.B1(n_945),
.B2(n_944),
.Y(n_1894)
);

CKINVDCx6p67_ASAP7_75t_R g1895 ( 
.A(n_1677),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1648),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1576),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1532),
.A2(n_943),
.B1(n_951),
.B2(n_948),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1665),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1453),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1684),
.B(n_1279),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1610),
.B(n_1279),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1416),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1543),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1640),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1669),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1655),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1482),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1417),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1539),
.B(n_1133),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1547),
.A2(n_968),
.B1(n_989),
.B2(n_952),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1468),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1418),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1420),
.A2(n_1149),
.B(n_1142),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1688),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1422),
.Y(n_1916)
);

OA21x2_ASAP7_75t_L g1917 ( 
.A1(n_1423),
.A2(n_1158),
.B(n_1149),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1520),
.B(n_1133),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1459),
.A2(n_1351),
.B1(n_1339),
.B2(n_958),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1429),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1432),
.B(n_1280),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1434),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1437),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1441),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1447),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1451),
.A2(n_1169),
.B(n_1158),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1469),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1452),
.B(n_1127),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1550),
.Y(n_1929)
);

OAI22x1_ASAP7_75t_L g1930 ( 
.A1(n_1702),
.A2(n_1232),
.B1(n_1240),
.B2(n_1198),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1553),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1459),
.A2(n_961),
.B1(n_962),
.B2(n_947),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1462),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1489),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1480),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1490),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1497),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1561),
.B(n_1159),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1504),
.Y(n_1939)
);

CKINVDCx11_ASAP7_75t_R g1940 ( 
.A(n_1460),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1505),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1511),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1514),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1522),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1523),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1526),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1528),
.B(n_1127),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1562),
.B(n_1280),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1536),
.B(n_1159),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1567),
.B(n_1208),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1568),
.Y(n_1951)
);

INVx4_ASAP7_75t_L g1952 ( 
.A(n_1577),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1578),
.Y(n_1953)
);

INVx5_ASAP7_75t_L g1954 ( 
.A(n_1600),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1583),
.Y(n_1955)
);

AND2x6_ASAP7_75t_L g1956 ( 
.A(n_1488),
.B(n_1169),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1584),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1587),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1589),
.A2(n_963),
.B1(n_967),
.B2(n_966),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1590),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1591),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1593),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1594),
.A2(n_995),
.B1(n_1035),
.B2(n_973),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1596),
.Y(n_1964)
);

AND2x6_ASAP7_75t_L g1965 ( 
.A(n_1491),
.B(n_1171),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1599),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1601),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1603),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1607),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1615),
.B(n_1127),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1617),
.B(n_1285),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1629),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1632),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1633),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1647),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1651),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1653),
.B(n_1208),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1654),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1659),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1660),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1662),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1667),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1670),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1671),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1672),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1678),
.B(n_1285),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1683),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1705),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1687),
.A2(n_965),
.B1(n_979),
.B2(n_977),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1472),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1692),
.Y(n_1991)
);

BUFx2_ASAP7_75t_L g1992 ( 
.A(n_1554),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1693),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1474),
.B(n_1394),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_SL g1995 ( 
.A1(n_1460),
.A2(n_980),
.B1(n_984),
.B2(n_974),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1899),
.B(n_1815),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1734),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1734),
.Y(n_1998)
);

CKINVDCx16_ASAP7_75t_R g1999 ( 
.A(n_1887),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1753),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1753),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1709),
.B(n_1224),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1839),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1743),
.B(n_1224),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_SL g2005 ( 
.A(n_1897),
.B(n_985),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1747),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1747),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1839),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1750),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1760),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1861),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1840),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1861),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1850),
.B(n_1127),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1840),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1850),
.B(n_1928),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1779),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1850),
.B(n_1127),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1797),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1775),
.B(n_1208),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1850),
.B(n_1127),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1863),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1815),
.B(n_1152),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1760),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1720),
.B(n_1224),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1928),
.B(n_1152),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1863),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1875),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1729),
.B(n_1267),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1865),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1760),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1875),
.Y(n_2032)
);

OA21x2_ASAP7_75t_L g2033 ( 
.A1(n_1713),
.A2(n_1798),
.B(n_1794),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1865),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1947),
.B(n_1152),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1849),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1779),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1876),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1799),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1876),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1849),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1763),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1879),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1778),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1778),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1879),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_1763),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1779),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1888),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1888),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1755),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1808),
.B(n_1267),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1947),
.B(n_1970),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1783),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1970),
.B(n_1152),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1788),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1788),
.Y(n_2057)
);

INVx6_ASAP7_75t_L g2058 ( 
.A(n_1954),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1891),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1775),
.B(n_994),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1891),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1752),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1809),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1822),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1752),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1825),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1828),
.Y(n_2067)
);

OA21x2_ASAP7_75t_L g2068 ( 
.A1(n_1794),
.A2(n_1183),
.B(n_1171),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1837),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1819),
.A2(n_1186),
.B(n_1183),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1735),
.B(n_1365),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1841),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1846),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1791),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1791),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1798),
.A2(n_1200),
.B(n_1186),
.Y(n_2076)
);

OA21x2_ASAP7_75t_L g2077 ( 
.A1(n_1804),
.A2(n_1207),
.B(n_1200),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1783),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1853),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1710),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1716),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1856),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1719),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1725),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1722),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1746),
.B(n_1152),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_SL g2087 ( 
.A1(n_1744),
.A2(n_1496),
.B1(n_1508),
.B2(n_1463),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1897),
.B(n_1152),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1857),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1726),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1735),
.B(n_1367),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1860),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1864),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1903),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_1725),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1783),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1869),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1756),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1913),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1872),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1810),
.B(n_1273),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1746),
.B(n_1152),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1859),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1878),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1757),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1756),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1882),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1795),
.Y(n_2108)
);

OA21x2_ASAP7_75t_L g2109 ( 
.A1(n_1804),
.A2(n_1862),
.B(n_1831),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1795),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1914),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1795),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1886),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1724),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1805),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1889),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1829),
.B(n_1185),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1896),
.Y(n_2118)
);

HB1xp67_ASAP7_75t_L g2119 ( 
.A(n_1921),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1803),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_1744),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_1833),
.B(n_1372),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_1915),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1852),
.B(n_1185),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1717),
.Y(n_2125)
);

INVxp67_ASAP7_75t_L g2126 ( 
.A(n_1880),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_1915),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1921),
.B(n_1273),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1829),
.B(n_1185),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1948),
.B(n_1287),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1805),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1733),
.Y(n_2132)
);

INVxp67_ASAP7_75t_L g2133 ( 
.A(n_1880),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1914),
.Y(n_2134)
);

INVx1_ASAP7_75t_SL g2135 ( 
.A(n_1759),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1917),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1736),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1852),
.B(n_1185),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1907),
.B(n_1185),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1917),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1948),
.B(n_1185),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1805),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1844),
.B(n_1185),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1844),
.B(n_1287),
.Y(n_2144)
);

INVx6_ASAP7_75t_L g2145 ( 
.A(n_1954),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1926),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1737),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1738),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1740),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1883),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1926),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1741),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1748),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1971),
.B(n_1207),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1884),
.B(n_1297),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1766),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1770),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1884),
.B(n_1297),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1883),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1971),
.B(n_1986),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1754),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1754),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1912),
.Y(n_2163)
);

INVxp67_ASAP7_75t_L g2164 ( 
.A(n_1727),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1986),
.B(n_1910),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1761),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1780),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1813),
.B(n_1210),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1784),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1786),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1796),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1885),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1801),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1823),
.B(n_1210),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1802),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1751),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1751),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1807),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1817),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1821),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1814),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1824),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_1885),
.B(n_1379),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1826),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1814),
.B(n_1209),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1842),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1814),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1764),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_1892),
.B(n_1380),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1867),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1765),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1868),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_1938),
.B(n_1381),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1827),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1892),
.Y(n_2195)
);

NAND2xp33_ASAP7_75t_SL g2196 ( 
.A(n_1767),
.B(n_996),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1790),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_1707),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_1774),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1832),
.B(n_1835),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1782),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1793),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1790),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1812),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1806),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1812),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1848),
.B(n_1210),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1806),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1776),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1831),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1862),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1827),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1776),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1771),
.B(n_1210),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1777),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1827),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1707),
.B(n_1383),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1830),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1830),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_1712),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_1712),
.B(n_1384),
.Y(n_2221)
);

INVx3_ASAP7_75t_L g2222 ( 
.A(n_1830),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1771),
.B(n_1902),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1834),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1777),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1834),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_1834),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1836),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1836),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1836),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_1800),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1838),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1838),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1838),
.B(n_1307),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1843),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1843),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1843),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1845),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1845),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1845),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1854),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_1811),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1854),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_SL g2244 ( 
.A1(n_1792),
.A2(n_1496),
.B1(n_1508),
.B2(n_1463),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1854),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_1858),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1858),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1858),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1871),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1871),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1871),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1874),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_1901),
.A2(n_1209),
.B(n_1307),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1874),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1874),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1881),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1881),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1708),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1902),
.B(n_1787),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1787),
.B(n_1221),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1881),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_1870),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1890),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1890),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1890),
.Y(n_2265)
);

INVx1_ASAP7_75t_SL g2266 ( 
.A(n_1769),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1727),
.B(n_1758),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1901),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1708),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_1758),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1708),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1714),
.Y(n_2272)
);

INVxp67_ASAP7_75t_L g2273 ( 
.A(n_1918),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1904),
.B(n_1309),
.Y(n_2274)
);

INVx6_ASAP7_75t_L g2275 ( 
.A(n_1954),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_1905),
.B(n_1309),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1787),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1787),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1900),
.B(n_1221),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1714),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1906),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_1714),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_1715),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_1934),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1908),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1715),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1715),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1732),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1732),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1732),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_1749),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1918),
.B(n_1312),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_SL g2293 ( 
.A(n_1895),
.B(n_1772),
.Y(n_2293)
);

INVxp33_ASAP7_75t_SL g2294 ( 
.A(n_1792),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_1923),
.B(n_1312),
.Y(n_2295)
);

INVx6_ASAP7_75t_L g2296 ( 
.A(n_1913),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1742),
.B(n_1221),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1927),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1749),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_1992),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_1749),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1956),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1956),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_1728),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1956),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1956),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1965),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_1789),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_1937),
.B(n_1316),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1965),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1965),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_1941),
.B(n_1316),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_1942),
.B(n_1333),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1949),
.B(n_1333),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1728),
.Y(n_2315)
);

INVx4_ASAP7_75t_L g2316 ( 
.A(n_1965),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2080),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_2114),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2080),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2000),
.Y(n_2320)
);

INVx5_ASAP7_75t_L g2321 ( 
.A(n_2007),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2001),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2099),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2081),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2234),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2161),
.B(n_1742),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2234),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2003),
.Y(n_2328)
);

NAND2xp33_ASAP7_75t_L g2329 ( 
.A(n_2017),
.B(n_1924),
.Y(n_2329)
);

INVx4_ASAP7_75t_L g2330 ( 
.A(n_2296),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2161),
.B(n_1711),
.Y(n_2331)
);

CKINVDCx16_ASAP7_75t_R g2332 ( 
.A(n_1999),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2081),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_2099),
.Y(n_2334)
);

INVx4_ASAP7_75t_L g2335 ( 
.A(n_2296),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2094),
.Y(n_2336)
);

INVx2_ASAP7_75t_SL g2337 ( 
.A(n_2114),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2008),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_SL g2339 ( 
.A(n_2009),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2083),
.Y(n_2340)
);

BUFx4f_ASAP7_75t_L g2341 ( 
.A(n_2296),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2012),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2009),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2083),
.Y(n_2344)
);

INVx1_ASAP7_75t_SL g2345 ( 
.A(n_2123),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2208),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2208),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2015),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2127),
.B(n_1887),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2022),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2027),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2085),
.Y(n_2352)
);

INVx3_ASAP7_75t_L g2353 ( 
.A(n_2017),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2085),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2002),
.B(n_1913),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2017),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2042),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2200),
.B(n_1916),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_SL g2359 ( 
.A(n_2051),
.Y(n_2359)
);

AND2x2_ASAP7_75t_SL g2360 ( 
.A(n_2293),
.B(n_1916),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_2198),
.Y(n_2361)
);

OAI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2162),
.A2(n_1718),
.B1(n_1711),
.B2(n_1762),
.Y(n_2362)
);

OAI22xp33_ASAP7_75t_L g2363 ( 
.A1(n_2162),
.A2(n_1718),
.B1(n_1762),
.B2(n_1911),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2030),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2051),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2034),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2017),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2210),
.B(n_1949),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2037),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2090),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2160),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2150),
.B(n_1916),
.Y(n_2372)
);

BUFx10_ASAP7_75t_L g2373 ( 
.A(n_2020),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2038),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2090),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2040),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2105),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2273),
.B(n_1929),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2037),
.Y(n_2379)
);

OR2x2_ASAP7_75t_L g2380 ( 
.A(n_2126),
.B(n_1847),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2043),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2105),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1997),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2150),
.B(n_1920),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_2209),
.A2(n_2213),
.B1(n_2225),
.B2(n_2215),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1997),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2004),
.B(n_1950),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2211),
.B(n_1945),
.Y(n_2388)
);

INVx3_ASAP7_75t_L g2389 ( 
.A(n_2037),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_2209),
.A2(n_1995),
.B1(n_1932),
.B2(n_1816),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_SL g2391 ( 
.A(n_2316),
.B(n_1772),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2046),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2159),
.B(n_1920),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2049),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2159),
.B(n_1920),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_2135),
.Y(n_2396)
);

BUFx3_ASAP7_75t_L g2397 ( 
.A(n_2284),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1998),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2050),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2053),
.B(n_1957),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2059),
.Y(n_2401)
);

NAND2xp33_ASAP7_75t_R g2402 ( 
.A(n_2300),
.B(n_1694),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2103),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1998),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2163),
.Y(n_2405)
);

INVx5_ASAP7_75t_L g2406 ( 
.A(n_2007),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2298),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2273),
.B(n_1929),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2087),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2213),
.A2(n_1995),
.B1(n_1932),
.B2(n_1816),
.Y(n_2410)
);

AND2x6_ASAP7_75t_L g2411 ( 
.A(n_2111),
.B(n_1924),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2215),
.B(n_1966),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2006),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2061),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2198),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2006),
.Y(n_2416)
);

INVxp33_ASAP7_75t_L g2417 ( 
.A(n_2025),
.Y(n_2417)
);

INVx4_ASAP7_75t_L g2418 ( 
.A(n_2037),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2042),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2225),
.B(n_1974),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2048),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2220),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2270),
.B(n_1781),
.Y(n_2423)
);

XNOR2xp5_ASAP7_75t_L g2424 ( 
.A(n_2244),
.B(n_1551),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2036),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2270),
.B(n_1781),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2164),
.A2(n_1911),
.B1(n_1963),
.B2(n_1962),
.Y(n_2427)
);

OR2x2_ASAP7_75t_L g2428 ( 
.A(n_2126),
.B(n_1990),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2164),
.B(n_1785),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2020),
.B(n_1785),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_SL g2431 ( 
.A(n_2172),
.B(n_1924),
.Y(n_2431)
);

INVx3_ASAP7_75t_L g2432 ( 
.A(n_2048),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2048),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_1996),
.B(n_1975),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2056),
.A2(n_2074),
.B1(n_2075),
.B2(n_2057),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2036),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2220),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2041),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2274),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2172),
.B(n_1925),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2041),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_1996),
.B(n_1978),
.Y(n_2442)
);

INVx5_ASAP7_75t_L g2443 ( 
.A(n_2007),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2274),
.Y(n_2444)
);

AO22x2_ASAP7_75t_L g2445 ( 
.A1(n_2267),
.A2(n_1773),
.B1(n_1768),
.B2(n_1894),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2276),
.Y(n_2446)
);

AND2x6_ASAP7_75t_L g2447 ( 
.A(n_2111),
.B(n_2134),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2276),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2056),
.A2(n_1768),
.B1(n_1773),
.B2(n_1894),
.Y(n_2449)
);

INVx2_ASAP7_75t_SL g2450 ( 
.A(n_2122),
.Y(n_2450)
);

AOI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2267),
.A2(n_2141),
.B1(n_2129),
.B2(n_2117),
.Y(n_2451)
);

NAND2xp33_ASAP7_75t_L g2452 ( 
.A(n_2048),
.B(n_1944),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2133),
.B(n_2060),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2057),
.A2(n_1851),
.B1(n_1855),
.B2(n_1877),
.Y(n_2454)
);

BUFx10_ASAP7_75t_L g2455 ( 
.A(n_2060),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2122),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_2165),
.B(n_1925),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2054),
.B(n_1925),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2054),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2054),
.B(n_1933),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2074),
.A2(n_1851),
.B1(n_1855),
.B2(n_1877),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2063),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2064),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2166),
.Y(n_2464)
);

OAI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_2133),
.A2(n_1963),
.B1(n_1933),
.B2(n_1944),
.Y(n_2465)
);

XNOR2xp5_ASAP7_75t_L g2466 ( 
.A(n_2231),
.B(n_1551),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2054),
.B(n_1933),
.Y(n_2467)
);

AOI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2141),
.A2(n_1723),
.B1(n_1922),
.B2(n_1909),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2078),
.B(n_1943),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2066),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_2295),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_SL g2472 ( 
.A(n_2281),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2067),
.Y(n_2473)
);

INVx4_ASAP7_75t_SL g2474 ( 
.A(n_2007),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2069),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2078),
.B(n_1943),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2166),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2072),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2188),
.Y(n_2479)
);

AOI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2075),
.A2(n_1919),
.B1(n_999),
.B2(n_1006),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2078),
.B(n_1943),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2073),
.Y(n_2482)
);

INVxp33_ASAP7_75t_L g2483 ( 
.A(n_2231),
.Y(n_2483)
);

BUFx10_ASAP7_75t_L g2484 ( 
.A(n_2058),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2029),
.B(n_1977),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2188),
.Y(n_2486)
);

INVx2_ASAP7_75t_SL g2487 ( 
.A(n_2295),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2078),
.B(n_1944),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2191),
.Y(n_2489)
);

BUFx10_ASAP7_75t_L g2490 ( 
.A(n_2058),
.Y(n_2490)
);

INVx8_ASAP7_75t_L g2491 ( 
.A(n_2096),
.Y(n_2491)
);

OR2x6_ASAP7_75t_L g2492 ( 
.A(n_2058),
.B(n_1946),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2191),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2079),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2201),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2266),
.B(n_2308),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2082),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2089),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2047),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2047),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2092),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2308),
.B(n_1952),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2093),
.Y(n_2503)
);

INVx4_ASAP7_75t_L g2504 ( 
.A(n_2096),
.Y(n_2504)
);

AOI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2117),
.A2(n_1723),
.B1(n_1983),
.B2(n_1981),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2124),
.B(n_1982),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2201),
.Y(n_2507)
);

AOI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2129),
.A2(n_1935),
.B1(n_1939),
.B2(n_1936),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2119),
.B(n_1952),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2138),
.B(n_1987),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2119),
.B(n_1931),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_2242),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2202),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2097),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_L g2515 ( 
.A1(n_2204),
.A2(n_1919),
.B1(n_1002),
.B2(n_1032),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2100),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2084),
.B(n_1951),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2202),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2242),
.Y(n_2519)
);

INVxp33_ASAP7_75t_L g2520 ( 
.A(n_2262),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2104),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2096),
.B(n_1946),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2086),
.B(n_1958),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2107),
.Y(n_2524)
);

INVx5_ASAP7_75t_L g2525 ( 
.A(n_2316),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2134),
.A2(n_2136),
.B1(n_2146),
.B2(n_2140),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2195),
.B(n_1946),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2113),
.Y(n_2528)
);

OAI22xp33_ASAP7_75t_SL g2529 ( 
.A1(n_2294),
.A2(n_1898),
.B1(n_1959),
.B2(n_1973),
.Y(n_2529)
);

HB1xp67_ASAP7_75t_L g2530 ( 
.A(n_2084),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2096),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2095),
.B(n_1960),
.Y(n_2532)
);

INVx3_ASAP7_75t_L g2533 ( 
.A(n_2108),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2108),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_2262),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2102),
.B(n_1961),
.Y(n_2536)
);

BUFx8_ASAP7_75t_SL g2537 ( 
.A(n_2121),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2011),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2011),
.Y(n_2539)
);

AOI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2204),
.A2(n_1011),
.B1(n_1034),
.B2(n_1898),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2154),
.A2(n_1964),
.B1(n_1968),
.B2(n_1967),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2176),
.B(n_1976),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2095),
.B(n_1953),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2177),
.B(n_1979),
.Y(n_2544)
);

BUFx4f_ASAP7_75t_L g2545 ( 
.A(n_2145),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2016),
.B(n_1980),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2013),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2013),
.Y(n_2548)
);

AND2x4_ASAP7_75t_L g2549 ( 
.A(n_2183),
.B(n_1953),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2028),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2116),
.Y(n_2551)
);

AND2x6_ASAP7_75t_L g2552 ( 
.A(n_2136),
.B(n_1953),
.Y(n_2552)
);

INVx5_ASAP7_75t_L g2553 ( 
.A(n_2108),
.Y(n_2553)
);

OR2x2_ASAP7_75t_L g2554 ( 
.A(n_2199),
.B(n_1962),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2206),
.A2(n_1959),
.B1(n_1893),
.B2(n_1337),
.Y(n_2555)
);

AND2x2_ASAP7_75t_SL g2556 ( 
.A(n_2128),
.B(n_1955),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2052),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2028),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2292),
.B(n_1988),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2314),
.B(n_1969),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2140),
.B(n_1955),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2032),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2146),
.B(n_1955),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2108),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2206),
.A2(n_1893),
.B1(n_1337),
.B2(n_1352),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2285),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2309),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2110),
.B(n_1972),
.Y(n_2568)
);

INVx5_ASAP7_75t_L g2569 ( 
.A(n_2110),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2193),
.B(n_1972),
.Y(n_2570)
);

INVx2_ASAP7_75t_SL g2571 ( 
.A(n_2309),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2110),
.Y(n_2572)
);

INVxp67_ASAP7_75t_SL g2573 ( 
.A(n_2282),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2118),
.Y(n_2574)
);

BUFx2_ASAP7_75t_L g2575 ( 
.A(n_2130),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2145),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2125),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2032),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2110),
.B(n_1972),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2112),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2101),
.B(n_1969),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2112),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2132),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2112),
.B(n_1984),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2183),
.B(n_1984),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2151),
.A2(n_1352),
.B1(n_1336),
.B2(n_1820),
.Y(n_2586)
);

INVx5_ASAP7_75t_L g2587 ( 
.A(n_2112),
.Y(n_2587)
);

INVx1_ASAP7_75t_SL g2588 ( 
.A(n_2005),
.Y(n_2588)
);

NOR2x1p5_ASAP7_75t_L g2589 ( 
.A(n_2137),
.B(n_1721),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2115),
.B(n_1984),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2151),
.B(n_1985),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2147),
.Y(n_2592)
);

INVx4_ASAP7_75t_L g2593 ( 
.A(n_2115),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2312),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2148),
.Y(n_2595)
);

AOI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2154),
.A2(n_1985),
.B1(n_1930),
.B2(n_1994),
.Y(n_2596)
);

AND2x6_ASAP7_75t_L g2597 ( 
.A(n_2302),
.B(n_1985),
.Y(n_2597)
);

BUFx3_ASAP7_75t_L g2598 ( 
.A(n_2312),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2149),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2217),
.B(n_1994),
.Y(n_2600)
);

OR2x2_ASAP7_75t_L g2601 ( 
.A(n_2221),
.B(n_1991),
.Y(n_2601)
);

AND2x6_ASAP7_75t_L g2602 ( 
.A(n_2303),
.B(n_1991),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2106),
.Y(n_2603)
);

AOI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2088),
.A2(n_1873),
.B1(n_1866),
.B2(n_1989),
.Y(n_2604)
);

OR2x2_ASAP7_75t_L g2605 ( 
.A(n_2221),
.B(n_1989),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2106),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2305),
.A2(n_1739),
.B1(n_1730),
.B2(n_1682),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2152),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2115),
.Y(n_2609)
);

OR2x6_ASAP7_75t_L g2610 ( 
.A(n_2145),
.B(n_1993),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2153),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2071),
.B(n_1993),
.Y(n_2612)
);

INVxp33_ASAP7_75t_L g2613 ( 
.A(n_2189),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2115),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2131),
.B(n_1993),
.Y(n_2615)
);

NOR3xp33_ASAP7_75t_L g2616 ( 
.A(n_2005),
.B(n_1940),
.C(n_1304),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2156),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2275),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2109),
.B(n_2197),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2157),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2131),
.Y(n_2621)
);

AND2x6_ASAP7_75t_L g2622 ( 
.A(n_2306),
.B(n_1336),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2044),
.A2(n_1364),
.B1(n_1529),
.B2(n_1517),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2167),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2044),
.A2(n_2045),
.B1(n_2278),
.B2(n_2277),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2313),
.Y(n_2626)
);

INVx3_ASAP7_75t_L g2627 ( 
.A(n_2131),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2071),
.B(n_1517),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_2297),
.B(n_1745),
.C(n_1818),
.Y(n_2629)
);

XOR2xp5_ASAP7_75t_L g2630 ( 
.A(n_2121),
.B(n_1529),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_L g2631 ( 
.A(n_2131),
.B(n_1221),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2169),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2142),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2109),
.B(n_1745),
.Y(n_2634)
);

INVx6_ASAP7_75t_L g2635 ( 
.A(n_2275),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2142),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2091),
.B(n_1544),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2196),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2170),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2142),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_2275),
.Y(n_2641)
);

NOR2x1p5_ASAP7_75t_L g2642 ( 
.A(n_2171),
.B(n_1866),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2173),
.Y(n_2643)
);

CKINVDCx6p67_ASAP7_75t_R g2644 ( 
.A(n_2189),
.Y(n_2644)
);

AOI22xp33_ASAP7_75t_L g2645 ( 
.A1(n_2045),
.A2(n_1364),
.B1(n_1552),
.B2(n_1544),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2175),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2019),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2039),
.Y(n_2648)
);

OR2x6_ASAP7_75t_L g2649 ( 
.A(n_2307),
.B(n_1818),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2120),
.Y(n_2650)
);

INVx4_ASAP7_75t_L g2651 ( 
.A(n_2142),
.Y(n_2651)
);

BUFx8_ASAP7_75t_SL g2652 ( 
.A(n_2313),
.Y(n_2652)
);

INVx4_ASAP7_75t_L g2653 ( 
.A(n_2181),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2253),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2253),
.Y(n_2655)
);

AND3x2_ASAP7_75t_L g2656 ( 
.A(n_2310),
.B(n_821),
.C(n_1552),
.Y(n_2656)
);

BUFx10_ASAP7_75t_L g2657 ( 
.A(n_2091),
.Y(n_2657)
);

INVx4_ASAP7_75t_L g2658 ( 
.A(n_2181),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2181),
.Y(n_2659)
);

OAI22xp33_ASAP7_75t_SL g2660 ( 
.A1(n_2297),
.A2(n_1364),
.B1(n_4),
.B2(n_2),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2268),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2181),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2109),
.B(n_1731),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2203),
.B(n_1731),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2178),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2187),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2253),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2179),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2180),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2062),
.Y(n_2670)
);

INVx1_ASAP7_75t_SL g2671 ( 
.A(n_2168),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2465),
.B(n_2570),
.Y(n_2672)
);

NAND3xp33_ASAP7_75t_SL g2673 ( 
.A(n_2515),
.B(n_1564),
.C(n_1559),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2465),
.B(n_2187),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2570),
.B(n_2187),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2400),
.B(n_2144),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2400),
.B(n_2155),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2383),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_2556),
.B(n_2187),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2386),
.Y(n_2680)
);

NAND2xp33_ASAP7_75t_L g2681 ( 
.A(n_2597),
.B(n_2194),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2462),
.Y(n_2682)
);

NOR3xp33_ASAP7_75t_L g2683 ( 
.A(n_2430),
.B(n_2196),
.C(n_2223),
.Y(n_2683)
);

NAND3xp33_ASAP7_75t_L g2684 ( 
.A(n_2453),
.B(n_2207),
.C(n_2174),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2463),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2378),
.A2(n_2218),
.B1(n_2219),
.B2(n_2212),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2455),
.B(n_2194),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_L g2688 ( 
.A(n_2323),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2470),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_L g2690 ( 
.A(n_2408),
.B(n_2368),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2455),
.B(n_2560),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2473),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2323),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2398),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2404),
.Y(n_2695)
);

INVx2_ASAP7_75t_SL g2696 ( 
.A(n_2535),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2519),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2368),
.B(n_2194),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2412),
.B(n_2158),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2412),
.B(n_2205),
.Y(n_2700)
);

NOR2xp67_ASAP7_75t_L g2701 ( 
.A(n_2336),
.B(n_2182),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2420),
.B(n_2226),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2413),
.Y(n_2703)
);

BUFx5_ASAP7_75t_L g2704 ( 
.A(n_2447),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2420),
.B(n_2226),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2475),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2478),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2600),
.A2(n_2229),
.B1(n_2232),
.B2(n_2224),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2482),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2427),
.A2(n_2240),
.B1(n_2241),
.B2(n_2235),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2543),
.B(n_2194),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2543),
.B(n_2423),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2426),
.B(n_1559),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_L g2714 ( 
.A(n_2427),
.B(n_2186),
.C(n_2184),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2397),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2494),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2523),
.B(n_2536),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2497),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2416),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2523),
.B(n_2230),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_L g2721 ( 
.A(n_2429),
.B(n_1564),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2498),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2388),
.B(n_1565),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_SL g2724 ( 
.A(n_2581),
.B(n_2216),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2323),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2501),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2559),
.B(n_2216),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2536),
.B(n_2230),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2334),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2388),
.B(n_2546),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2559),
.B(n_2216),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2387),
.B(n_2190),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2503),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_SL g2734 ( 
.A(n_2360),
.B(n_2311),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2345),
.B(n_1565),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2345),
.B(n_1579),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2425),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2436),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2438),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2514),
.Y(n_2740)
);

BUFx8_ASAP7_75t_L g2741 ( 
.A(n_2339),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_2371),
.B(n_1579),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2516),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2521),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_SL g2745 ( 
.A(n_2391),
.B(n_2216),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_L g2746 ( 
.A(n_2371),
.B(n_1586),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2549),
.B(n_2228),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2385),
.B(n_2088),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_2417),
.B(n_1586),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2441),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2483),
.B(n_1608),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2546),
.B(n_2233),
.Y(n_2752)
);

INVx2_ASAP7_75t_SL g2753 ( 
.A(n_2318),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2326),
.B(n_2233),
.Y(n_2754)
);

NOR2xp67_ASAP7_75t_L g2755 ( 
.A(n_2554),
.B(n_2192),
.Y(n_2755)
);

INVxp67_ASAP7_75t_L g2756 ( 
.A(n_2357),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2520),
.B(n_1608),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2326),
.B(n_2237),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2549),
.B(n_2228),
.Y(n_2759)
);

INVx2_ASAP7_75t_SL g2760 ( 
.A(n_2337),
.Y(n_2760)
);

NOR3xp33_ASAP7_75t_L g2761 ( 
.A(n_2363),
.B(n_2227),
.C(n_2222),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2385),
.B(n_2237),
.Y(n_2762)
);

INVxp33_ASAP7_75t_L g2763 ( 
.A(n_2349),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2524),
.Y(n_2764)
);

NOR3xp33_ASAP7_75t_L g2765 ( 
.A(n_2363),
.B(n_2227),
.C(n_2222),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2528),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2671),
.B(n_2238),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2585),
.B(n_2228),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2671),
.B(n_2238),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2317),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2540),
.B(n_2362),
.C(n_2542),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2506),
.B(n_2239),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2319),
.Y(n_2773)
);

NOR2xp67_ASAP7_75t_L g2774 ( 
.A(n_2629),
.B(n_2239),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2557),
.B(n_1613),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2506),
.B(n_2245),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2324),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2510),
.B(n_2245),
.Y(n_2778)
);

NOR2xp67_ASAP7_75t_L g2779 ( 
.A(n_2629),
.B(n_2248),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2557),
.B(n_1613),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2334),
.Y(n_2781)
);

INVx8_ASAP7_75t_L g2782 ( 
.A(n_2491),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2551),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2333),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2340),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2510),
.B(n_2248),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2574),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2331),
.B(n_2251),
.Y(n_2788)
);

NOR2xp67_ASAP7_75t_L g2789 ( 
.A(n_2407),
.B(n_2251),
.Y(n_2789)
);

NAND2xp33_ASAP7_75t_L g2790 ( 
.A(n_2597),
.B(n_2228),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2380),
.B(n_1626),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2585),
.B(n_2236),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2512),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2331),
.B(n_2249),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2434),
.B(n_2249),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2396),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2344),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2434),
.B(n_2252),
.Y(n_2798)
);

NOR3xp33_ASAP7_75t_L g2799 ( 
.A(n_2355),
.B(n_2254),
.C(n_2252),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2352),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2442),
.B(n_2254),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2577),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2354),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2396),
.B(n_1626),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2485),
.B(n_1628),
.Y(n_2805)
);

INVxp33_ASAP7_75t_L g2806 ( 
.A(n_2466),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2370),
.Y(n_2807)
);

NAND2xp33_ASAP7_75t_L g2808 ( 
.A(n_2597),
.B(n_2236),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2496),
.B(n_1628),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2375),
.Y(n_2810)
);

BUFx5_ASAP7_75t_L g2811 ( 
.A(n_2447),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2491),
.Y(n_2812)
);

BUFx8_ASAP7_75t_L g2813 ( 
.A(n_2339),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2583),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2377),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2382),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2464),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2442),
.B(n_2243),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2454),
.B(n_2255),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2508),
.B(n_2236),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2592),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2595),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2454),
.B(n_2256),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2461),
.B(n_2257),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_SL g2825 ( 
.A(n_2391),
.B(n_2236),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2461),
.B(n_2561),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2561),
.B(n_2261),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2477),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2599),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2435),
.B(n_2246),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2620),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2496),
.B(n_1634),
.Y(n_2832)
);

AND2x6_ASAP7_75t_SL g2833 ( 
.A(n_2649),
.B(n_1634),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2632),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2479),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2563),
.B(n_2263),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_SL g2837 ( 
.A(n_2541),
.B(n_2246),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2639),
.Y(n_2838)
);

BUFx6f_ASAP7_75t_L g2839 ( 
.A(n_2334),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2486),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2563),
.B(n_2264),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2435),
.B(n_2246),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2591),
.B(n_2246),
.Y(n_2843)
);

NOR2xp67_ASAP7_75t_L g2844 ( 
.A(n_2505),
.B(n_2279),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_L g2845 ( 
.A(n_2356),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2489),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2637),
.B(n_1635),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2591),
.B(n_2247),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2646),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2493),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2511),
.B(n_2247),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2495),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2507),
.Y(n_2853)
);

INVxp33_ASAP7_75t_L g2854 ( 
.A(n_2628),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2320),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2513),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2588),
.B(n_2247),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2449),
.B(n_2247),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2449),
.B(n_2250),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2527),
.B(n_2250),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2428),
.B(n_1635),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2588),
.B(n_2250),
.Y(n_2862)
);

NOR3xp33_ASAP7_75t_L g2863 ( 
.A(n_2607),
.B(n_2362),
.C(n_2529),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2575),
.B(n_1636),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2518),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2612),
.B(n_1636),
.Y(n_2866)
);

NAND3xp33_ASAP7_75t_L g2867 ( 
.A(n_2540),
.B(n_2139),
.C(n_2185),
.Y(n_2867)
);

BUFx6f_ASAP7_75t_L g2868 ( 
.A(n_2356),
.Y(n_2868)
);

AOI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2358),
.A2(n_2259),
.B1(n_2265),
.B2(n_2250),
.Y(n_2869)
);

A2O1A1Ixp33_ASAP7_75t_L g2870 ( 
.A1(n_2451),
.A2(n_2021),
.B(n_2018),
.C(n_2014),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2468),
.B(n_2265),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2322),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2373),
.B(n_1657),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2502),
.B(n_2265),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2608),
.B(n_2265),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2502),
.B(n_2304),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2611),
.B(n_2304),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2617),
.B(n_2624),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2538),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2643),
.B(n_2026),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2539),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2527),
.B(n_2282),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2547),
.B(n_2035),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2548),
.B(n_2055),
.Y(n_2884)
);

A2O1A1Ixp33_ASAP7_75t_L g2885 ( 
.A1(n_2542),
.A2(n_2143),
.B(n_2023),
.C(n_2076),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2328),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2357),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2550),
.B(n_2023),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2373),
.B(n_2517),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2532),
.B(n_2282),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2558),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2562),
.B(n_2068),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2509),
.B(n_2282),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_2544),
.B(n_2283),
.Y(n_2894)
);

NAND2x1_ASAP7_75t_L g2895 ( 
.A(n_2418),
.B(n_2010),
.Y(n_2895)
);

AO221x1_ASAP7_75t_L g2896 ( 
.A1(n_2445),
.A2(n_2010),
.B1(n_2031),
.B2(n_2024),
.C(n_2291),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2419),
.B(n_1657),
.Y(n_2897)
);

INVx2_ASAP7_75t_SL g2898 ( 
.A(n_2419),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2338),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2578),
.B(n_2068),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2499),
.B(n_1661),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2499),
.B(n_1661),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2603),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_L g2904 ( 
.A(n_2500),
.B(n_1674),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2544),
.B(n_2301),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2606),
.Y(n_2906)
);

NAND3xp33_ASAP7_75t_L g2907 ( 
.A(n_2515),
.B(n_2185),
.C(n_2214),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2346),
.B(n_2068),
.Y(n_2908)
);

AND2x6_ASAP7_75t_L g2909 ( 
.A(n_2654),
.B(n_2269),
.Y(n_2909)
);

INVx3_ASAP7_75t_L g2910 ( 
.A(n_2491),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2342),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2348),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2350),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2346),
.B(n_2077),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2351),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2364),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_SL g2917 ( 
.A(n_2545),
.B(n_1676),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2347),
.B(n_2077),
.Y(n_2918)
);

NOR2xp67_ASAP7_75t_L g2919 ( 
.A(n_2601),
.B(n_2258),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2366),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2374),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2347),
.B(n_2077),
.Y(n_2922)
);

CKINVDCx20_ASAP7_75t_R g2923 ( 
.A(n_2332),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2376),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_SL g2925 ( 
.A(n_2545),
.B(n_1676),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2566),
.B(n_2301),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2596),
.B(n_2301),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2381),
.Y(n_2928)
);

INVxp67_ASAP7_75t_L g2929 ( 
.A(n_2500),
.Y(n_2929)
);

INVxp67_ASAP7_75t_L g2930 ( 
.A(n_2530),
.Y(n_2930)
);

NAND2xp33_ASAP7_75t_L g2931 ( 
.A(n_2597),
.B(n_2411),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2447),
.B(n_2062),
.Y(n_2932)
);

NOR2xp67_ASAP7_75t_L g2933 ( 
.A(n_2576),
.B(n_2280),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2392),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2394),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2399),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2401),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2414),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_2321),
.B(n_2443),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2661),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2343),
.Y(n_2941)
);

INVx2_ASAP7_75t_SL g2942 ( 
.A(n_2365),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2321),
.B(n_2283),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2361),
.B(n_1674),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2647),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2665),
.Y(n_2946)
);

NAND2xp33_ASAP7_75t_L g2947 ( 
.A(n_2411),
.B(n_2283),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2668),
.Y(n_2948)
);

BUFx3_ASAP7_75t_L g2949 ( 
.A(n_2403),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2447),
.B(n_2065),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2321),
.B(n_2283),
.Y(n_2951)
);

NAND2xp33_ASAP7_75t_SL g2952 ( 
.A(n_2641),
.B(n_1682),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2321),
.B(n_2301),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2669),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2555),
.B(n_2065),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2555),
.B(n_2098),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2439),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2648),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2406),
.B(n_2098),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2650),
.Y(n_2960)
);

BUFx6f_ASAP7_75t_L g2961 ( 
.A(n_2356),
.Y(n_2961)
);

NOR2xp67_ASAP7_75t_L g2962 ( 
.A(n_2450),
.B(n_2286),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2670),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2361),
.B(n_1691),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2796),
.B(n_2341),
.Y(n_2965)
);

AND2x6_ASAP7_75t_SL g2966 ( 
.A(n_2804),
.B(n_2735),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2682),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2916),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_SL g2969 ( 
.A(n_2723),
.B(n_2341),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2690),
.B(n_2605),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2717),
.B(n_2445),
.Y(n_2971)
);

NAND2xp33_ASAP7_75t_L g2972 ( 
.A(n_2771),
.B(n_2602),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2730),
.B(n_2445),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2676),
.B(n_2677),
.Y(n_2974)
);

INVx2_ASAP7_75t_SL g2975 ( 
.A(n_2715),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2685),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2949),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2689),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2699),
.B(n_2415),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2789),
.B(n_2594),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2713),
.B(n_1691),
.Y(n_2981)
);

OAI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2771),
.A2(n_2619),
.B(n_2634),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2692),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2706),
.Y(n_2984)
);

INVxp67_ASAP7_75t_L g2985 ( 
.A(n_2864),
.Y(n_2985)
);

BUFx8_ASAP7_75t_L g2986 ( 
.A(n_2793),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2707),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2754),
.B(n_2422),
.Y(n_2988)
);

AOI22xp33_ASAP7_75t_L g2989 ( 
.A1(n_2863),
.A2(n_2410),
.B1(n_2390),
.B2(n_2480),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2936),
.Y(n_2990)
);

OR2x6_ASAP7_75t_L g2991 ( 
.A(n_2782),
.B(n_2492),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2673),
.A2(n_2410),
.B1(n_2390),
.B2(n_2480),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2758),
.B(n_2437),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2709),
.Y(n_2994)
);

INVx8_ASAP7_75t_L g2995 ( 
.A(n_2782),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2826),
.B(n_2325),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2805),
.B(n_2530),
.Y(n_2997)
);

OAI221xp5_ASAP7_75t_L g2998 ( 
.A1(n_2809),
.A2(n_2604),
.B1(n_2832),
.B2(n_2847),
.C(n_2721),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2672),
.A2(n_2714),
.B1(n_2638),
.B2(n_2742),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2732),
.B(n_2720),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2866),
.B(n_2746),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2716),
.Y(n_3002)
);

AO22x1_ASAP7_75t_L g3003 ( 
.A1(n_2889),
.A2(n_2409),
.B1(n_2616),
.B2(n_2405),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2755),
.B(n_2623),
.Y(n_3004)
);

NOR2xp67_ASAP7_75t_SL g3005 ( 
.A(n_2812),
.B(n_2525),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2917),
.B(n_2623),
.Y(n_3006)
);

INVx4_ASAP7_75t_L g3007 ( 
.A(n_2782),
.Y(n_3007)
);

NAND2x1p5_ASAP7_75t_L g3008 ( 
.A(n_2812),
.B(n_2406),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2718),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2728),
.B(n_2327),
.Y(n_3010)
);

INVx2_ASAP7_75t_SL g3011 ( 
.A(n_2697),
.Y(n_3011)
);

INVxp67_ASAP7_75t_SL g3012 ( 
.A(n_2756),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2722),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2775),
.B(n_2780),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_2683),
.A2(n_2616),
.B1(n_2598),
.B2(n_2471),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2678),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2917),
.B(n_2645),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2944),
.A2(n_2487),
.B1(n_2571),
.B2(n_2567),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2726),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2858),
.A2(n_2625),
.B1(n_2586),
.B2(n_2645),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2854),
.B(n_2613),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2788),
.B(n_2626),
.Y(n_3022)
);

CKINVDCx6p67_ASAP7_75t_R g3023 ( 
.A(n_2923),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2791),
.A2(n_2457),
.B1(n_2607),
.B2(n_2402),
.Y(n_3024)
);

O2A1O1Ixp5_ASAP7_75t_L g3025 ( 
.A1(n_2674),
.A2(n_2460),
.B(n_2467),
.C(n_2458),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2733),
.Y(n_3026)
);

AND2x4_ASAP7_75t_L g3027 ( 
.A(n_2860),
.B(n_2456),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2925),
.B(n_2657),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2763),
.B(n_2964),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_2736),
.B(n_2444),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2700),
.B(n_2586),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2767),
.B(n_2446),
.Y(n_3032)
);

NAND2xp33_ASAP7_75t_L g3033 ( 
.A(n_2704),
.B(n_2602),
.Y(n_3033)
);

AOI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2751),
.A2(n_2757),
.B1(n_2749),
.B2(n_2861),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2897),
.B(n_1703),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2740),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2769),
.B(n_2448),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2859),
.A2(n_2625),
.B1(n_2406),
.B2(n_2443),
.Y(n_3038)
);

AO22x1_ASAP7_75t_L g3039 ( 
.A1(n_2806),
.A2(n_2618),
.B1(n_2602),
.B2(n_2330),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2860),
.B(n_2492),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2712),
.B(n_2372),
.Y(n_3041)
);

NOR3xp33_ASAP7_75t_SL g3042 ( 
.A(n_2873),
.B(n_2424),
.C(n_2615),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2933),
.B(n_2492),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2794),
.B(n_2752),
.Y(n_3044)
);

O2A1O1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_2691),
.A2(n_2660),
.B(n_2384),
.C(n_2395),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_SL g3046 ( 
.A(n_2925),
.B(n_2657),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_2761),
.A2(n_2642),
.B1(n_2393),
.B2(n_2440),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2743),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2744),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2745),
.A2(n_2443),
.B(n_2406),
.Y(n_3050)
);

NOR2x2_ASAP7_75t_L g3051 ( 
.A(n_2945),
.B(n_2649),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2772),
.B(n_2431),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2901),
.B(n_1703),
.Y(n_3053)
);

AOI22xp33_ASAP7_75t_L g3054 ( 
.A1(n_2765),
.A2(n_2644),
.B1(n_2472),
.B2(n_2359),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2776),
.B(n_2469),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2680),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2734),
.A2(n_2472),
.B1(n_2359),
.B2(n_2476),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2902),
.B(n_2630),
.Y(n_3058)
);

BUFx6f_ASAP7_75t_L g3059 ( 
.A(n_2688),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2741),
.Y(n_3060)
);

AOI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_2734),
.A2(n_2481),
.B1(n_2522),
.B2(n_2488),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_L g3062 ( 
.A(n_2904),
.B(n_2618),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2694),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_SL g3064 ( 
.A1(n_2696),
.A2(n_2610),
.B1(n_2649),
.B2(n_2537),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2778),
.B(n_2579),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2786),
.B(n_2568),
.Y(n_3066)
);

OR2x2_ASAP7_75t_L g3067 ( 
.A(n_2887),
.B(n_2610),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2818),
.B(n_2584),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2702),
.B(n_2590),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2764),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2705),
.B(n_2329),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2766),
.B(n_2452),
.Y(n_3072)
);

INVx2_ASAP7_75t_SL g3073 ( 
.A(n_2941),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2783),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2787),
.B(n_2619),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2701),
.B(n_2330),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2952),
.A2(n_2589),
.B1(n_2610),
.B2(n_2602),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2802),
.B(n_2335),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2929),
.B(n_2652),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2679),
.A2(n_2335),
.B1(n_2552),
.B2(n_2411),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2814),
.B(n_2573),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2898),
.B(n_2484),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2821),
.Y(n_3083)
);

AND2x4_ASAP7_75t_L g3084 ( 
.A(n_2942),
.B(n_2656),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2822),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2753),
.B(n_2760),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2930),
.B(n_2635),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2829),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2741),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2745),
.A2(n_2443),
.B(n_2553),
.Y(n_3090)
);

OR2x2_ASAP7_75t_L g3091 ( 
.A(n_2878),
.B(n_2565),
.Y(n_3091)
);

NAND2xp33_ASAP7_75t_L g3092 ( 
.A(n_2704),
.B(n_2411),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2831),
.Y(n_3093)
);

BUFx8_ASAP7_75t_L g3094 ( 
.A(n_2688),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2834),
.B(n_2573),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_SL g3096 ( 
.A1(n_2838),
.A2(n_2635),
.B1(n_2565),
.B2(n_2504),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_2813),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2849),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2695),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2819),
.B(n_2526),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2724),
.B(n_2635),
.Y(n_3101)
);

O2A1O1Ixp5_ASAP7_75t_L g3102 ( 
.A1(n_2820),
.A2(n_2634),
.B(n_2663),
.C(n_2260),
.Y(n_3102)
);

INVx5_ASAP7_75t_L g3103 ( 
.A(n_2845),
.Y(n_3103)
);

AOI221xp5_ASAP7_75t_L g3104 ( 
.A1(n_2855),
.A2(n_2526),
.B1(n_2664),
.B2(n_2299),
.C(n_2290),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2872),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2886),
.B(n_2552),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2899),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2911),
.B(n_2552),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2912),
.B(n_2552),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2913),
.B(n_2656),
.Y(n_3110)
);

BUFx2_ASAP7_75t_L g3111 ( 
.A(n_2688),
.Y(n_3111)
);

AND2x6_ASAP7_75t_SL g3112 ( 
.A(n_2813),
.B(n_2664),
.Y(n_3112)
);

NAND3xp33_ASAP7_75t_L g3113 ( 
.A(n_2684),
.B(n_2033),
.C(n_2631),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2693),
.B(n_2484),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2693),
.B(n_2490),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2915),
.B(n_2920),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2957),
.A2(n_2622),
.B1(n_2369),
.B2(n_2379),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2703),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2693),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2921),
.B(n_2474),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2725),
.B(n_2490),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2924),
.B(n_2928),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2934),
.B(n_2474),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_2725),
.B(n_2525),
.Y(n_3124)
);

INVx2_ASAP7_75t_SL g3125 ( 
.A(n_2725),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2935),
.B(n_2937),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2938),
.B(n_2474),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2825),
.A2(n_2569),
.B(n_2553),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2940),
.B(n_2823),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2946),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_2896),
.A2(n_2622),
.B1(n_2369),
.B2(n_2379),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2824),
.B(n_2353),
.Y(n_3132)
);

AND2x6_ASAP7_75t_SL g3133 ( 
.A(n_2833),
.B(n_2288),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2948),
.B(n_2353),
.Y(n_3134)
);

CKINVDCx5p33_ASAP7_75t_R g3135 ( 
.A(n_2833),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_2729),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2954),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2880),
.B(n_2389),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2927),
.A2(n_2622),
.B1(n_2421),
.B2(n_2432),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_SL g3140 ( 
.A(n_2825),
.B(n_2525),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2795),
.B(n_2389),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2729),
.B(n_2525),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2729),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2798),
.B(n_2421),
.Y(n_3144)
);

AOI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2919),
.A2(n_2622),
.B1(n_2662),
.B2(n_2659),
.Y(n_3145)
);

INVx2_ASAP7_75t_SL g3146 ( 
.A(n_2781),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2719),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2801),
.B(n_2432),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_R g3149 ( 
.A(n_2910),
.B(n_2666),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2958),
.A2(n_2459),
.B1(n_2533),
.B2(n_2433),
.Y(n_3150)
);

O2A1O1Ixp5_ASAP7_75t_L g3151 ( 
.A1(n_2837),
.A2(n_2663),
.B(n_2667),
.C(n_2655),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2827),
.B(n_2433),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2737),
.Y(n_3153)
);

HB1xp67_ASAP7_75t_L g3154 ( 
.A(n_2781),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2675),
.B(n_2459),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_SL g3156 ( 
.A(n_2781),
.B(n_2553),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2839),
.B(n_2553),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_SL g3158 ( 
.A(n_2839),
.B(n_2569),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_2839),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_2845),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2738),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2836),
.B(n_2533),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2841),
.B(n_2534),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2960),
.B(n_2534),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2962),
.B(n_2569),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2883),
.B(n_2564),
.Y(n_3166)
);

NAND2xp33_ASAP7_75t_L g3167 ( 
.A(n_2704),
.B(n_2367),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2883),
.B(n_2564),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2884),
.B(n_2572),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_2708),
.B(n_2569),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2884),
.B(n_2572),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2955),
.B(n_2614),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_2963),
.B(n_2614),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2739),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2956),
.B(n_2876),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2877),
.B(n_2627),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2686),
.B(n_2587),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2843),
.B(n_2627),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2848),
.B(n_2633),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_SL g3180 ( 
.A(n_2845),
.B(n_2587),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_2747),
.A2(n_2662),
.B1(n_2666),
.B2(n_2659),
.Y(n_3181)
);

OR2x6_ASAP7_75t_L g3182 ( 
.A(n_2910),
.B(n_2367),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2770),
.B(n_2633),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2750),
.Y(n_3184)
);

A2O1A1Ixp33_ASAP7_75t_L g3185 ( 
.A1(n_2844),
.A2(n_2907),
.B(n_2867),
.C(n_2871),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2879),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2881),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_2868),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2974),
.B(n_2773),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3140),
.A2(n_2947),
.B(n_2790),
.Y(n_3190)
);

INVx2_ASAP7_75t_SL g3191 ( 
.A(n_2986),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3014),
.B(n_2777),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2968),
.Y(n_3193)
);

INVx2_ASAP7_75t_SL g3194 ( 
.A(n_2986),
.Y(n_3194)
);

BUFx8_ASAP7_75t_L g3195 ( 
.A(n_3060),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2990),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2998),
.B(n_2687),
.Y(n_3197)
);

CKINVDCx8_ASAP7_75t_R g3198 ( 
.A(n_3112),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3000),
.B(n_2784),
.Y(n_3199)
);

BUFx6f_ASAP7_75t_L g3200 ( 
.A(n_3103),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_3140),
.A2(n_2808),
.B(n_2681),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2997),
.B(n_2903),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2992),
.A2(n_2989),
.B1(n_2999),
.B2(n_3024),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_3006),
.A2(n_2907),
.B1(n_2799),
.B2(n_2851),
.Y(n_3204)
);

NOR2x2_ASAP7_75t_L g3205 ( 
.A(n_3182),
.B(n_2785),
.Y(n_3205)
);

INVx2_ASAP7_75t_SL g3206 ( 
.A(n_2977),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2970),
.B(n_2797),
.Y(n_3207)
);

O2A1O1Ixp33_ASAP7_75t_L g3208 ( 
.A1(n_3017),
.A2(n_2874),
.B(n_2905),
.C(n_2894),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3001),
.B(n_2985),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_3045),
.A2(n_2779),
.B(n_2774),
.C(n_2710),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2981),
.B(n_2759),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_3030),
.B(n_3034),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_3103),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2979),
.B(n_2800),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_3050),
.A2(n_2870),
.B(n_2931),
.Y(n_3215)
);

O2A1O1Ixp33_ASAP7_75t_SL g3216 ( 
.A1(n_3004),
.A2(n_2973),
.B(n_2971),
.C(n_2969),
.Y(n_3216)
);

OA21x2_ASAP7_75t_L g3217 ( 
.A1(n_3113),
.A2(n_2070),
.B(n_2885),
.Y(n_3217)
);

CKINVDCx20_ASAP7_75t_R g3218 ( 
.A(n_3023),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2988),
.B(n_2803),
.Y(n_3219)
);

INVx2_ASAP7_75t_SL g3220 ( 
.A(n_2975),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3021),
.B(n_3042),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_3092),
.A2(n_3033),
.B(n_3090),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2993),
.B(n_2807),
.Y(n_3223)
);

AND2x2_ASAP7_75t_SL g3224 ( 
.A(n_2972),
.B(n_2875),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_3029),
.B(n_2906),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_3047),
.A2(n_2869),
.B1(n_2711),
.B2(n_2792),
.Y(n_3226)
);

A2O1A1Ixp33_ASAP7_75t_L g3227 ( 
.A1(n_3185),
.A2(n_2684),
.B(n_2867),
.C(n_2731),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3128),
.A2(n_2748),
.B(n_2587),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_3062),
.B(n_2926),
.Y(n_3229)
);

OAI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_3025),
.A2(n_2727),
.B(n_2893),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_3035),
.B(n_2704),
.Y(n_3231)
);

AND2x4_ASAP7_75t_L g3232 ( 
.A(n_3040),
.B(n_2768),
.Y(n_3232)
);

BUFx2_ASAP7_75t_L g3233 ( 
.A(n_3159),
.Y(n_3233)
);

NAND2xp33_ASAP7_75t_L g3234 ( 
.A(n_2995),
.B(n_2704),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3167),
.A2(n_2748),
.B(n_2587),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3032),
.B(n_2810),
.Y(n_3236)
);

BUFx2_ASAP7_75t_L g3237 ( 
.A(n_3188),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3044),
.A2(n_2939),
.B(n_2842),
.Y(n_3238)
);

OR2x2_ASAP7_75t_L g3239 ( 
.A(n_3116),
.B(n_2815),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3037),
.B(n_2816),
.Y(n_3240)
);

NOR2x1p5_ASAP7_75t_SL g3241 ( 
.A(n_3091),
.B(n_2811),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3016),
.Y(n_3242)
);

INVx1_ASAP7_75t_SL g3243 ( 
.A(n_3011),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3027),
.B(n_2817),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3071),
.A2(n_2842),
.B(n_2830),
.Y(n_3245)
);

NOR2x1_ASAP7_75t_R g3246 ( 
.A(n_3089),
.B(n_2961),
.Y(n_3246)
);

INVx2_ASAP7_75t_SL g3247 ( 
.A(n_3094),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_SL g3248 ( 
.A(n_3007),
.B(n_2418),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3031),
.A2(n_2830),
.B(n_2762),
.Y(n_3249)
);

BUFx2_ASAP7_75t_L g3250 ( 
.A(n_3094),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3022),
.B(n_2828),
.Y(n_3251)
);

OAI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3175),
.A2(n_2890),
.B(n_2698),
.Y(n_3252)
);

NAND2x1p5_ASAP7_75t_L g3253 ( 
.A(n_3007),
.B(n_2868),
.Y(n_3253)
);

O2A1O1Ixp33_ASAP7_75t_L g3254 ( 
.A1(n_3028),
.A2(n_2862),
.B(n_2857),
.C(n_2882),
.Y(n_3254)
);

OAI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_2996),
.A2(n_2950),
.B(n_2932),
.Y(n_3255)
);

AOI21x1_ASAP7_75t_L g3256 ( 
.A1(n_3177),
.A2(n_2914),
.B(n_2908),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3129),
.B(n_2835),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2973),
.B(n_2840),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3010),
.B(n_2846),
.Y(n_3259)
);

OR2x6_ASAP7_75t_L g3260 ( 
.A(n_2995),
.B(n_2868),
.Y(n_3260)
);

AOI21x1_ASAP7_75t_L g3261 ( 
.A1(n_3170),
.A2(n_2914),
.B(n_2908),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3056),
.Y(n_3262)
);

AOI21xp33_ASAP7_75t_L g3263 ( 
.A1(n_3053),
.A2(n_2950),
.B(n_2932),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_3058),
.B(n_2850),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_3068),
.B(n_2852),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3122),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3126),
.Y(n_3267)
);

O2A1O1Ixp33_ASAP7_75t_L g3268 ( 
.A1(n_3046),
.A2(n_2959),
.B(n_2853),
.C(n_2865),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3063),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3052),
.B(n_2856),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2967),
.Y(n_3271)
);

NAND2xp33_ASAP7_75t_L g3272 ( 
.A(n_2995),
.B(n_2811),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3113),
.A2(n_2888),
.B(n_2918),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_SL g3274 ( 
.A(n_3057),
.B(n_2811),
.Y(n_3274)
);

OAI22xp5_ASAP7_75t_SL g3275 ( 
.A1(n_3135),
.A2(n_2961),
.B1(n_2895),
.B2(n_2891),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2976),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_3103),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3027),
.B(n_2961),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_SL g3279 ( 
.A(n_3041),
.B(n_2811),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_2982),
.A2(n_2888),
.B(n_2918),
.Y(n_3280)
);

A2O1A1Ixp33_ASAP7_75t_L g3281 ( 
.A1(n_3015),
.A2(n_2640),
.B(n_2951),
.C(n_2943),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2982),
.A2(n_2922),
.B(n_2900),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_2980),
.B(n_2811),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3012),
.B(n_2922),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_3073),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3100),
.A2(n_2900),
.B(n_2892),
.Y(n_3286)
);

O2A1O1Ixp33_ASAP7_75t_L g3287 ( 
.A1(n_2965),
.A2(n_2953),
.B(n_2640),
.C(n_2315),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_3100),
.A2(n_2892),
.B(n_2593),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3038),
.A2(n_2593),
.B(n_2504),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3075),
.B(n_2367),
.Y(n_3290)
);

AOI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3054),
.A2(n_2909),
.B1(n_2653),
.B2(n_2658),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3099),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_3038),
.A2(n_2653),
.B(n_2651),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2966),
.B(n_2531),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3118),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_3008),
.Y(n_3296)
);

INVxp67_ASAP7_75t_L g3297 ( 
.A(n_3086),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3161),
.Y(n_3298)
);

OR2x6_ASAP7_75t_SL g3299 ( 
.A(n_3110),
.B(n_2269),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3055),
.B(n_3065),
.Y(n_3300)
);

O2A1O1Ixp5_ASAP7_75t_L g3301 ( 
.A1(n_3039),
.A2(n_2658),
.B(n_2651),
.C(n_2031),
.Y(n_3301)
);

INVxp67_ASAP7_75t_L g3302 ( 
.A(n_3087),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3102),
.A2(n_2580),
.B(n_2531),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3066),
.A2(n_2580),
.B(n_2531),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3069),
.A2(n_2582),
.B(n_2580),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3020),
.A2(n_2609),
.B(n_2582),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_3020),
.A2(n_2609),
.B(n_2582),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_3079),
.B(n_2609),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3081),
.B(n_2621),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_3172),
.A2(n_2024),
.B(n_2033),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3095),
.B(n_2621),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3040),
.B(n_2978),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3174),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_3003),
.B(n_2621),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_3103),
.Y(n_3315)
);

AOI21x1_ASAP7_75t_L g3316 ( 
.A1(n_3132),
.A2(n_2033),
.B(n_2271),
.Y(n_3316)
);

AND2x2_ASAP7_75t_SL g3317 ( 
.A(n_3061),
.B(n_2636),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_3138),
.A2(n_2636),
.B(n_2272),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_2980),
.B(n_2636),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2983),
.Y(n_3320)
);

AND2x4_ASAP7_75t_L g3321 ( 
.A(n_3043),
.B(n_2271),
.Y(n_3321)
);

OR2x6_ASAP7_75t_L g3322 ( 
.A(n_2991),
.B(n_2272),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3184),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2984),
.B(n_2909),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3096),
.A2(n_2289),
.B(n_2287),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_3166),
.A2(n_2289),
.B(n_2287),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_L g3327 ( 
.A(n_3059),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2987),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2994),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3018),
.A2(n_2909),
.B1(n_2291),
.B2(n_1295),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3168),
.A2(n_2909),
.B(n_1295),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_3067),
.B(n_545),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3002),
.B(n_2),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3009),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3169),
.A2(n_1295),
.B(n_1252),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3013),
.B(n_3),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_3101),
.B(n_547),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3019),
.B(n_5),
.Y(n_3338)
);

CKINVDCx5p33_ASAP7_75t_R g3339 ( 
.A(n_3097),
.Y(n_3339)
);

A2O1A1Ixp33_ASAP7_75t_L g3340 ( 
.A1(n_3077),
.A2(n_1295),
.B(n_1252),
.C(n_7),
.Y(n_3340)
);

OAI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3072),
.A2(n_1731),
.B(n_5),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3026),
.B(n_6),
.Y(n_3342)
);

HB1xp67_ASAP7_75t_L g3343 ( 
.A(n_3154),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3036),
.B(n_6),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3008),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3171),
.A2(n_1252),
.B(n_549),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3147),
.B(n_7),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3048),
.Y(n_3348)
);

O2A1O1Ixp5_ASAP7_75t_L g3349 ( 
.A1(n_3165),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_3151),
.A2(n_1252),
.B(n_685),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3049),
.B(n_9),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3078),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_3352)
);

OAI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3155),
.A2(n_11),
.B(n_12),
.Y(n_3353)
);

O2A1O1Ixp33_ASAP7_75t_L g3354 ( 
.A1(n_3076),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_3354)
);

O2A1O1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_3114),
.A2(n_17),
.B(n_14),
.C(n_15),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3070),
.B(n_17),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3152),
.A2(n_698),
.B(n_696),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_3059),
.Y(n_3358)
);

HB1xp67_ASAP7_75t_L g3359 ( 
.A(n_3111),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3162),
.A2(n_700),
.B(n_550),
.Y(n_3360)
);

OAI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3141),
.A2(n_19),
.B(n_20),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3074),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3083),
.B(n_3085),
.Y(n_3363)
);

OAI21x1_ASAP7_75t_L g3364 ( 
.A1(n_3144),
.A2(n_551),
.B(n_548),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3088),
.B(n_19),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3139),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3163),
.A2(n_683),
.B(n_682),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_3059),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3093),
.Y(n_3369)
);

AND2x4_ASAP7_75t_L g3370 ( 
.A(n_3043),
.B(n_553),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3098),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_R g3372 ( 
.A(n_3133),
.B(n_555),
.Y(n_3372)
);

BUFx6f_ASAP7_75t_L g3373 ( 
.A(n_3136),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3124),
.A2(n_689),
.B(n_688),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3105),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3107),
.Y(n_3376)
);

NOR2xp67_ASAP7_75t_L g3377 ( 
.A(n_3153),
.B(n_556),
.Y(n_3377)
);

OAI21xp33_ASAP7_75t_L g3378 ( 
.A1(n_3130),
.A2(n_21),
.B(n_23),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_3119),
.Y(n_3379)
);

AOI22x1_ASAP7_75t_L g3380 ( 
.A1(n_3137),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3187),
.B(n_28),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_3082),
.B(n_557),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3186),
.B(n_28),
.Y(n_3383)
);

HB1xp67_ASAP7_75t_L g3384 ( 
.A(n_3160),
.Y(n_3384)
);

AND2x4_ASAP7_75t_L g3385 ( 
.A(n_2991),
.B(n_559),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_3142),
.A2(n_3148),
.B(n_3176),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_3115),
.B(n_560),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3178),
.A2(n_672),
.B(n_670),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3084),
.B(n_30),
.Y(n_3389)
);

BUFx6f_ASAP7_75t_L g3390 ( 
.A(n_3136),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3134),
.B(n_30),
.Y(n_3391)
);

OAI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3173),
.A2(n_31),
.B(n_32),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3179),
.B(n_31),
.Y(n_3393)
);

OAI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3106),
.A2(n_32),
.B(n_34),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3164),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3183),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3125),
.B(n_34),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3143),
.B(n_35),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3300),
.B(n_3121),
.Y(n_3399)
);

AND2x4_ASAP7_75t_L g3400 ( 
.A(n_3385),
.B(n_2991),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3341),
.A2(n_3109),
.B(n_3108),
.Y(n_3401)
);

HB1xp67_ASAP7_75t_L g3402 ( 
.A(n_3343),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3328),
.Y(n_3403)
);

INVxp67_ASAP7_75t_L g3404 ( 
.A(n_3209),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3212),
.B(n_3146),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3329),
.Y(n_3406)
);

XOR2xp5_ASAP7_75t_L g3407 ( 
.A(n_3218),
.B(n_3064),
.Y(n_3407)
);

OA22x2_ASAP7_75t_L g3408 ( 
.A1(n_3353),
.A2(n_3084),
.B1(n_3123),
.B2(n_3120),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3266),
.B(n_3136),
.Y(n_3409)
);

BUFx4f_ASAP7_75t_L g3410 ( 
.A(n_3200),
.Y(n_3410)
);

CKINVDCx5p33_ASAP7_75t_R g3411 ( 
.A(n_3195),
.Y(n_3411)
);

INVx3_ASAP7_75t_L g3412 ( 
.A(n_3200),
.Y(n_3412)
);

BUFx3_ASAP7_75t_L g3413 ( 
.A(n_3233),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3202),
.B(n_3127),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3267),
.B(n_3104),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_SL g3416 ( 
.A1(n_3203),
.A2(n_3051),
.B1(n_3149),
.B2(n_3182),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3348),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3197),
.A2(n_3145),
.B1(n_3080),
.B2(n_3117),
.Y(n_3418)
);

AND3x1_ASAP7_75t_SL g3419 ( 
.A(n_3271),
.B(n_35),
.C(n_36),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3222),
.A2(n_3157),
.B(n_3156),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_3302),
.B(n_3158),
.Y(n_3421)
);

BUFx2_ASAP7_75t_L g3422 ( 
.A(n_3379),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3276),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3199),
.B(n_3180),
.Y(n_3424)
);

BUFx6f_ASAP7_75t_L g3425 ( 
.A(n_3200),
.Y(n_3425)
);

AND2x4_ASAP7_75t_L g3426 ( 
.A(n_3385),
.B(n_3182),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3214),
.B(n_3181),
.Y(n_3427)
);

AND3x1_ASAP7_75t_SL g3428 ( 
.A(n_3320),
.B(n_36),
.C(n_37),
.Y(n_3428)
);

BUFx2_ASAP7_75t_L g3429 ( 
.A(n_3205),
.Y(n_3429)
);

CKINVDCx20_ASAP7_75t_R g3430 ( 
.A(n_3195),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3213),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3334),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3211),
.A2(n_3131),
.B1(n_3150),
.B2(n_3005),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3362),
.Y(n_3434)
);

INVx1_ASAP7_75t_SL g3435 ( 
.A(n_3243),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3371),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3337),
.B(n_562),
.Y(n_3437)
);

BUFx6f_ASAP7_75t_L g3438 ( 
.A(n_3213),
.Y(n_3438)
);

BUFx6f_ASAP7_75t_L g3439 ( 
.A(n_3213),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3193),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3369),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3221),
.B(n_3225),
.Y(n_3442)
);

AOI221xp5_ASAP7_75t_SL g3443 ( 
.A1(n_3392),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.C(n_42),
.Y(n_3443)
);

INVx5_ASAP7_75t_L g3444 ( 
.A(n_3277),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3375),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3196),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_3277),
.Y(n_3447)
);

INVxp67_ASAP7_75t_SL g3448 ( 
.A(n_3284),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_3312),
.B(n_564),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_L g3450 ( 
.A(n_3264),
.B(n_565),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3244),
.B(n_568),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3242),
.Y(n_3452)
);

INVxp67_ASAP7_75t_L g3453 ( 
.A(n_3359),
.Y(n_3453)
);

INVx1_ASAP7_75t_SL g3454 ( 
.A(n_3237),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3251),
.B(n_38),
.Y(n_3455)
);

OAI21xp33_ASAP7_75t_SL g3456 ( 
.A1(n_3317),
.A2(n_39),
.B(n_40),
.Y(n_3456)
);

BUFx2_ASAP7_75t_L g3457 ( 
.A(n_3384),
.Y(n_3457)
);

BUFx3_ASAP7_75t_L g3458 ( 
.A(n_3250),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3262),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3376),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3232),
.B(n_569),
.Y(n_3461)
);

BUFx3_ASAP7_75t_L g3462 ( 
.A(n_3206),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3347),
.B(n_570),
.Y(n_3463)
);

BUFx2_ASAP7_75t_L g3464 ( 
.A(n_3327),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3192),
.B(n_571),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_L g3466 ( 
.A1(n_3215),
.A2(n_576),
.B(n_574),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3327),
.Y(n_3467)
);

NOR2xp67_ASAP7_75t_L g3468 ( 
.A(n_3297),
.B(n_686),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3332),
.B(n_579),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3363),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3219),
.B(n_42),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3278),
.B(n_580),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3275),
.B(n_581),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3269),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3258),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3223),
.B(n_43),
.Y(n_3476)
);

AOI22x1_ASAP7_75t_L g3477 ( 
.A1(n_3361),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3189),
.B(n_3236),
.Y(n_3478)
);

INVx3_ASAP7_75t_L g3479 ( 
.A(n_3277),
.Y(n_3479)
);

AND2x4_ASAP7_75t_L g3480 ( 
.A(n_3232),
.B(n_583),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3292),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3256),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3261),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3316),
.Y(n_3484)
);

BUFx6f_ASAP7_75t_L g3485 ( 
.A(n_3315),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3240),
.B(n_47),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3239),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3389),
.B(n_584),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3241),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3259),
.B(n_47),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3295),
.Y(n_3491)
);

OR2x6_ASAP7_75t_L g3492 ( 
.A(n_3201),
.B(n_585),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3322),
.B(n_589),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_L g3494 ( 
.A1(n_3378),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3494)
);

NOR2x1_ASAP7_75t_L g3495 ( 
.A(n_3229),
.B(n_51),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_R g3496 ( 
.A(n_3339),
.B(n_591),
.Y(n_3496)
);

INVx2_ASAP7_75t_SL g3497 ( 
.A(n_3220),
.Y(n_3497)
);

BUFx3_ASAP7_75t_L g3498 ( 
.A(n_3285),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_3224),
.B(n_593),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3327),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3227),
.Y(n_3501)
);

AOI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3294),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3382),
.B(n_595),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3282),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3257),
.B(n_54),
.Y(n_3505)
);

A2O1A1Ixp33_ASAP7_75t_L g3506 ( 
.A1(n_3340),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_3506)
);

BUFx2_ASAP7_75t_SL g3507 ( 
.A(n_3191),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3370),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3265),
.B(n_58),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3270),
.B(n_3207),
.Y(n_3510)
);

HB1xp67_ASAP7_75t_L g3511 ( 
.A(n_3324),
.Y(n_3511)
);

INVx1_ASAP7_75t_SL g3512 ( 
.A(n_3308),
.Y(n_3512)
);

OR2x2_ASAP7_75t_L g3513 ( 
.A(n_3393),
.B(n_3298),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3190),
.A2(n_597),
.B(n_596),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3395),
.B(n_58),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3321),
.B(n_599),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3280),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3396),
.B(n_59),
.Y(n_3518)
);

A2O1A1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_3210),
.A2(n_62),
.B(n_59),
.C(n_61),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3313),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3323),
.B(n_61),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3315),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3391),
.B(n_3383),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3245),
.B(n_62),
.Y(n_3524)
);

BUFx3_ASAP7_75t_L g3525 ( 
.A(n_3247),
.Y(n_3525)
);

INVx3_ASAP7_75t_L g3526 ( 
.A(n_3315),
.Y(n_3526)
);

INVx2_ASAP7_75t_SL g3527 ( 
.A(n_3358),
.Y(n_3527)
);

CKINVDCx20_ASAP7_75t_R g3528 ( 
.A(n_3198),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3333),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3321),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3336),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3370),
.B(n_600),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_3358),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_SL g3534 ( 
.A(n_3314),
.B(n_601),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3358),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3322),
.B(n_602),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3380),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3309),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3290),
.B(n_63),
.Y(n_3539)
);

A2O1A1Ixp33_ASAP7_75t_L g3540 ( 
.A1(n_3394),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_3540)
);

NOR2x1_ASAP7_75t_L g3541 ( 
.A(n_3296),
.B(n_68),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3311),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3226),
.B(n_603),
.Y(n_3543)
);

INVxp67_ASAP7_75t_L g3544 ( 
.A(n_3246),
.Y(n_3544)
);

AOI211xp5_ASAP7_75t_L g3545 ( 
.A1(n_3352),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3545)
);

INVxp67_ASAP7_75t_SL g3546 ( 
.A(n_3208),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3338),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3368),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3249),
.B(n_70),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3342),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3344),
.B(n_71),
.Y(n_3551)
);

AND2x4_ASAP7_75t_L g3552 ( 
.A(n_3283),
.B(n_606),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3351),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_3356),
.B(n_607),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_3194),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3365),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3387),
.B(n_72),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3368),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3368),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3381),
.B(n_3299),
.Y(n_3560)
);

NOR2xp67_ASAP7_75t_L g3561 ( 
.A(n_3296),
.B(n_610),
.Y(n_3561)
);

OR2x6_ASAP7_75t_L g3562 ( 
.A(n_3260),
.B(n_3253),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3216),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3319),
.B(n_611),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3373),
.Y(n_3565)
);

AND2x4_ASAP7_75t_L g3566 ( 
.A(n_3345),
.B(n_612),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3238),
.B(n_72),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3273),
.Y(n_3568)
);

OR2x2_ASAP7_75t_SL g3569 ( 
.A(n_3397),
.B(n_73),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3279),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3217),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3217),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3252),
.Y(n_3573)
);

OR2x2_ASAP7_75t_L g3574 ( 
.A(n_3231),
.B(n_73),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3398),
.B(n_3263),
.Y(n_3575)
);

INVx2_ASAP7_75t_SL g3576 ( 
.A(n_3373),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3230),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3390),
.Y(n_3578)
);

BUFx3_ASAP7_75t_L g3579 ( 
.A(n_3373),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3390),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3255),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3390),
.Y(n_3582)
);

HB1xp67_ASAP7_75t_L g3583 ( 
.A(n_3274),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3386),
.B(n_74),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3204),
.B(n_74),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3254),
.B(n_76),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3268),
.Y(n_3587)
);

OR2x2_ASAP7_75t_L g3588 ( 
.A(n_3286),
.B(n_76),
.Y(n_3588)
);

AOI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3366),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3589)
);

INVx4_ASAP7_75t_L g3590 ( 
.A(n_3260),
.Y(n_3590)
);

BUFx2_ASAP7_75t_L g3591 ( 
.A(n_3345),
.Y(n_3591)
);

INVx4_ASAP7_75t_L g3592 ( 
.A(n_3248),
.Y(n_3592)
);

AND3x1_ASAP7_75t_SL g3593 ( 
.A(n_3372),
.B(n_77),
.C(n_78),
.Y(n_3593)
);

INVxp67_ASAP7_75t_SL g3594 ( 
.A(n_3288),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3355),
.B(n_80),
.Y(n_3595)
);

AO22x1_ASAP7_75t_L g3596 ( 
.A1(n_3354),
.A2(n_3310),
.B1(n_3349),
.B2(n_3272),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3377),
.B(n_3281),
.Y(n_3597)
);

INVxp67_ASAP7_75t_SL g3598 ( 
.A(n_3304),
.Y(n_3598)
);

AND2x4_ASAP7_75t_L g3599 ( 
.A(n_3291),
.B(n_613),
.Y(n_3599)
);

CKINVDCx5p33_ASAP7_75t_R g3600 ( 
.A(n_3305),
.Y(n_3600)
);

NOR2xp67_ASAP7_75t_L g3601 ( 
.A(n_3346),
.B(n_615),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3364),
.Y(n_3602)
);

CKINVDCx5p33_ASAP7_75t_R g3603 ( 
.A(n_3374),
.Y(n_3603)
);

A2O1A1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_3357),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3306),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_SL g3606 ( 
.A(n_3360),
.B(n_618),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3330),
.B(n_619),
.Y(n_3607)
);

AOI22xp5_ASAP7_75t_L g3608 ( 
.A1(n_3543),
.A2(n_3367),
.B1(n_3388),
.B2(n_3234),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3594),
.A2(n_3228),
.B(n_3235),
.Y(n_3609)
);

BUFx3_ASAP7_75t_L g3610 ( 
.A(n_3462),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_3487),
.B(n_3307),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3423),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3403),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_SL g3614 ( 
.A(n_3603),
.B(n_3287),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3402),
.Y(n_3615)
);

HB1xp67_ASAP7_75t_L g3616 ( 
.A(n_3457),
.Y(n_3616)
);

BUFx6f_ASAP7_75t_L g3617 ( 
.A(n_3533),
.Y(n_3617)
);

INVx1_ASAP7_75t_SL g3618 ( 
.A(n_3512),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3406),
.Y(n_3619)
);

O2A1O1Ixp33_ASAP7_75t_L g3620 ( 
.A1(n_3540),
.A2(n_3331),
.B(n_3325),
.C(n_3301),
.Y(n_3620)
);

OAI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3416),
.A2(n_3293),
.B1(n_3289),
.B2(n_3303),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3432),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3434),
.Y(n_3623)
);

O2A1O1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3519),
.A2(n_3350),
.B(n_3335),
.C(n_3318),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3417),
.Y(n_3625)
);

BUFx2_ASAP7_75t_L g3626 ( 
.A(n_3422),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3436),
.Y(n_3627)
);

AOI21xp33_ASAP7_75t_L g3628 ( 
.A1(n_3575),
.A2(n_3326),
.B(n_82),
.Y(n_3628)
);

AOI21x1_ASAP7_75t_L g3629 ( 
.A1(n_3596),
.A2(n_83),
.B(n_84),
.Y(n_3629)
);

BUFx3_ASAP7_75t_L g3630 ( 
.A(n_3413),
.Y(n_3630)
);

AOI22x1_ASAP7_75t_L g3631 ( 
.A1(n_3600),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3631)
);

BUFx6f_ASAP7_75t_L g3632 ( 
.A(n_3533),
.Y(n_3632)
);

BUFx3_ASAP7_75t_L g3633 ( 
.A(n_3498),
.Y(n_3633)
);

BUFx8_ASAP7_75t_L g3634 ( 
.A(n_3464),
.Y(n_3634)
);

CKINVDCx5p33_ASAP7_75t_R g3635 ( 
.A(n_3411),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3469),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3441),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3445),
.Y(n_3638)
);

INVx1_ASAP7_75t_SL g3639 ( 
.A(n_3435),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3460),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_3528),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3481),
.Y(n_3642)
);

BUFx3_ASAP7_75t_L g3643 ( 
.A(n_3458),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3570),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3470),
.Y(n_3645)
);

CKINVDCx5p33_ASAP7_75t_R g3646 ( 
.A(n_3430),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3592),
.B(n_620),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3570),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3489),
.B(n_695),
.Y(n_3649)
);

OR2x6_ASAP7_75t_SL g3650 ( 
.A(n_3555),
.B(n_88),
.Y(n_3650)
);

HAxp5_ASAP7_75t_L g3651 ( 
.A(n_3569),
.B(n_89),
.CON(n_3651),
.SN(n_3651)
);

INVx4_ASAP7_75t_L g3652 ( 
.A(n_3444),
.Y(n_3652)
);

BUFx6f_ASAP7_75t_L g3653 ( 
.A(n_3533),
.Y(n_3653)
);

BUFx3_ASAP7_75t_L g3654 ( 
.A(n_3525),
.Y(n_3654)
);

OAI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3545),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_3655)
);

INVxp67_ASAP7_75t_SL g3656 ( 
.A(n_3448),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3440),
.Y(n_3657)
);

INVx4_ASAP7_75t_L g3658 ( 
.A(n_3425),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3517),
.A2(n_622),
.B(n_621),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_3507),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_3579),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_3425),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3475),
.B(n_91),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3583),
.Y(n_3664)
);

AND2x4_ASAP7_75t_L g3665 ( 
.A(n_3489),
.B(n_693),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3478),
.B(n_3510),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3517),
.A2(n_625),
.B(n_624),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_3496),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3504),
.A2(n_627),
.B(n_626),
.Y(n_3669)
);

AND2x4_ASAP7_75t_L g3670 ( 
.A(n_3511),
.B(n_628),
.Y(n_3670)
);

INVx1_ASAP7_75t_SL g3671 ( 
.A(n_3454),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3442),
.B(n_92),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3581),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3482),
.Y(n_3674)
);

INVx2_ASAP7_75t_SL g3675 ( 
.A(n_3497),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3482),
.Y(n_3676)
);

INVxp67_ASAP7_75t_L g3677 ( 
.A(n_3421),
.Y(n_3677)
);

BUFx6f_ASAP7_75t_L g3678 ( 
.A(n_3425),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3591),
.B(n_3429),
.Y(n_3679)
);

INVx2_ASAP7_75t_SL g3680 ( 
.A(n_3535),
.Y(n_3680)
);

INVx1_ASAP7_75t_SL g3681 ( 
.A(n_3405),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3504),
.A2(n_632),
.B(n_631),
.Y(n_3682)
);

AO22x1_ASAP7_75t_L g3683 ( 
.A1(n_3495),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_3494),
.A2(n_97),
.B1(n_93),
.B2(n_96),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3592),
.B(n_633),
.Y(n_3685)
);

BUFx6f_ASAP7_75t_L g3686 ( 
.A(n_3438),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3560),
.B(n_97),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3483),
.Y(n_3688)
);

BUFx3_ASAP7_75t_L g3689 ( 
.A(n_3467),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3538),
.B(n_98),
.Y(n_3690)
);

INVx2_ASAP7_75t_SL g3691 ( 
.A(n_3535),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3446),
.Y(n_3692)
);

O2A1O1Ixp33_ASAP7_75t_L g3693 ( 
.A1(n_3506),
.A2(n_3604),
.B(n_3595),
.C(n_3557),
.Y(n_3693)
);

INVx4_ASAP7_75t_L g3694 ( 
.A(n_3444),
.Y(n_3694)
);

OR2x6_ASAP7_75t_SL g3695 ( 
.A(n_3574),
.B(n_98),
.Y(n_3695)
);

O2A1O1Ixp33_ASAP7_75t_L g3696 ( 
.A1(n_3585),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_3696)
);

NAND3xp33_ASAP7_75t_SL g3697 ( 
.A(n_3502),
.B(n_99),
.C(n_100),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3542),
.B(n_101),
.Y(n_3698)
);

OAI22xp5_ASAP7_75t_L g3699 ( 
.A1(n_3508),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3483),
.Y(n_3700)
);

BUFx6f_ASAP7_75t_L g3701 ( 
.A(n_3438),
.Y(n_3701)
);

AOI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3606),
.A2(n_637),
.B(n_636),
.Y(n_3702)
);

AND2x6_ASAP7_75t_L g3703 ( 
.A(n_3599),
.B(n_638),
.Y(n_3703)
);

INVx3_ASAP7_75t_L g3704 ( 
.A(n_3438),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3452),
.Y(n_3705)
);

BUFx6f_ASAP7_75t_L g3706 ( 
.A(n_3439),
.Y(n_3706)
);

OR2x6_ASAP7_75t_L g3707 ( 
.A(n_3492),
.B(n_640),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3529),
.B(n_102),
.Y(n_3708)
);

BUFx6f_ASAP7_75t_L g3709 ( 
.A(n_3439),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3531),
.B(n_103),
.Y(n_3710)
);

BUFx2_ASAP7_75t_L g3711 ( 
.A(n_3453),
.Y(n_3711)
);

BUFx12f_ASAP7_75t_L g3712 ( 
.A(n_3488),
.Y(n_3712)
);

BUFx2_ASAP7_75t_L g3713 ( 
.A(n_3404),
.Y(n_3713)
);

OAI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3589),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3547),
.B(n_105),
.Y(n_3715)
);

INVx4_ASAP7_75t_L g3716 ( 
.A(n_3439),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3459),
.Y(n_3717)
);

AOI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3599),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3550),
.B(n_107),
.Y(n_3719)
);

A2O1A1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3443),
.A2(n_3450),
.B(n_3586),
.C(n_3501),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3474),
.Y(n_3721)
);

NAND2xp33_ASAP7_75t_L g3722 ( 
.A(n_3477),
.B(n_108),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_3485),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3414),
.B(n_3530),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3491),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3553),
.B(n_110),
.Y(n_3726)
);

AOI21x1_ASAP7_75t_SL g3727 ( 
.A1(n_3584),
.A2(n_111),
.B(n_112),
.Y(n_3727)
);

A2O1A1Ixp33_ASAP7_75t_L g3728 ( 
.A1(n_3501),
.A2(n_114),
.B(n_111),
.C(n_113),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3568),
.Y(n_3729)
);

CKINVDCx14_ASAP7_75t_R g3730 ( 
.A(n_3407),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3513),
.B(n_113),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3568),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3485),
.Y(n_3733)
);

A2O1A1Ixp33_ASAP7_75t_SL g3734 ( 
.A1(n_3577),
.A2(n_118),
.B(n_114),
.C(n_115),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3408),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3548),
.Y(n_3736)
);

CKINVDCx16_ASAP7_75t_R g3737 ( 
.A(n_3400),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3520),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3573),
.Y(n_3739)
);

INVx5_ASAP7_75t_L g3740 ( 
.A(n_3492),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3556),
.B(n_119),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3409),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3399),
.B(n_120),
.Y(n_3743)
);

BUFx2_ASAP7_75t_L g3744 ( 
.A(n_3400),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3588),
.Y(n_3745)
);

INVx1_ASAP7_75t_SL g3746 ( 
.A(n_3558),
.Y(n_3746)
);

INVxp67_ASAP7_75t_SL g3747 ( 
.A(n_3546),
.Y(n_3747)
);

AOI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3473),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_3748)
);

INVx3_ASAP7_75t_L g3749 ( 
.A(n_3485),
.Y(n_3749)
);

INVx2_ASAP7_75t_SL g3750 ( 
.A(n_3559),
.Y(n_3750)
);

O2A1O1Ixp5_ASAP7_75t_L g3751 ( 
.A1(n_3499),
.A2(n_125),
.B(n_122),
.C(n_124),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3565),
.Y(n_3752)
);

AOI22xp33_ASAP7_75t_L g3753 ( 
.A1(n_3537),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3532),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3424),
.B(n_128),
.Y(n_3755)
);

BUFx3_ASAP7_75t_L g3756 ( 
.A(n_3578),
.Y(n_3756)
);

AOI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_3597),
.A2(n_643),
.B(n_642),
.Y(n_3757)
);

AOI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_3549),
.A2(n_648),
.B(n_647),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3580),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3582),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3605),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3455),
.B(n_129),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_SL g3763 ( 
.A(n_3523),
.B(n_649),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3418),
.A2(n_132),
.B1(n_129),
.B2(n_131),
.Y(n_3764)
);

O2A1O1Ixp33_ASAP7_75t_L g3765 ( 
.A1(n_3456),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_3765)
);

OR2x2_ASAP7_75t_L g3766 ( 
.A(n_3539),
.B(n_133),
.Y(n_3766)
);

BUFx2_ASAP7_75t_L g3767 ( 
.A(n_3590),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3471),
.B(n_134),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3605),
.Y(n_3769)
);

A2O1A1Ixp33_ASAP7_75t_L g3770 ( 
.A1(n_3514),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3587),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3500),
.Y(n_3772)
);

BUFx6f_ASAP7_75t_L g3773 ( 
.A(n_3410),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3527),
.Y(n_3774)
);

NAND2x1_ASAP7_75t_SL g3775 ( 
.A(n_3563),
.B(n_135),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3576),
.Y(n_3776)
);

BUFx4f_ASAP7_75t_L g3777 ( 
.A(n_3562),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3451),
.B(n_3463),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3476),
.B(n_136),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3503),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_3780)
);

NOR2xp67_ASAP7_75t_L g3781 ( 
.A(n_3509),
.B(n_138),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3598),
.Y(n_3782)
);

AOI21x1_ASAP7_75t_L g3783 ( 
.A1(n_3484),
.A2(n_139),
.B(n_141),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3524),
.B(n_141),
.Y(n_3784)
);

AND2x4_ASAP7_75t_L g3785 ( 
.A(n_3590),
.B(n_692),
.Y(n_3785)
);

AOI22xp33_ASAP7_75t_L g3786 ( 
.A1(n_3437),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_3786)
);

INVx4_ASAP7_75t_L g3787 ( 
.A(n_3444),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3412),
.Y(n_3788)
);

INVx1_ASAP7_75t_SL g3789 ( 
.A(n_3426),
.Y(n_3789)
);

INVx3_ASAP7_75t_L g3790 ( 
.A(n_3412),
.Y(n_3790)
);

AND2x4_ASAP7_75t_L g3791 ( 
.A(n_3431),
.B(n_650),
.Y(n_3791)
);

INVx8_ASAP7_75t_L g3792 ( 
.A(n_3562),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3484),
.Y(n_3793)
);

BUFx2_ASAP7_75t_L g3794 ( 
.A(n_3431),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3486),
.B(n_142),
.Y(n_3795)
);

BUFx3_ASAP7_75t_L g3796 ( 
.A(n_3447),
.Y(n_3796)
);

INVx4_ASAP7_75t_L g3797 ( 
.A(n_3410),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3567),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3447),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3479),
.Y(n_3800)
);

OAI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3544),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3479),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3522),
.Y(n_3803)
);

A2O1A1Ixp33_ASAP7_75t_L g3804 ( 
.A1(n_3601),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_3804)
);

OAI22xp5_ASAP7_75t_SL g3805 ( 
.A1(n_3551),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_3805)
);

BUFx2_ASAP7_75t_L g3806 ( 
.A(n_3522),
.Y(n_3806)
);

INVx4_ASAP7_75t_L g3807 ( 
.A(n_3526),
.Y(n_3807)
);

AOI22xp5_ASAP7_75t_SL g3808 ( 
.A1(n_3426),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3808)
);

OR2x6_ASAP7_75t_L g3809 ( 
.A(n_3420),
.B(n_651),
.Y(n_3809)
);

NOR2xp33_ASAP7_75t_L g3810 ( 
.A(n_3490),
.B(n_149),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3571),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3415),
.B(n_150),
.Y(n_3812)
);

BUFx2_ASAP7_75t_L g3813 ( 
.A(n_3526),
.Y(n_3813)
);

BUFx3_ASAP7_75t_L g3814 ( 
.A(n_3472),
.Y(n_3814)
);

INVx5_ASAP7_75t_L g3815 ( 
.A(n_3493),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3461),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3461),
.Y(n_3817)
);

OR2x2_ASAP7_75t_L g3818 ( 
.A(n_3505),
.B(n_151),
.Y(n_3818)
);

AND2x4_ASAP7_75t_L g3819 ( 
.A(n_3480),
.B(n_691),
.Y(n_3819)
);

OR2x6_ASAP7_75t_L g3820 ( 
.A(n_3493),
.B(n_652),
.Y(n_3820)
);

O2A1O1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3433),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_3821)
);

BUFx6f_ASAP7_75t_L g3822 ( 
.A(n_3480),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3521),
.Y(n_3823)
);

BUFx3_ASAP7_75t_L g3824 ( 
.A(n_3566),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3518),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3602),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3427),
.B(n_152),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3515),
.A2(n_156),
.B1(n_153),
.B2(n_154),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3534),
.A2(n_159),
.B1(n_154),
.B2(n_158),
.Y(n_3829)
);

AND2x4_ASAP7_75t_SL g3830 ( 
.A(n_3536),
.B(n_654),
.Y(n_3830)
);

INVxp67_ASAP7_75t_SL g3831 ( 
.A(n_3571),
.Y(n_3831)
);

HB1xp67_ASAP7_75t_L g3832 ( 
.A(n_3572),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3572),
.Y(n_3833)
);

NAND2x1p5_ASAP7_75t_L g3834 ( 
.A(n_3815),
.B(n_3536),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3644),
.Y(n_3835)
);

BUFx6f_ASAP7_75t_L g3836 ( 
.A(n_3617),
.Y(n_3836)
);

OR2x2_ASAP7_75t_L g3837 ( 
.A(n_3664),
.B(n_3401),
.Y(n_3837)
);

BUFx6f_ASAP7_75t_L g3838 ( 
.A(n_3617),
.Y(n_3838)
);

BUFx6f_ASAP7_75t_L g3839 ( 
.A(n_3617),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3640),
.Y(n_3840)
);

A2O1A1Ixp33_ASAP7_75t_L g3841 ( 
.A1(n_3693),
.A2(n_3541),
.B(n_3468),
.C(n_3564),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3645),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3718),
.A2(n_3465),
.B1(n_3552),
.B2(n_3607),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3648),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3656),
.B(n_3449),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3612),
.Y(n_3846)
);

OAI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3636),
.A2(n_3552),
.B1(n_3561),
.B2(n_3516),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3622),
.Y(n_3848)
);

BUFx6f_ASAP7_75t_L g3849 ( 
.A(n_3632),
.Y(n_3849)
);

CKINVDCx8_ASAP7_75t_R g3850 ( 
.A(n_3641),
.Y(n_3850)
);

BUFx6f_ASAP7_75t_L g3851 ( 
.A(n_3632),
.Y(n_3851)
);

INVx8_ASAP7_75t_L g3852 ( 
.A(n_3820),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3677),
.B(n_3554),
.Y(n_3853)
);

INVx2_ASAP7_75t_SL g3854 ( 
.A(n_3643),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3681),
.B(n_3566),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3623),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3637),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3638),
.Y(n_3858)
);

BUFx3_ASAP7_75t_L g3859 ( 
.A(n_3654),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_3782),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3722),
.A2(n_3466),
.B(n_3428),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3642),
.Y(n_3862)
);

AND2x4_ASAP7_75t_L g3863 ( 
.A(n_3744),
.B(n_655),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3616),
.B(n_160),
.Y(n_3864)
);

BUFx6f_ASAP7_75t_L g3865 ( 
.A(n_3632),
.Y(n_3865)
);

OAI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3655),
.A2(n_3748),
.B1(n_3735),
.B2(n_3720),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3674),
.Y(n_3867)
);

AND2x4_ASAP7_75t_L g3868 ( 
.A(n_3626),
.B(n_656),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3615),
.B(n_160),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_3618),
.B(n_161),
.Y(n_3870)
);

AOI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3703),
.A2(n_3593),
.B1(n_3419),
.B2(n_164),
.Y(n_3871)
);

O2A1O1Ixp33_ASAP7_75t_L g3872 ( 
.A1(n_3821),
.A2(n_164),
.B(n_161),
.C(n_162),
.Y(n_3872)
);

INVx1_ASAP7_75t_SL g3873 ( 
.A(n_3671),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_L g3874 ( 
.A(n_3639),
.B(n_162),
.Y(n_3874)
);

BUFx12f_ASAP7_75t_L g3875 ( 
.A(n_3646),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3613),
.Y(n_3876)
);

OR2x2_ASAP7_75t_L g3877 ( 
.A(n_3729),
.B(n_165),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3676),
.Y(n_3878)
);

INVxp67_ASAP7_75t_L g3879 ( 
.A(n_3711),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3611),
.Y(n_3880)
);

OR2x6_ASAP7_75t_L g3881 ( 
.A(n_3792),
.B(n_657),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_L g3882 ( 
.A1(n_3697),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3619),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3737),
.B(n_167),
.Y(n_3884)
);

BUFx6f_ASAP7_75t_L g3885 ( 
.A(n_3653),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3666),
.B(n_168),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3630),
.Y(n_3887)
);

NAND2xp33_ASAP7_75t_L g3888 ( 
.A(n_3703),
.B(n_168),
.Y(n_3888)
);

INVx2_ASAP7_75t_SL g3889 ( 
.A(n_3610),
.Y(n_3889)
);

INVx5_ASAP7_75t_L g3890 ( 
.A(n_3809),
.Y(n_3890)
);

BUFx3_ASAP7_75t_L g3891 ( 
.A(n_3633),
.Y(n_3891)
);

NAND2x1p5_ASAP7_75t_L g3892 ( 
.A(n_3815),
.B(n_659),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3745),
.B(n_171),
.Y(n_3893)
);

AOI22xp33_ASAP7_75t_L g3894 ( 
.A1(n_3703),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_3894)
);

OAI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3770),
.A2(n_172),
.B(n_174),
.Y(n_3895)
);

AND2x4_ASAP7_75t_L g3896 ( 
.A(n_3689),
.B(n_660),
.Y(n_3896)
);

NAND2x1_ASAP7_75t_L g3897 ( 
.A(n_3732),
.B(n_3652),
.Y(n_3897)
);

NOR2xp33_ASAP7_75t_L g3898 ( 
.A(n_3695),
.B(n_174),
.Y(n_3898)
);

INVx5_ASAP7_75t_L g3899 ( 
.A(n_3809),
.Y(n_3899)
);

INVx3_ASAP7_75t_L g3900 ( 
.A(n_3796),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_SL g3901 ( 
.A(n_3635),
.Y(n_3901)
);

BUFx6f_ASAP7_75t_L g3902 ( 
.A(n_3653),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3631),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3798),
.B(n_175),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3679),
.B(n_177),
.Y(n_3905)
);

NAND2x1p5_ASAP7_75t_L g3906 ( 
.A(n_3815),
.B(n_662),
.Y(n_3906)
);

INVx5_ASAP7_75t_L g3907 ( 
.A(n_3707),
.Y(n_3907)
);

NOR2xp67_ASAP7_75t_L g3908 ( 
.A(n_3673),
.B(n_178),
.Y(n_3908)
);

BUFx12f_ASAP7_75t_L g3909 ( 
.A(n_3668),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3688),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3700),
.Y(n_3911)
);

BUFx2_ASAP7_75t_L g3912 ( 
.A(n_3832),
.Y(n_3912)
);

BUFx12f_ASAP7_75t_L g3913 ( 
.A(n_3660),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3679),
.B(n_179),
.Y(n_3914)
);

INVx5_ASAP7_75t_L g3915 ( 
.A(n_3707),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3793),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3625),
.Y(n_3917)
);

INVx2_ASAP7_75t_SL g3918 ( 
.A(n_3634),
.Y(n_3918)
);

BUFx12f_ASAP7_75t_L g3919 ( 
.A(n_3731),
.Y(n_3919)
);

AOI22xp33_ASAP7_75t_L g3920 ( 
.A1(n_3805),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3920)
);

OAI21xp33_ASAP7_75t_SL g3921 ( 
.A1(n_3775),
.A2(n_180),
.B(n_181),
.Y(n_3921)
);

BUFx3_ASAP7_75t_L g3922 ( 
.A(n_3634),
.Y(n_3922)
);

BUFx2_ASAP7_75t_L g3923 ( 
.A(n_3833),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3811),
.Y(n_3924)
);

INVx5_ASAP7_75t_L g3925 ( 
.A(n_3820),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3747),
.B(n_3742),
.Y(n_3926)
);

INVx1_ASAP7_75t_SL g3927 ( 
.A(n_3713),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3739),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3825),
.B(n_3823),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3771),
.B(n_182),
.Y(n_3930)
);

INVx3_ASAP7_75t_L g3931 ( 
.A(n_3756),
.Y(n_3931)
);

BUFx2_ASAP7_75t_L g3932 ( 
.A(n_3831),
.Y(n_3932)
);

INVx6_ASAP7_75t_L g3933 ( 
.A(n_3773),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3738),
.B(n_183),
.Y(n_3934)
);

INVx2_ASAP7_75t_SL g3935 ( 
.A(n_3675),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3827),
.B(n_185),
.Y(n_3936)
);

INVx2_ASAP7_75t_SL g3937 ( 
.A(n_3792),
.Y(n_3937)
);

AOI222xp33_ASAP7_75t_L g3938 ( 
.A1(n_3684),
.A2(n_189),
.B1(n_191),
.B2(n_186),
.C1(n_187),
.C2(n_190),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3761),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3794),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3627),
.Y(n_3941)
);

OAI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_3754),
.A2(n_192),
.B1(n_189),
.B2(n_190),
.Y(n_3942)
);

AO21x2_ASAP7_75t_L g3943 ( 
.A1(n_3629),
.A2(n_192),
.B(n_193),
.Y(n_3943)
);

INVxp67_ASAP7_75t_L g3944 ( 
.A(n_3803),
.Y(n_3944)
);

OR2x6_ASAP7_75t_L g3945 ( 
.A(n_3817),
.B(n_3652),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3806),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3724),
.B(n_193),
.Y(n_3947)
);

INVx3_ASAP7_75t_L g3948 ( 
.A(n_3653),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3769),
.B(n_194),
.Y(n_3949)
);

BUFx6f_ASAP7_75t_L g3950 ( 
.A(n_3662),
.Y(n_3950)
);

BUFx2_ASAP7_75t_L g3951 ( 
.A(n_3813),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3752),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_L g3953 ( 
.A(n_3762),
.B(n_195),
.Y(n_3953)
);

OR2x2_ASAP7_75t_L g3954 ( 
.A(n_3789),
.B(n_195),
.Y(n_3954)
);

INVx4_ASAP7_75t_L g3955 ( 
.A(n_3662),
.Y(n_3955)
);

INVx1_ASAP7_75t_SL g3956 ( 
.A(n_3661),
.Y(n_3956)
);

INVx3_ASAP7_75t_L g3957 ( 
.A(n_3662),
.Y(n_3957)
);

BUFx6f_ASAP7_75t_L g3958 ( 
.A(n_3678),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3759),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3657),
.Y(n_3960)
);

AOI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_3740),
.A2(n_197),
.B(n_198),
.Y(n_3961)
);

OAI22xp5_ASAP7_75t_SL g3962 ( 
.A1(n_3730),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_L g3963 ( 
.A1(n_3764),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3760),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3692),
.B(n_200),
.Y(n_3965)
);

NOR2xp67_ASAP7_75t_L g3966 ( 
.A(n_3740),
.B(n_3708),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3705),
.Y(n_3967)
);

OR2x2_ASAP7_75t_L g3968 ( 
.A(n_3826),
.B(n_201),
.Y(n_3968)
);

INVx1_ASAP7_75t_SL g3969 ( 
.A(n_3746),
.Y(n_3969)
);

AND2x4_ASAP7_75t_L g3970 ( 
.A(n_3767),
.B(n_664),
.Y(n_3970)
);

OR2x6_ASAP7_75t_L g3971 ( 
.A(n_3694),
.B(n_667),
.Y(n_3971)
);

OAI22xp5_ASAP7_75t_L g3972 ( 
.A1(n_3753),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3717),
.Y(n_3973)
);

BUFx6f_ASAP7_75t_L g3974 ( 
.A(n_3678),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3721),
.Y(n_3975)
);

A2O1A1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3696),
.A2(n_205),
.B(n_202),
.C(n_203),
.Y(n_3976)
);

BUFx10_ASAP7_75t_L g3977 ( 
.A(n_3773),
.Y(n_3977)
);

AND2x4_ASAP7_75t_L g3978 ( 
.A(n_3788),
.B(n_678),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_3712),
.Y(n_3979)
);

INVx3_ASAP7_75t_L g3980 ( 
.A(n_3678),
.Y(n_3980)
);

BUFx2_ASAP7_75t_L g3981 ( 
.A(n_3807),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3725),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3799),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3736),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3750),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3802),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3755),
.B(n_205),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3772),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3814),
.B(n_206),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3699),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_3686),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3783),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3783),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3743),
.B(n_210),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3768),
.B(n_211),
.Y(n_3995)
);

INVx4_ASAP7_75t_L g3996 ( 
.A(n_3686),
.Y(n_3996)
);

INVxp67_ASAP7_75t_L g3997 ( 
.A(n_3774),
.Y(n_3997)
);

AND2x4_ASAP7_75t_L g3998 ( 
.A(n_3824),
.B(n_680),
.Y(n_3998)
);

CKINVDCx5p33_ASAP7_75t_R g3999 ( 
.A(n_3686),
.Y(n_3999)
);

OAI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3829),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3714),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_4001)
);

INVx5_ASAP7_75t_L g4002 ( 
.A(n_3694),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3776),
.Y(n_4003)
);

AND2x4_ASAP7_75t_L g4004 ( 
.A(n_3790),
.B(n_684),
.Y(n_4004)
);

CKINVDCx20_ASAP7_75t_R g4005 ( 
.A(n_3777),
.Y(n_4005)
);

BUFx2_ASAP7_75t_L g4006 ( 
.A(n_3807),
.Y(n_4006)
);

AO22x1_ASAP7_75t_L g4007 ( 
.A1(n_3740),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3690),
.Y(n_4008)
);

INVx2_ASAP7_75t_SL g4009 ( 
.A(n_3701),
.Y(n_4009)
);

NOR2x1_ASAP7_75t_SL g4010 ( 
.A(n_3787),
.B(n_216),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3779),
.B(n_217),
.Y(n_4011)
);

NAND2xp33_ASAP7_75t_L g4012 ( 
.A(n_3804),
.B(n_217),
.Y(n_4012)
);

BUFx4_ASAP7_75t_SL g4013 ( 
.A(n_3784),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3628),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3880),
.B(n_3687),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3940),
.B(n_3778),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3888),
.A2(n_3624),
.B(n_3614),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3940),
.B(n_3672),
.Y(n_4018)
);

BUFx2_ASAP7_75t_L g4019 ( 
.A(n_3945),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3945),
.B(n_3680),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3924),
.Y(n_4021)
);

O2A1O1Ixp33_ASAP7_75t_SL g4022 ( 
.A1(n_3898),
.A2(n_3728),
.B(n_3734),
.C(n_3812),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3946),
.Y(n_4023)
);

OAI21x1_ASAP7_75t_L g4024 ( 
.A1(n_3897),
.A2(n_3609),
.B(n_3629),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3867),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3897),
.A2(n_3993),
.B(n_3992),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3866),
.A2(n_3810),
.B1(n_3795),
.B2(n_3621),
.Y(n_4027)
);

INVxp67_ASAP7_75t_L g4028 ( 
.A(n_3988),
.Y(n_4028)
);

OAI21x1_ASAP7_75t_L g4029 ( 
.A1(n_3861),
.A2(n_3727),
.B(n_3620),
.Y(n_4029)
);

AND2x4_ASAP7_75t_L g4030 ( 
.A(n_3946),
.B(n_3691),
.Y(n_4030)
);

NAND2x1_ASAP7_75t_L g4031 ( 
.A(n_3932),
.B(n_3787),
.Y(n_4031)
);

O2A1O1Ixp33_ASAP7_75t_L g4032 ( 
.A1(n_3976),
.A2(n_3801),
.B(n_3828),
.C(n_3651),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3860),
.B(n_3818),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3951),
.B(n_3800),
.Y(n_4034)
);

OAI21x1_ASAP7_75t_L g4035 ( 
.A1(n_3834),
.A2(n_3837),
.B(n_3878),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3937),
.B(n_3650),
.Y(n_4036)
);

CKINVDCx6p67_ASAP7_75t_R g4037 ( 
.A(n_3922),
.Y(n_4037)
);

HB1xp67_ASAP7_75t_L g4038 ( 
.A(n_3912),
.Y(n_4038)
);

HB1xp67_ASAP7_75t_L g4039 ( 
.A(n_3912),
.Y(n_4039)
);

AND2x6_ASAP7_75t_L g4040 ( 
.A(n_3871),
.B(n_3816),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3951),
.Y(n_4041)
);

NAND2x1p5_ASAP7_75t_L g4042 ( 
.A(n_3907),
.B(n_3816),
.Y(n_4042)
);

HB1xp67_ASAP7_75t_L g4043 ( 
.A(n_3932),
.Y(n_4043)
);

OA21x2_ASAP7_75t_L g4044 ( 
.A1(n_3910),
.A2(n_3663),
.B(n_3775),
.Y(n_4044)
);

BUFx3_ASAP7_75t_L g4045 ( 
.A(n_3875),
.Y(n_4045)
);

OAI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3841),
.A2(n_3758),
.B(n_3757),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_SL g4047 ( 
.A1(n_3918),
.A2(n_4005),
.B(n_4011),
.C(n_3995),
.Y(n_4047)
);

BUFx10_ASAP7_75t_L g4048 ( 
.A(n_3870),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_SL g4049 ( 
.A1(n_3907),
.A2(n_3808),
.B1(n_3822),
.B2(n_3816),
.Y(n_4049)
);

OAI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_3907),
.A2(n_3786),
.B1(n_3780),
.B2(n_3608),
.Y(n_4050)
);

OAI21x1_ASAP7_75t_L g4051 ( 
.A1(n_3911),
.A2(n_3667),
.B(n_3659),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3923),
.Y(n_4052)
);

O2A1O1Ixp33_ASAP7_75t_SL g4053 ( 
.A1(n_3895),
.A2(n_3766),
.B(n_3710),
.C(n_3719),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3944),
.B(n_3658),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3926),
.B(n_3781),
.Y(n_4055)
);

AO31x2_ASAP7_75t_L g4056 ( 
.A1(n_3981),
.A2(n_3716),
.A3(n_3797),
.B(n_3682),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3916),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3927),
.B(n_3704),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3969),
.B(n_3715),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3923),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3961),
.A2(n_3669),
.B(n_3765),
.Y(n_4061)
);

BUFx2_ASAP7_75t_L g4062 ( 
.A(n_3981),
.Y(n_4062)
);

AO31x2_ASAP7_75t_L g4063 ( 
.A1(n_4006),
.A2(n_3797),
.A3(n_3698),
.B(n_3741),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3846),
.Y(n_4064)
);

AO21x1_ASAP7_75t_L g4065 ( 
.A1(n_3929),
.A2(n_3726),
.B(n_3670),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_4012),
.A2(n_3685),
.B1(n_3647),
.B2(n_3665),
.Y(n_4066)
);

A2O1A1Ixp33_ASAP7_75t_L g4067 ( 
.A1(n_3872),
.A2(n_3751),
.B(n_3830),
.C(n_3702),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3835),
.Y(n_4068)
);

OAI21x1_ASAP7_75t_L g4069 ( 
.A1(n_3930),
.A2(n_3763),
.B(n_3749),
.Y(n_4069)
);

OAI22xp5_ASAP7_75t_L g4070 ( 
.A1(n_3915),
.A2(n_3822),
.B1(n_3665),
.B2(n_3649),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3844),
.Y(n_4071)
);

AOI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_3890),
.A2(n_3683),
.B(n_3670),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_SL g4073 ( 
.A1(n_4010),
.A2(n_3822),
.B(n_3706),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3962),
.A2(n_3649),
.B1(n_3819),
.B2(n_3785),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3879),
.B(n_4008),
.Y(n_4075)
);

INVx3_ASAP7_75t_L g4076 ( 
.A(n_4006),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3845),
.A2(n_3706),
.B(n_3701),
.Y(n_4077)
);

OAI21x1_ASAP7_75t_L g4078 ( 
.A1(n_3949),
.A2(n_3706),
.B(n_3701),
.Y(n_4078)
);

AND2x4_ASAP7_75t_L g4079 ( 
.A(n_3984),
.B(n_3709),
.Y(n_4079)
);

OAI21x1_ASAP7_75t_L g4080 ( 
.A1(n_3939),
.A2(n_3723),
.B(n_3709),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_3953),
.A2(n_3819),
.B1(n_3785),
.B2(n_3791),
.Y(n_4081)
);

OA21x2_ASAP7_75t_L g4082 ( 
.A1(n_3928),
.A2(n_3791),
.B(n_3723),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3848),
.Y(n_4083)
);

OAI21x1_ASAP7_75t_L g4084 ( 
.A1(n_3877),
.A2(n_3723),
.B(n_3709),
.Y(n_4084)
);

OAI21x1_ASAP7_75t_L g4085 ( 
.A1(n_3892),
.A2(n_3733),
.B(n_3773),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3856),
.Y(n_4086)
);

OAI21x1_ASAP7_75t_L g4087 ( 
.A1(n_3906),
.A2(n_3733),
.B(n_220),
.Y(n_4087)
);

OA21x2_ASAP7_75t_L g4088 ( 
.A1(n_3857),
.A2(n_3733),
.B(n_221),
.Y(n_4088)
);

BUFx2_ASAP7_75t_L g4089 ( 
.A(n_3931),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3858),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3840),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3862),
.Y(n_4092)
);

NOR2xp33_ASAP7_75t_L g4093 ( 
.A(n_3873),
.B(n_221),
.Y(n_4093)
);

NAND3xp33_ASAP7_75t_L g4094 ( 
.A(n_3938),
.B(n_222),
.C(n_223),
.Y(n_4094)
);

AOI22xp33_ASAP7_75t_SL g4095 ( 
.A1(n_3915),
.A2(n_225),
.B1(n_222),
.B2(n_224),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_3850),
.B(n_225),
.Y(n_4096)
);

OAI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_3921),
.A2(n_226),
.B(n_227),
.Y(n_4097)
);

AOI22xp33_ASAP7_75t_SL g4098 ( 
.A1(n_3915),
.A2(n_230),
.B1(n_226),
.B2(n_229),
.Y(n_4098)
);

HB1xp67_ASAP7_75t_L g4099 ( 
.A(n_4003),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3960),
.B(n_230),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3975),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3952),
.Y(n_4102)
);

OAI21x1_ASAP7_75t_L g4103 ( 
.A1(n_3966),
.A2(n_231),
.B(n_232),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3982),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3900),
.A2(n_233),
.B(n_234),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3959),
.Y(n_4106)
);

CKINVDCx5p33_ASAP7_75t_R g4107 ( 
.A(n_3901),
.Y(n_4107)
);

OA21x2_ASAP7_75t_L g4108 ( 
.A1(n_3869),
.A2(n_233),
.B(n_234),
.Y(n_4108)
);

OR2x6_ASAP7_75t_L g4109 ( 
.A(n_3852),
.B(n_235),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3842),
.Y(n_4110)
);

OAI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3936),
.A2(n_235),
.B(n_236),
.Y(n_4111)
);

AND2x4_ASAP7_75t_L g4112 ( 
.A(n_3985),
.B(n_236),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3876),
.Y(n_4113)
);

OAI21x1_ASAP7_75t_L g4114 ( 
.A1(n_3934),
.A2(n_237),
.B(n_238),
.Y(n_4114)
);

INVx1_ASAP7_75t_SL g4115 ( 
.A(n_3956),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3964),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3983),
.Y(n_4117)
);

OAI21x1_ASAP7_75t_L g4118 ( 
.A1(n_3965),
.A2(n_237),
.B(n_238),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3986),
.Y(n_4119)
);

OA21x2_ASAP7_75t_L g4120 ( 
.A1(n_3904),
.A2(n_239),
.B(n_240),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_3997),
.B(n_240),
.Y(n_4121)
);

OAI221xp5_ASAP7_75t_SL g4122 ( 
.A1(n_3920),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.C(n_244),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3883),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3917),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_3968),
.A2(n_241),
.B(n_242),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3941),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3887),
.B(n_244),
.Y(n_4127)
);

BUFx2_ASAP7_75t_L g4128 ( 
.A(n_3955),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3967),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_3886),
.B(n_3913),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3973),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3854),
.B(n_246),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3893),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3855),
.B(n_529),
.Y(n_4134)
);

AOI22xp33_ASAP7_75t_L g4135 ( 
.A1(n_3890),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_4135)
);

AOI222xp33_ASAP7_75t_L g4136 ( 
.A1(n_3942),
.A2(n_4000),
.B1(n_3882),
.B2(n_3972),
.C1(n_4014),
.C2(n_4001),
.Y(n_4136)
);

AO21x2_ASAP7_75t_L g4137 ( 
.A1(n_3943),
.A2(n_247),
.B(n_249),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3890),
.A2(n_250),
.B(n_251),
.Y(n_4138)
);

AOI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_3899),
.A2(n_254),
.B1(n_251),
.B2(n_253),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4002),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3864),
.B(n_528),
.Y(n_4141)
);

OAI21x1_ASAP7_75t_L g4142 ( 
.A1(n_3948),
.A2(n_253),
.B(n_256),
.Y(n_4142)
);

NAND2x1p5_ASAP7_75t_L g4143 ( 
.A(n_3925),
.B(n_256),
.Y(n_4143)
);

AND2x4_ASAP7_75t_L g4144 ( 
.A(n_4002),
.B(n_258),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3947),
.B(n_528),
.Y(n_4145)
);

AOI22xp33_ASAP7_75t_L g4146 ( 
.A1(n_3899),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4146)
);

OAI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3847),
.A2(n_259),
.B(n_260),
.Y(n_4147)
);

AOI22xp5_ASAP7_75t_L g4148 ( 
.A1(n_3899),
.A2(n_3925),
.B1(n_3843),
.B2(n_3894),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4002),
.Y(n_4149)
);

AOI21x1_ASAP7_75t_L g4150 ( 
.A1(n_4007),
.A2(n_261),
.B(n_262),
.Y(n_4150)
);

AND2x4_ASAP7_75t_L g4151 ( 
.A(n_4009),
.B(n_261),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3935),
.B(n_262),
.Y(n_4152)
);

O2A1O1Ixp33_ASAP7_75t_L g4153 ( 
.A1(n_3987),
.A2(n_3994),
.B(n_3903),
.C(n_3990),
.Y(n_4153)
);

OR2x2_ASAP7_75t_L g4154 ( 
.A(n_3954),
.B(n_527),
.Y(n_4154)
);

A2O1A1Ixp33_ASAP7_75t_L g4155 ( 
.A1(n_3925),
.A2(n_527),
.B(n_265),
.C(n_263),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_3957),
.Y(n_4156)
);

CKINVDCx16_ASAP7_75t_R g4157 ( 
.A(n_3909),
.Y(n_4157)
);

BUFx2_ASAP7_75t_L g4158 ( 
.A(n_3996),
.Y(n_4158)
);

INVx1_ASAP7_75t_SL g4159 ( 
.A(n_3859),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3980),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3908),
.Y(n_4161)
);

OAI21x1_ASAP7_75t_L g4162 ( 
.A1(n_3884),
.A2(n_264),
.B(n_265),
.Y(n_4162)
);

AND2x4_ASAP7_75t_L g4163 ( 
.A(n_3889),
.B(n_266),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3853),
.B(n_526),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3836),
.Y(n_4165)
);

BUFx4f_ASAP7_75t_SL g4166 ( 
.A(n_3891),
.Y(n_4166)
);

OA21x2_ASAP7_75t_L g4167 ( 
.A1(n_4026),
.A2(n_3999),
.B(n_3874),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_4076),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_4107),
.B(n_3979),
.Y(n_4169)
);

INVx5_ASAP7_75t_L g4170 ( 
.A(n_4109),
.Y(n_4170)
);

OAI21x1_ASAP7_75t_L g4171 ( 
.A1(n_4035),
.A2(n_3914),
.B(n_3905),
.Y(n_4171)
);

OR2x2_ASAP7_75t_L g4172 ( 
.A(n_4033),
.B(n_3989),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_4076),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_4040),
.A2(n_4046),
.B1(n_4094),
.B2(n_4017),
.Y(n_4174)
);

NAND2x1p5_ASAP7_75t_L g4175 ( 
.A(n_4082),
.B(n_3863),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4021),
.Y(n_4176)
);

OR2x6_ASAP7_75t_L g4177 ( 
.A(n_4072),
.B(n_3852),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_SL g4178 ( 
.A1(n_4040),
.A2(n_3919),
.B1(n_3971),
.B2(n_3868),
.Y(n_4178)
);

BUFx2_ASAP7_75t_R g4179 ( 
.A(n_4045),
.Y(n_4179)
);

OAI21x1_ASAP7_75t_L g4180 ( 
.A1(n_4024),
.A2(n_3963),
.B(n_4013),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4021),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_4077),
.Y(n_4182)
);

BUFx2_ASAP7_75t_SL g4183 ( 
.A(n_4163),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4133),
.B(n_3836),
.Y(n_4184)
);

BUFx6f_ASAP7_75t_L g4185 ( 
.A(n_4037),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4025),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4025),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_4019),
.B(n_3838),
.Y(n_4188)
);

INVxp67_ASAP7_75t_SL g4189 ( 
.A(n_4065),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4057),
.Y(n_4190)
);

NAND2x1p5_ASAP7_75t_L g4191 ( 
.A(n_4082),
.B(n_3896),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_4038),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4063),
.B(n_3838),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_4063),
.B(n_3839),
.Y(n_4194)
);

AOI21x1_ASAP7_75t_L g4195 ( 
.A1(n_4140),
.A2(n_4149),
.B(n_4031),
.Y(n_4195)
);

AOI21x1_ASAP7_75t_L g4196 ( 
.A1(n_4140),
.A2(n_3971),
.B(n_3970),
.Y(n_4196)
);

OAI21x1_ASAP7_75t_L g4197 ( 
.A1(n_4080),
.A2(n_3977),
.B(n_3933),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4057),
.Y(n_4198)
);

INVx3_ASAP7_75t_L g4199 ( 
.A(n_4030),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4090),
.Y(n_4200)
);

BUFx12f_ASAP7_75t_L g4201 ( 
.A(n_4109),
.Y(n_4201)
);

BUFx2_ASAP7_75t_L g4202 ( 
.A(n_4062),
.Y(n_4202)
);

AND2x4_ASAP7_75t_L g4203 ( 
.A(n_4149),
.B(n_3839),
.Y(n_4203)
);

AOI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_4040),
.A2(n_3881),
.B1(n_3998),
.B2(n_3933),
.Y(n_4204)
);

INVx5_ASAP7_75t_L g4205 ( 
.A(n_4144),
.Y(n_4205)
);

CKINVDCx20_ASAP7_75t_R g4206 ( 
.A(n_4166),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4090),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4068),
.Y(n_4208)
);

OAI22xp5_ASAP7_75t_L g4209 ( 
.A1(n_4049),
.A2(n_3881),
.B1(n_3851),
.B2(n_3865),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4148),
.A2(n_3851),
.B1(n_3865),
.B2(n_3849),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4071),
.Y(n_4211)
);

OA21x2_ASAP7_75t_L g4212 ( 
.A1(n_4060),
.A2(n_3978),
.B(n_4004),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_4084),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_SL g4214 ( 
.A1(n_4040),
.A2(n_3885),
.B1(n_3902),
.B2(n_3849),
.Y(n_4214)
);

OAI21x1_ASAP7_75t_L g4215 ( 
.A1(n_4042),
.A2(n_3991),
.B(n_3902),
.Y(n_4215)
);

CKINVDCx11_ASAP7_75t_R g4216 ( 
.A(n_4048),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4083),
.Y(n_4217)
);

OAI21x1_ASAP7_75t_L g4218 ( 
.A1(n_4078),
.A2(n_3950),
.B(n_3885),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4099),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4064),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4086),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4016),
.B(n_3950),
.Y(n_4222)
);

BUFx6f_ASAP7_75t_L g4223 ( 
.A(n_4163),
.Y(n_4223)
);

INVx4_ASAP7_75t_L g4224 ( 
.A(n_4157),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4101),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4104),
.Y(n_4226)
);

CKINVDCx20_ASAP7_75t_R g4227 ( 
.A(n_4159),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4091),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4052),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4063),
.B(n_3958),
.Y(n_4230)
);

CKINVDCx5p33_ASAP7_75t_R g4231 ( 
.A(n_4115),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4091),
.Y(n_4232)
);

AOI22xp5_ASAP7_75t_L g4233 ( 
.A1(n_4050),
.A2(n_3974),
.B1(n_3991),
.B2(n_3958),
.Y(n_4233)
);

BUFx6f_ASAP7_75t_L g4234 ( 
.A(n_4151),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4018),
.B(n_3974),
.Y(n_4235)
);

OAI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_4147),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_4028),
.B(n_267),
.Y(n_4237)
);

AND2x4_ASAP7_75t_L g4238 ( 
.A(n_4020),
.B(n_269),
.Y(n_4238)
);

INVx4_ASAP7_75t_L g4239 ( 
.A(n_4151),
.Y(n_4239)
);

OAI22xp33_ASAP7_75t_L g4240 ( 
.A1(n_4070),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_4240)
);

AOI22xp33_ASAP7_75t_L g4241 ( 
.A1(n_4027),
.A2(n_526),
.B1(n_272),
.B2(n_270),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_4023),
.Y(n_4242)
);

OAI22xp33_ASAP7_75t_L g4243 ( 
.A1(n_4143),
.A2(n_4161),
.B1(n_4097),
.B2(n_4088),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_SL g4244 ( 
.A1(n_4111),
.A2(n_274),
.B1(n_271),
.B2(n_272),
.Y(n_4244)
);

AOI22xp33_ASAP7_75t_SL g4245 ( 
.A1(n_4029),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_4245)
);

BUFx12f_ASAP7_75t_L g4246 ( 
.A(n_4048),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4092),
.Y(n_4247)
);

OAI21x1_ASAP7_75t_L g4248 ( 
.A1(n_4051),
.A2(n_278),
.B(n_279),
.Y(n_4248)
);

OAI21xp5_ASAP7_75t_SL g4249 ( 
.A1(n_4032),
.A2(n_280),
.B(n_281),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4092),
.Y(n_4250)
);

BUFx2_ASAP7_75t_L g4251 ( 
.A(n_4039),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4060),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4110),
.Y(n_4253)
);

INVx2_ASAP7_75t_SL g4254 ( 
.A(n_4034),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4041),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4117),
.Y(n_4256)
);

NOR2xp33_ASAP7_75t_L g4257 ( 
.A(n_4055),
.B(n_280),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4119),
.Y(n_4258)
);

BUFx6f_ASAP7_75t_L g4259 ( 
.A(n_4112),
.Y(n_4259)
);

INVx2_ASAP7_75t_SL g4260 ( 
.A(n_4089),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4113),
.Y(n_4261)
);

OAI22xp33_ASAP7_75t_L g4262 ( 
.A1(n_4161),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4123),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4124),
.Y(n_4264)
);

OAI22xp33_ASAP7_75t_L g4265 ( 
.A1(n_4088),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4131),
.Y(n_4266)
);

CKINVDCx20_ASAP7_75t_R g4267 ( 
.A(n_4058),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4043),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4102),
.Y(n_4269)
);

OAI22xp33_ASAP7_75t_L g4270 ( 
.A1(n_4108),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4106),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_4066),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_4272)
);

AOI21x1_ASAP7_75t_L g4273 ( 
.A1(n_4128),
.A2(n_288),
.B(n_289),
.Y(n_4273)
);

AOI22xp33_ASAP7_75t_L g4274 ( 
.A1(n_4136),
.A2(n_525),
.B1(n_292),
.B2(n_290),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4116),
.Y(n_4275)
);

AOI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4137),
.A2(n_295),
.B1(n_291),
.B2(n_293),
.Y(n_4276)
);

INVx2_ASAP7_75t_SL g4277 ( 
.A(n_4030),
.Y(n_4277)
);

INVx5_ASAP7_75t_L g4278 ( 
.A(n_4144),
.Y(n_4278)
);

AND2x4_ASAP7_75t_L g4279 ( 
.A(n_4020),
.B(n_291),
.Y(n_4279)
);

HB1xp67_ASAP7_75t_L g4280 ( 
.A(n_4044),
.Y(n_4280)
);

AOI22xp33_ASAP7_75t_SL g4281 ( 
.A1(n_4061),
.A2(n_297),
.B1(n_293),
.B2(n_296),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4126),
.Y(n_4282)
);

BUFx12f_ASAP7_75t_L g4283 ( 
.A(n_4154),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4158),
.B(n_296),
.Y(n_4284)
);

AO21x2_ASAP7_75t_L g4285 ( 
.A1(n_4137),
.A2(n_297),
.B(n_298),
.Y(n_4285)
);

BUFx4f_ASAP7_75t_SL g4286 ( 
.A(n_4121),
.Y(n_4286)
);

CKINVDCx5p33_ASAP7_75t_R g4287 ( 
.A(n_4096),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4129),
.Y(n_4288)
);

AOI22xp33_ASAP7_75t_SL g4289 ( 
.A1(n_4108),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_4289)
);

BUFx4_ASAP7_75t_R g4290 ( 
.A(n_4156),
.Y(n_4290)
);

HB1xp67_ASAP7_75t_SL g4291 ( 
.A(n_4121),
.Y(n_4291)
);

BUFx10_ASAP7_75t_L g4292 ( 
.A(n_4093),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4160),
.Y(n_4293)
);

AOI22xp33_ASAP7_75t_SL g4294 ( 
.A1(n_4120),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_4294)
);

CKINVDCx11_ASAP7_75t_R g4295 ( 
.A(n_4112),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4075),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4054),
.B(n_4015),
.Y(n_4297)
);

BUFx3_ASAP7_75t_L g4298 ( 
.A(n_4079),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4069),
.A2(n_302),
.B(n_303),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4100),
.Y(n_4300)
);

NAND2x1p5_ASAP7_75t_L g4301 ( 
.A(n_4085),
.B(n_303),
.Y(n_4301)
);

INVx3_ASAP7_75t_L g4302 ( 
.A(n_4079),
.Y(n_4302)
);

CKINVDCx20_ASAP7_75t_R g4303 ( 
.A(n_4036),
.Y(n_4303)
);

OAI21x1_ASAP7_75t_L g4304 ( 
.A1(n_4044),
.A2(n_304),
.B(n_305),
.Y(n_4304)
);

BUFx8_ASAP7_75t_L g4305 ( 
.A(n_4132),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4160),
.Y(n_4306)
);

AO21x1_ASAP7_75t_SL g4307 ( 
.A1(n_4074),
.A2(n_306),
.B(n_307),
.Y(n_4307)
);

BUFx12f_ASAP7_75t_L g4308 ( 
.A(n_4127),
.Y(n_4308)
);

INVx2_ASAP7_75t_SL g4309 ( 
.A(n_4165),
.Y(n_4309)
);

AND2x4_ASAP7_75t_L g4310 ( 
.A(n_4165),
.B(n_307),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4120),
.Y(n_4311)
);

AOI21x1_ASAP7_75t_L g4312 ( 
.A1(n_4134),
.A2(n_308),
.B(n_310),
.Y(n_4312)
);

OAI21x1_ASAP7_75t_L g4313 ( 
.A1(n_4073),
.A2(n_308),
.B(n_311),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4059),
.Y(n_4314)
);

AO21x1_ASAP7_75t_SL g4315 ( 
.A1(n_4135),
.A2(n_312),
.B(n_313),
.Y(n_4315)
);

AO21x2_ASAP7_75t_L g4316 ( 
.A1(n_4189),
.A2(n_4138),
.B(n_4155),
.Y(n_4316)
);

OAI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_4174),
.A2(n_4153),
.B(n_4022),
.Y(n_4317)
);

INVxp67_ASAP7_75t_SL g4318 ( 
.A(n_4280),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4177),
.B(n_4302),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_4274),
.A2(n_4095),
.B1(n_4098),
.B2(n_4139),
.Y(n_4320)
);

INVx4_ASAP7_75t_L g4321 ( 
.A(n_4185),
.Y(n_4321)
);

AO21x2_ASAP7_75t_L g4322 ( 
.A1(n_4311),
.A2(n_4150),
.B(n_4152),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4293),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4176),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_4203),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4181),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4186),
.Y(n_4327)
);

INVx3_ASAP7_75t_L g4328 ( 
.A(n_4195),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4203),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4187),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4306),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4177),
.B(n_4130),
.Y(n_4332)
);

BUFx2_ASAP7_75t_SL g4333 ( 
.A(n_4206),
.Y(n_4333)
);

A2O1A1Ixp33_ASAP7_75t_L g4334 ( 
.A1(n_4249),
.A2(n_4122),
.B(n_4067),
.C(n_4103),
.Y(n_4334)
);

OR2x6_ASAP7_75t_L g4335 ( 
.A(n_4224),
.B(n_4087),
.Y(n_4335)
);

INVx3_ASAP7_75t_L g4336 ( 
.A(n_4205),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4190),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4198),
.Y(n_4338)
);

INVx3_ASAP7_75t_L g4339 ( 
.A(n_4205),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4200),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4207),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4225),
.Y(n_4342)
);

BUFx2_ASAP7_75t_L g4343 ( 
.A(n_4246),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_4216),
.Y(n_4344)
);

INVxp67_ASAP7_75t_L g4345 ( 
.A(n_4291),
.Y(n_4345)
);

HB1xp67_ASAP7_75t_L g4346 ( 
.A(n_4192),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4226),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4208),
.Y(n_4348)
);

BUFx2_ASAP7_75t_L g4349 ( 
.A(n_4202),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4244),
.A2(n_4146),
.B1(n_4164),
.B2(n_4162),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_SL g4351 ( 
.A1(n_4170),
.A2(n_4141),
.B1(n_4145),
.B2(n_4114),
.Y(n_4351)
);

HB1xp67_ASAP7_75t_L g4352 ( 
.A(n_4252),
.Y(n_4352)
);

AOI21x1_ASAP7_75t_L g4353 ( 
.A1(n_4273),
.A2(n_4125),
.B(n_4118),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4211),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4217),
.Y(n_4355)
);

AOI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4236),
.A2(n_4053),
.B(n_4047),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4253),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4261),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4251),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4263),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4199),
.B(n_4056),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4304),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4228),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4232),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4264),
.Y(n_4365)
);

CKINVDCx11_ASAP7_75t_R g4366 ( 
.A(n_4201),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4247),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4266),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4250),
.Y(n_4369)
);

INVxp33_ASAP7_75t_L g4370 ( 
.A(n_4185),
.Y(n_4370)
);

HB1xp67_ASAP7_75t_L g4371 ( 
.A(n_4219),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4309),
.Y(n_4372)
);

BUFx3_ASAP7_75t_L g4373 ( 
.A(n_4170),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_4260),
.Y(n_4374)
);

BUFx3_ASAP7_75t_L g4375 ( 
.A(n_4170),
.Y(n_4375)
);

INVx4_ASAP7_75t_L g4376 ( 
.A(n_4205),
.Y(n_4376)
);

OAI21x1_ASAP7_75t_L g4377 ( 
.A1(n_4191),
.A2(n_4197),
.B(n_4194),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4220),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4221),
.Y(n_4379)
);

CKINVDCx6p67_ASAP7_75t_R g4380 ( 
.A(n_4278),
.Y(n_4380)
);

INVxp33_ASAP7_75t_L g4381 ( 
.A(n_4167),
.Y(n_4381)
);

AOI211xp5_ASAP7_75t_L g4382 ( 
.A1(n_4243),
.A2(n_4105),
.B(n_4142),
.C(n_4056),
.Y(n_4382)
);

OAI22xp5_ASAP7_75t_L g4383 ( 
.A1(n_4214),
.A2(n_4081),
.B1(n_4056),
.B2(n_314),
.Y(n_4383)
);

AND2x2_ASAP7_75t_L g4384 ( 
.A(n_4188),
.B(n_312),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4256),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4258),
.Y(n_4386)
);

AND2x4_ASAP7_75t_L g4387 ( 
.A(n_4278),
.B(n_313),
.Y(n_4387)
);

HB1xp67_ASAP7_75t_L g4388 ( 
.A(n_4268),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4269),
.Y(n_4389)
);

AO21x2_ASAP7_75t_L g4390 ( 
.A1(n_4270),
.A2(n_315),
.B(n_316),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4229),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_4231),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4242),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4271),
.Y(n_4394)
);

OR2x2_ASAP7_75t_L g4395 ( 
.A(n_4296),
.B(n_4314),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_4255),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_4227),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4282),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4298),
.B(n_315),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_4278),
.Y(n_4400)
);

OR2x2_ASAP7_75t_L g4401 ( 
.A(n_4300),
.B(n_316),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4288),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4275),
.Y(n_4403)
);

OA21x2_ASAP7_75t_L g4404 ( 
.A1(n_4182),
.A2(n_317),
.B(n_318),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4171),
.B(n_317),
.Y(n_4405)
);

AOI22xp33_ASAP7_75t_SL g4406 ( 
.A1(n_4285),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4218),
.Y(n_4407)
);

INVx4_ASAP7_75t_L g4408 ( 
.A(n_4290),
.Y(n_4408)
);

BUFx3_ASAP7_75t_L g4409 ( 
.A(n_4305),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4193),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4168),
.Y(n_4411)
);

HB1xp67_ASAP7_75t_L g4412 ( 
.A(n_4167),
.Y(n_4412)
);

NOR2x1_ASAP7_75t_SL g4413 ( 
.A(n_4277),
.B(n_319),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4230),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4237),
.Y(n_4415)
);

OR2x6_ASAP7_75t_L g4416 ( 
.A(n_4301),
.B(n_321),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4173),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4184),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4213),
.Y(n_4419)
);

INVx3_ASAP7_75t_L g4420 ( 
.A(n_4239),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4175),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4248),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4254),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4259),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4259),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4212),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4234),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4212),
.Y(n_4428)
);

INVx5_ASAP7_75t_L g4429 ( 
.A(n_4284),
.Y(n_4429)
);

BUFx3_ASAP7_75t_L g4430 ( 
.A(n_4305),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4299),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4172),
.Y(n_4432)
);

OAI21x1_ASAP7_75t_L g4433 ( 
.A1(n_4215),
.A2(n_4210),
.B(n_4209),
.Y(n_4433)
);

INVx2_ASAP7_75t_SL g4434 ( 
.A(n_4223),
.Y(n_4434)
);

INVx1_ASAP7_75t_SL g4435 ( 
.A(n_4179),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4310),
.Y(n_4436)
);

BUFx3_ASAP7_75t_L g4437 ( 
.A(n_4284),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4310),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4312),
.Y(n_4439)
);

AO21x2_ASAP7_75t_L g4440 ( 
.A1(n_4265),
.A2(n_321),
.B(n_322),
.Y(n_4440)
);

INVx3_ASAP7_75t_L g4441 ( 
.A(n_4223),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4312),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4234),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4297),
.Y(n_4444)
);

AOI22xp33_ASAP7_75t_L g4445 ( 
.A1(n_4272),
.A2(n_325),
.B1(n_322),
.B2(n_324),
.Y(n_4445)
);

HB1xp67_ASAP7_75t_SL g4446 ( 
.A(n_4238),
.Y(n_4446)
);

AND2x4_ASAP7_75t_L g4447 ( 
.A(n_4180),
.B(n_4196),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4313),
.Y(n_4448)
);

BUFx3_ASAP7_75t_L g4449 ( 
.A(n_4283),
.Y(n_4449)
);

AOI22xp33_ASAP7_75t_L g4450 ( 
.A1(n_4281),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4238),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4183),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4279),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4235),
.B(n_330),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4233),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4303),
.B(n_330),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4222),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4279),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_4295),
.Y(n_4459)
);

INVx2_ASAP7_75t_L g4460 ( 
.A(n_4286),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4276),
.Y(n_4461)
);

BUFx3_ASAP7_75t_L g4462 ( 
.A(n_4308),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4196),
.Y(n_4463)
);

NAND3xp33_ASAP7_75t_L g4464 ( 
.A(n_4317),
.B(n_4289),
.C(n_4294),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4376),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4351),
.B(n_4257),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4352),
.Y(n_4467)
);

AOI222xp33_ASAP7_75t_L g4468 ( 
.A1(n_4461),
.A2(n_4241),
.B1(n_4262),
.B2(n_4240),
.C1(n_4292),
.C2(n_4287),
.Y(n_4468)
);

OAI22xp33_ASAP7_75t_L g4469 ( 
.A1(n_4408),
.A2(n_4267),
.B1(n_4307),
.B2(n_4178),
.Y(n_4469)
);

AND2x2_ASAP7_75t_SL g4470 ( 
.A(n_4408),
.B(n_4204),
.Y(n_4470)
);

AOI22xp33_ASAP7_75t_L g4471 ( 
.A1(n_4316),
.A2(n_4245),
.B1(n_4315),
.B2(n_4307),
.Y(n_4471)
);

INVx3_ASAP7_75t_L g4472 ( 
.A(n_4376),
.Y(n_4472)
);

OR2x2_ASAP7_75t_L g4473 ( 
.A(n_4444),
.B(n_4169),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_4345),
.Y(n_4474)
);

OAI211xp5_ASAP7_75t_L g4475 ( 
.A1(n_4356),
.A2(n_4315),
.B(n_4292),
.C(n_333),
.Y(n_4475)
);

BUFx6f_ASAP7_75t_L g4476 ( 
.A(n_4366),
.Y(n_4476)
);

OAI221xp5_ASAP7_75t_L g4477 ( 
.A1(n_4356),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.C(n_334),
.Y(n_4477)
);

OAI211xp5_ASAP7_75t_L g4478 ( 
.A1(n_4334),
.A2(n_331),
.B(n_334),
.C(n_335),
.Y(n_4478)
);

NAND2x1_ASAP7_75t_L g4479 ( 
.A(n_4336),
.B(n_335),
.Y(n_4479)
);

AOI22xp33_ASAP7_75t_L g4480 ( 
.A1(n_4316),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_4480)
);

AOI22xp33_ASAP7_75t_L g4481 ( 
.A1(n_4383),
.A2(n_4432),
.B1(n_4447),
.B2(n_4320),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_L g4482 ( 
.A(n_4435),
.B(n_336),
.Y(n_4482)
);

OAI21xp5_ASAP7_75t_L g4483 ( 
.A1(n_4334),
.A2(n_339),
.B(n_340),
.Y(n_4483)
);

AOI22xp33_ASAP7_75t_L g4484 ( 
.A1(n_4447),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_4484)
);

AOI221xp5_ASAP7_75t_L g4485 ( 
.A1(n_4381),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.C(n_345),
.Y(n_4485)
);

OAI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4345),
.A2(n_344),
.B1(n_347),
.B2(n_349),
.Y(n_4486)
);

AOI22xp33_ASAP7_75t_L g4487 ( 
.A1(n_4320),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_4487)
);

AOI22xp33_ASAP7_75t_SL g4488 ( 
.A1(n_4373),
.A2(n_350),
.B1(n_351),
.B2(n_353),
.Y(n_4488)
);

AOI22xp33_ASAP7_75t_SL g4489 ( 
.A1(n_4373),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_4489)
);

OAI22xp33_ASAP7_75t_L g4490 ( 
.A1(n_4381),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_4490)
);

NOR2x1_ASAP7_75t_L g4491 ( 
.A(n_4375),
.B(n_4400),
.Y(n_4491)
);

AOI22xp33_ASAP7_75t_SL g4492 ( 
.A1(n_4375),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4352),
.Y(n_4493)
);

AOI221xp5_ASAP7_75t_L g4494 ( 
.A1(n_4382),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.C(n_360),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_4380),
.A2(n_359),
.B1(n_361),
.B2(n_363),
.Y(n_4495)
);

AOI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_4444),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_4496)
);

OAI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_4349),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_4497)
);

OAI221xp5_ASAP7_75t_L g4498 ( 
.A1(n_4351),
.A2(n_4350),
.B1(n_4406),
.B2(n_4400),
.C(n_4335),
.Y(n_4498)
);

AOI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_4439),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_4415),
.B(n_367),
.Y(n_4500)
);

AOI21xp33_ASAP7_75t_L g4501 ( 
.A1(n_4322),
.A2(n_368),
.B(n_369),
.Y(n_4501)
);

AOI21xp33_ASAP7_75t_L g4502 ( 
.A1(n_4322),
.A2(n_370),
.B(n_372),
.Y(n_4502)
);

OAI221xp5_ASAP7_75t_L g4503 ( 
.A1(n_4350),
.A2(n_370),
.B1(n_374),
.B2(n_375),
.C(n_376),
.Y(n_4503)
);

OR2x2_ASAP7_75t_L g4504 ( 
.A(n_4359),
.B(n_374),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_4446),
.A2(n_375),
.B1(n_376),
.B2(n_378),
.Y(n_4505)
);

AOI221xp5_ASAP7_75t_L g4506 ( 
.A1(n_4439),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.C(n_381),
.Y(n_4506)
);

OR2x2_ASAP7_75t_L g4507 ( 
.A(n_4359),
.B(n_379),
.Y(n_4507)
);

BUFx12f_ASAP7_75t_L g4508 ( 
.A(n_4366),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4448),
.B(n_380),
.Y(n_4509)
);

AOI22xp33_ASAP7_75t_SL g4510 ( 
.A1(n_4413),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_4510)
);

AOI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4440),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_4511)
);

AOI22xp33_ASAP7_75t_SL g4512 ( 
.A1(n_4412),
.A2(n_387),
.B1(n_389),
.B2(n_390),
.Y(n_4512)
);

AOI22xp33_ASAP7_75t_L g4513 ( 
.A1(n_4440),
.A2(n_387),
.B1(n_389),
.B2(n_391),
.Y(n_4513)
);

OA21x2_ASAP7_75t_L g4514 ( 
.A1(n_4318),
.A2(n_392),
.B(n_393),
.Y(n_4514)
);

AOI22xp5_ASAP7_75t_L g4515 ( 
.A1(n_4452),
.A2(n_392),
.B1(n_394),
.B2(n_395),
.Y(n_4515)
);

AOI221xp5_ASAP7_75t_L g4516 ( 
.A1(n_4442),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.C(n_397),
.Y(n_4516)
);

OAI21xp33_ASAP7_75t_L g4517 ( 
.A1(n_4406),
.A2(n_396),
.B(n_397),
.Y(n_4517)
);

AOI221xp5_ASAP7_75t_L g4518 ( 
.A1(n_4442),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.C(n_401),
.Y(n_4518)
);

OAI22xp5_ASAP7_75t_L g4519 ( 
.A1(n_4446),
.A2(n_398),
.B1(n_399),
.B2(n_401),
.Y(n_4519)
);

AOI22xp33_ASAP7_75t_SL g4520 ( 
.A1(n_4412),
.A2(n_402),
.B1(n_403),
.B2(n_405),
.Y(n_4520)
);

NAND3xp33_ASAP7_75t_L g4521 ( 
.A(n_4450),
.B(n_402),
.C(n_403),
.Y(n_4521)
);

AOI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4390),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_4333),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4364),
.Y(n_4524)
);

O2A1O1Ixp33_ASAP7_75t_L g4525 ( 
.A1(n_4416),
.A2(n_406),
.B(n_407),
.C(n_408),
.Y(n_4525)
);

OR2x6_ASAP7_75t_L g4526 ( 
.A(n_4416),
.B(n_409),
.Y(n_4526)
);

AOI22xp33_ASAP7_75t_L g4527 ( 
.A1(n_4390),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_4527)
);

OAI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_4429),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_4528)
);

HB1xp67_ASAP7_75t_L g4529 ( 
.A(n_4346),
.Y(n_4529)
);

INVxp67_ASAP7_75t_L g4530 ( 
.A(n_4387),
.Y(n_4530)
);

AO21x2_ASAP7_75t_L g4531 ( 
.A1(n_4318),
.A2(n_413),
.B(n_414),
.Y(n_4531)
);

AOI22xp33_ASAP7_75t_L g4532 ( 
.A1(n_4319),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_4532)
);

OAI22xp5_ASAP7_75t_L g4533 ( 
.A1(n_4429),
.A2(n_415),
.B1(n_416),
.B2(n_419),
.Y(n_4533)
);

OAI21x1_ASAP7_75t_SL g4534 ( 
.A1(n_4436),
.A2(n_420),
.B(n_421),
.Y(n_4534)
);

OAI22xp5_ASAP7_75t_L g4535 ( 
.A1(n_4429),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_4535)
);

INVx5_ASAP7_75t_SL g4536 ( 
.A(n_4416),
.Y(n_4536)
);

NOR2xp33_ASAP7_75t_L g4537 ( 
.A(n_4370),
.B(n_422),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4420),
.B(n_424),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4364),
.Y(n_4539)
);

AOI22xp33_ASAP7_75t_L g4540 ( 
.A1(n_4420),
.A2(n_4460),
.B1(n_4455),
.B2(n_4459),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4324),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4326),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4327),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4448),
.B(n_425),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4330),
.Y(n_4545)
);

OR2x2_ASAP7_75t_L g4546 ( 
.A(n_4395),
.B(n_426),
.Y(n_4546)
);

CKINVDCx20_ASAP7_75t_R g4547 ( 
.A(n_4397),
.Y(n_4547)
);

OA21x2_ASAP7_75t_L g4548 ( 
.A1(n_4377),
.A2(n_426),
.B(n_427),
.Y(n_4548)
);

AOI22xp33_ASAP7_75t_L g4549 ( 
.A1(n_4460),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4332),
.B(n_429),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4405),
.B(n_4443),
.Y(n_4551)
);

OAI22xp5_ASAP7_75t_L g4552 ( 
.A1(n_4429),
.A2(n_430),
.B1(n_431),
.B2(n_434),
.Y(n_4552)
);

OAI221xp5_ASAP7_75t_L g4553 ( 
.A1(n_4335),
.A2(n_431),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4459),
.Y(n_4554)
);

INVx4_ASAP7_75t_SL g4555 ( 
.A(n_4409),
.Y(n_4555)
);

AOI21xp5_ASAP7_75t_L g4556 ( 
.A1(n_4456),
.A2(n_435),
.B(n_436),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_4456),
.A2(n_438),
.B(n_439),
.Y(n_4557)
);

AOI22xp33_ASAP7_75t_L g4558 ( 
.A1(n_4343),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_4558)
);

INVx4_ASAP7_75t_SL g4559 ( 
.A(n_4409),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_4449),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_4560)
);

AOI22xp33_ASAP7_75t_SL g4561 ( 
.A1(n_4433),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4325),
.B(n_443),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4329),
.B(n_444),
.Y(n_4563)
);

AND2x4_ASAP7_75t_L g4564 ( 
.A(n_4336),
.B(n_445),
.Y(n_4564)
);

AOI21xp33_ASAP7_75t_L g4565 ( 
.A1(n_4422),
.A2(n_446),
.B(n_447),
.Y(n_4565)
);

BUFx3_ASAP7_75t_L g4566 ( 
.A(n_4430),
.Y(n_4566)
);

AOI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_4449),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4337),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4436),
.B(n_448),
.Y(n_4569)
);

AOI22xp33_ASAP7_75t_L g4570 ( 
.A1(n_4431),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_4570)
);

AOI221xp5_ASAP7_75t_L g4571 ( 
.A1(n_4426),
.A2(n_450),
.B1(n_451),
.B2(n_453),
.C(n_454),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4340),
.Y(n_4572)
);

AOI221xp5_ASAP7_75t_L g4573 ( 
.A1(n_4428),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.C(n_457),
.Y(n_4573)
);

OAI221xp5_ASAP7_75t_L g4574 ( 
.A1(n_4335),
.A2(n_455),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_4574)
);

OAI221xp5_ASAP7_75t_L g4575 ( 
.A1(n_4450),
.A2(n_458),
.B1(n_459),
.B2(n_460),
.C(n_461),
.Y(n_4575)
);

AOI222xp33_ASAP7_75t_L g4576 ( 
.A1(n_4445),
.A2(n_4387),
.B1(n_4431),
.B2(n_4362),
.C1(n_4346),
.C2(n_4430),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4341),
.Y(n_4577)
);

OAI22xp5_ASAP7_75t_L g4578 ( 
.A1(n_4437),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4438),
.B(n_462),
.Y(n_4579)
);

OAI221xp5_ASAP7_75t_L g4580 ( 
.A1(n_4339),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.C(n_466),
.Y(n_4580)
);

AO21x1_ASAP7_75t_L g4581 ( 
.A1(n_4463),
.A2(n_463),
.B(n_465),
.Y(n_4581)
);

AOI22xp33_ASAP7_75t_L g4582 ( 
.A1(n_4418),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.Y(n_4582)
);

OR2x2_ASAP7_75t_L g4583 ( 
.A(n_4403),
.B(n_467),
.Y(n_4583)
);

AOI221xp5_ASAP7_75t_L g4584 ( 
.A1(n_4362),
.A2(n_4410),
.B1(n_4414),
.B2(n_4445),
.C(n_4371),
.Y(n_4584)
);

AOI22xp5_ASAP7_75t_L g4585 ( 
.A1(n_4374),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_4585)
);

OAI211xp5_ASAP7_75t_L g4586 ( 
.A1(n_4339),
.A2(n_471),
.B(n_472),
.C(n_473),
.Y(n_4586)
);

AOI22xp33_ASAP7_75t_L g4587 ( 
.A1(n_4457),
.A2(n_473),
.B1(n_474),
.B2(n_475),
.Y(n_4587)
);

OAI211xp5_ASAP7_75t_L g4588 ( 
.A1(n_4353),
.A2(n_474),
.B(n_475),
.C(n_476),
.Y(n_4588)
);

AOI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4370),
.A2(n_476),
.B(n_477),
.Y(n_4589)
);

BUFx3_ASAP7_75t_L g4590 ( 
.A(n_4344),
.Y(n_4590)
);

AOI222xp33_ASAP7_75t_L g4591 ( 
.A1(n_4462),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.C1(n_482),
.C2(n_483),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4438),
.B(n_479),
.Y(n_4592)
);

CKINVDCx20_ASAP7_75t_R g4593 ( 
.A(n_4392),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4371),
.Y(n_4594)
);

BUFx6f_ASAP7_75t_L g4595 ( 
.A(n_4321),
.Y(n_4595)
);

AO21x2_ASAP7_75t_L g4596 ( 
.A1(n_4407),
.A2(n_480),
.B(n_481),
.Y(n_4596)
);

AOI221xp5_ASAP7_75t_L g4597 ( 
.A1(n_4388),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.C(n_487),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4342),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4474),
.B(n_4421),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4470),
.B(n_4411),
.Y(n_4600)
);

BUFx2_ASAP7_75t_L g4601 ( 
.A(n_4508),
.Y(n_4601)
);

INVxp67_ASAP7_75t_L g4602 ( 
.A(n_4491),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4529),
.Y(n_4603)
);

HB1xp67_ASAP7_75t_L g4604 ( 
.A(n_4530),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4595),
.Y(n_4605)
);

BUFx8_ASAP7_75t_L g4606 ( 
.A(n_4476),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4554),
.B(n_4451),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4594),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4576),
.B(n_4481),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4467),
.Y(n_4610)
);

HB1xp67_ASAP7_75t_L g4611 ( 
.A(n_4514),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4540),
.B(n_4465),
.Y(n_4612)
);

BUFx2_ASAP7_75t_R g4613 ( 
.A(n_4523),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4493),
.Y(n_4614)
);

BUFx3_ASAP7_75t_L g4615 ( 
.A(n_4476),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4472),
.B(n_4536),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4472),
.B(n_4411),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4524),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4536),
.B(n_4417),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4548),
.B(n_4417),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4539),
.B(n_4388),
.Y(n_4621)
);

INVx2_ASAP7_75t_SL g4622 ( 
.A(n_4595),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4548),
.B(n_4361),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4595),
.Y(n_4624)
);

BUFx3_ASAP7_75t_L g4625 ( 
.A(n_4476),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4566),
.Y(n_4626)
);

INVx2_ASAP7_75t_L g4627 ( 
.A(n_4479),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4514),
.Y(n_4628)
);

OR2x2_ASAP7_75t_L g4629 ( 
.A(n_4546),
.B(n_4338),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_4596),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4561),
.B(n_4441),
.Y(n_4631)
);

BUFx3_ASAP7_75t_L g4632 ( 
.A(n_4590),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4541),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4555),
.B(n_4441),
.Y(n_4634)
);

BUFx2_ASAP7_75t_L g4635 ( 
.A(n_4526),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4542),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4494),
.B(n_4451),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4555),
.B(n_4372),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4543),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4559),
.B(n_4391),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4545),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4531),
.Y(n_4642)
);

AND2x2_ASAP7_75t_SL g4643 ( 
.A(n_4466),
.B(n_4321),
.Y(n_4643)
);

NOR2xp33_ASAP7_75t_L g4644 ( 
.A(n_4559),
.B(n_4462),
.Y(n_4644)
);

AND2x4_ASAP7_75t_L g4645 ( 
.A(n_4473),
.B(n_4437),
.Y(n_4645)
);

INVx2_ASAP7_75t_L g4646 ( 
.A(n_4564),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4568),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4564),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4572),
.Y(n_4649)
);

INVxp67_ASAP7_75t_L g4650 ( 
.A(n_4526),
.Y(n_4650)
);

OR2x2_ASAP7_75t_L g4651 ( 
.A(n_4598),
.B(n_4338),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4551),
.B(n_4391),
.Y(n_4652)
);

AND2x4_ASAP7_75t_SL g4653 ( 
.A(n_4471),
.B(n_4453),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4577),
.Y(n_4654)
);

AND2x4_ASAP7_75t_SL g4655 ( 
.A(n_4538),
.B(n_4453),
.Y(n_4655)
);

NOR2xp33_ASAP7_75t_R g4656 ( 
.A(n_4593),
.B(n_4401),
.Y(n_4656)
);

AND2x4_ASAP7_75t_L g4657 ( 
.A(n_4483),
.B(n_4328),
.Y(n_4657)
);

NOR2x1_ASAP7_75t_SL g4658 ( 
.A(n_4475),
.B(n_4434),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4550),
.B(n_4393),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4504),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4569),
.B(n_4393),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4468),
.B(n_4443),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4583),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4507),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4579),
.B(n_4396),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4509),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4592),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4464),
.B(n_4424),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4500),
.Y(n_4669)
);

BUFx6f_ASAP7_75t_L g4670 ( 
.A(n_4562),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4563),
.B(n_4396),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4534),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4584),
.B(n_4423),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4544),
.B(n_4589),
.Y(n_4674)
);

AND2x4_ASAP7_75t_SL g4675 ( 
.A(n_4547),
.B(n_4458),
.Y(n_4675)
);

INVx2_ASAP7_75t_L g4676 ( 
.A(n_4498),
.Y(n_4676)
);

BUFx3_ASAP7_75t_L g4677 ( 
.A(n_4537),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4581),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4501),
.B(n_4323),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4522),
.Y(n_4680)
);

BUFx2_ASAP7_75t_L g4681 ( 
.A(n_4469),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4588),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4502),
.B(n_4323),
.Y(n_4683)
);

INVx3_ASAP7_75t_L g4684 ( 
.A(n_4478),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4477),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4490),
.Y(n_4686)
);

BUFx2_ASAP7_75t_L g4687 ( 
.A(n_4505),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4482),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4528),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4519),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4533),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4553),
.Y(n_4692)
);

BUFx3_ASAP7_75t_L g4693 ( 
.A(n_4515),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4480),
.B(n_4331),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4535),
.Y(n_4695)
);

BUFx3_ASAP7_75t_L g4696 ( 
.A(n_4585),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4574),
.Y(n_4697)
);

HB1xp67_ASAP7_75t_L g4698 ( 
.A(n_4552),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4525),
.Y(n_4699)
);

INVxp67_ASAP7_75t_SL g4700 ( 
.A(n_4556),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4510),
.B(n_4331),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4503),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4484),
.B(n_4425),
.Y(n_4703)
);

INVx2_ASAP7_75t_SL g4704 ( 
.A(n_4486),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4511),
.B(n_4427),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4604),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4621),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4615),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4634),
.B(n_4328),
.Y(n_4709)
);

OR2x2_ASAP7_75t_L g4710 ( 
.A(n_4642),
.B(n_4357),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4615),
.Y(n_4711)
);

HB1xp67_ASAP7_75t_L g4712 ( 
.A(n_4635),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4634),
.B(n_4363),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4616),
.B(n_4363),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4621),
.Y(n_4715)
);

NAND2x1_ASAP7_75t_L g4716 ( 
.A(n_4642),
.B(n_4367),
.Y(n_4716)
);

BUFx3_ASAP7_75t_L g4717 ( 
.A(n_4606),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4684),
.B(n_4557),
.Y(n_4718)
);

NAND4xp25_ASAP7_75t_L g4719 ( 
.A(n_4609),
.B(n_4487),
.C(n_4591),
.D(n_4485),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4625),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4616),
.B(n_4367),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4627),
.B(n_4378),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4611),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4627),
.B(n_4379),
.Y(n_4724)
);

OAI21xp33_ASAP7_75t_SL g4725 ( 
.A1(n_4628),
.A2(n_4527),
.B(n_4513),
.Y(n_4725)
);

AND2x2_ASAP7_75t_L g4726 ( 
.A(n_4675),
.B(n_4385),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4628),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4651),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4675),
.B(n_4386),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4626),
.B(n_4389),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4626),
.B(n_4394),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4651),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4629),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4638),
.B(n_4398),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4625),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4629),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4670),
.Y(n_4737)
);

INVx2_ASAP7_75t_SL g4738 ( 
.A(n_4606),
.Y(n_4738)
);

AOI22xp33_ASAP7_75t_L g4739 ( 
.A1(n_4681),
.A2(n_4517),
.B1(n_4521),
.B2(n_4575),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4670),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4638),
.B(n_4402),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4603),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4670),
.Y(n_4743)
);

AND2x4_ASAP7_75t_L g4744 ( 
.A(n_4622),
.B(n_4419),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4660),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4678),
.B(n_4358),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4660),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4684),
.B(n_4497),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4684),
.B(n_4384),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4670),
.Y(n_4750)
);

INVxp33_ASAP7_75t_L g4751 ( 
.A(n_4644),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4622),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4599),
.B(n_4360),
.Y(n_4753)
);

AOI22xp33_ASAP7_75t_L g4754 ( 
.A1(n_4681),
.A2(n_4499),
.B1(n_4506),
.B2(n_4516),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4599),
.B(n_4600),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4664),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4600),
.B(n_4365),
.Y(n_4757)
);

INVx2_ASAP7_75t_SL g4758 ( 
.A(n_4606),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4650),
.B(n_4512),
.Y(n_4759)
);

AOI22xp33_ASAP7_75t_SL g4760 ( 
.A1(n_4653),
.A2(n_4586),
.B1(n_4580),
.B2(n_4578),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4601),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4664),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4601),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_L g4764 ( 
.A(n_4658),
.B(n_4520),
.Y(n_4764)
);

HB1xp67_ASAP7_75t_L g4765 ( 
.A(n_4646),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_4645),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4663),
.Y(n_4767)
);

OR2x2_ASAP7_75t_L g4768 ( 
.A(n_4667),
.B(n_4368),
.Y(n_4768)
);

AND2x4_ASAP7_75t_L g4769 ( 
.A(n_4602),
.B(n_4419),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4645),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4755),
.B(n_4643),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4765),
.Y(n_4772)
);

AOI22xp5_ASAP7_75t_L g4773 ( 
.A1(n_4754),
.A2(n_4676),
.B1(n_4687),
.B2(n_4680),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4755),
.B(n_4643),
.Y(n_4774)
);

INVx3_ASAP7_75t_L g4775 ( 
.A(n_4716),
.Y(n_4775)
);

INVxp67_ASAP7_75t_L g4776 ( 
.A(n_4717),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4723),
.Y(n_4777)
);

CKINVDCx6p67_ASAP7_75t_R g4778 ( 
.A(n_4717),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4716),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4761),
.B(n_4687),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4766),
.Y(n_4781)
);

NOR2xp33_ASAP7_75t_L g4782 ( 
.A(n_4751),
.B(n_4613),
.Y(n_4782)
);

INVx4_ASAP7_75t_L g4783 ( 
.A(n_4738),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4723),
.Y(n_4784)
);

AND2x2_ASAP7_75t_L g4785 ( 
.A(n_4761),
.B(n_4612),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4763),
.B(n_4612),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4763),
.B(n_4646),
.Y(n_4787)
);

INVx2_ASAP7_75t_SL g4788 ( 
.A(n_4738),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4766),
.Y(n_4789)
);

INVx3_ASAP7_75t_L g4790 ( 
.A(n_4770),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4727),
.Y(n_4791)
);

BUFx2_ASAP7_75t_L g4792 ( 
.A(n_4737),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4770),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4708),
.B(n_4648),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4708),
.B(n_4711),
.Y(n_4795)
);

BUFx2_ASAP7_75t_L g4796 ( 
.A(n_4737),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4740),
.Y(n_4797)
);

INVx2_ASAP7_75t_L g4798 ( 
.A(n_4740),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4711),
.B(n_4682),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4743),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4720),
.B(n_4648),
.Y(n_4801)
);

HB1xp67_ASAP7_75t_L g4802 ( 
.A(n_4712),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4727),
.Y(n_4803)
);

OR2x2_ASAP7_75t_L g4804 ( 
.A(n_4706),
.B(n_4630),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4728),
.Y(n_4805)
);

AOI22xp33_ASAP7_75t_L g4806 ( 
.A1(n_4719),
.A2(n_4676),
.B1(n_4693),
.B2(n_4657),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4728),
.Y(n_4807)
);

INVx3_ASAP7_75t_L g4808 ( 
.A(n_4744),
.Y(n_4808)
);

OR2x2_ASAP7_75t_L g4809 ( 
.A(n_4748),
.B(n_4607),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_L g4810 ( 
.A(n_4751),
.B(n_4758),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4720),
.B(n_4619),
.Y(n_4811)
);

INVx4_ASAP7_75t_L g4812 ( 
.A(n_4758),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4732),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4735),
.B(n_4619),
.Y(n_4814)
);

AO21x2_ASAP7_75t_L g4815 ( 
.A1(n_4718),
.A2(n_4700),
.B(n_4673),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4735),
.B(n_4605),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4709),
.B(n_4605),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4743),
.Y(n_4818)
);

INVx5_ASAP7_75t_SL g4819 ( 
.A(n_4750),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4750),
.Y(n_4820)
);

CKINVDCx11_ASAP7_75t_R g4821 ( 
.A(n_4752),
.Y(n_4821)
);

AND2x4_ASAP7_75t_L g4822 ( 
.A(n_4752),
.B(n_4645),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4709),
.Y(n_4823)
);

INVx1_ASAP7_75t_SL g4824 ( 
.A(n_4726),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4732),
.Y(n_4825)
);

AND2x2_ASAP7_75t_L g4826 ( 
.A(n_4726),
.B(n_4624),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4815),
.B(n_4739),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_SL g4828 ( 
.A(n_4773),
.B(n_4760),
.Y(n_4828)
);

NAND2x1p5_ASAP7_75t_L g4829 ( 
.A(n_4783),
.B(n_4632),
.Y(n_4829)
);

NOR2xp33_ASAP7_75t_SL g4830 ( 
.A(n_4771),
.B(n_4688),
.Y(n_4830)
);

OR2x2_ASAP7_75t_L g4831 ( 
.A(n_4780),
.B(n_4759),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4808),
.Y(n_4832)
);

AND2x2_ASAP7_75t_L g4833 ( 
.A(n_4778),
.B(n_4632),
.Y(n_4833)
);

AND2x2_ASAP7_75t_L g4834 ( 
.A(n_4778),
.B(n_4655),
.Y(n_4834)
);

BUFx2_ASAP7_75t_L g4835 ( 
.A(n_4808),
.Y(n_4835)
);

OR2x2_ASAP7_75t_L g4836 ( 
.A(n_4824),
.B(n_4749),
.Y(n_4836)
);

NAND3xp33_ASAP7_75t_L g4837 ( 
.A(n_4806),
.B(n_4725),
.C(n_4764),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4771),
.B(n_4655),
.Y(n_4838)
);

INVx2_ASAP7_75t_L g4839 ( 
.A(n_4808),
.Y(n_4839)
);

AND2x4_ASAP7_75t_L g4840 ( 
.A(n_4822),
.B(n_4624),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4774),
.B(n_4672),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4792),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4774),
.B(n_4672),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4792),
.Y(n_4844)
);

NAND2x1_ASAP7_75t_L g4845 ( 
.A(n_4822),
.B(n_4744),
.Y(n_4845)
);

NAND2x1p5_ASAP7_75t_L g4846 ( 
.A(n_4783),
.B(n_4756),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4796),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4796),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4785),
.B(n_4653),
.Y(n_4849)
);

CKINVDCx14_ASAP7_75t_R g4850 ( 
.A(n_4821),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4815),
.B(n_4680),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4775),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4815),
.B(n_4698),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4775),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4785),
.B(n_4729),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4786),
.B(n_4729),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4775),
.Y(n_4857)
);

OR2x6_ASAP7_75t_L g4858 ( 
.A(n_4783),
.B(n_4688),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4790),
.Y(n_4859)
);

OR2x2_ASAP7_75t_L g4860 ( 
.A(n_4802),
.B(n_4704),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4790),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4812),
.B(n_4699),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4790),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_4786),
.B(n_4631),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4787),
.Y(n_4865)
);

BUFx3_ASAP7_75t_L g4866 ( 
.A(n_4822),
.Y(n_4866)
);

OR2x2_ASAP7_75t_L g4867 ( 
.A(n_4799),
.B(n_4704),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4819),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4811),
.B(n_4631),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_4811),
.B(n_4667),
.Y(n_4870)
);

INVxp67_ASAP7_75t_L g4871 ( 
.A(n_4810),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4787),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4781),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4835),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4832),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4869),
.B(n_4788),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4866),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4832),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4866),
.Y(n_4879)
);

BUFx2_ASAP7_75t_L g4880 ( 
.A(n_4850),
.Y(n_4880)
);

NOR2xp33_ASAP7_75t_L g4881 ( 
.A(n_4850),
.B(n_4776),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4839),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4846),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4839),
.Y(n_4884)
);

INVx5_ASAP7_75t_L g4885 ( 
.A(n_4858),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_4846),
.Y(n_4886)
);

BUFx2_ASAP7_75t_L g4887 ( 
.A(n_4829),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4842),
.Y(n_4888)
);

AND2x4_ASAP7_75t_L g4889 ( 
.A(n_4844),
.B(n_4823),
.Y(n_4889)
);

INVx1_ASAP7_75t_SL g4890 ( 
.A(n_4849),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4864),
.B(n_4817),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4833),
.B(n_4817),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4855),
.B(n_4788),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4856),
.B(n_4826),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4834),
.B(n_4826),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4847),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4840),
.B(n_4812),
.Y(n_4897)
);

AND2x2_ASAP7_75t_SL g4898 ( 
.A(n_4827),
.B(n_4782),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4848),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4841),
.B(n_4812),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4843),
.B(n_4814),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4859),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4838),
.B(n_4814),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4829),
.B(n_4795),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4845),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4870),
.B(n_4795),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4840),
.B(n_4816),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4861),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4885),
.B(n_4794),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4880),
.B(n_4794),
.Y(n_4910)
);

BUFx2_ASAP7_75t_L g4911 ( 
.A(n_4880),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4892),
.B(n_4801),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4885),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4885),
.B(n_4801),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_L g4915 ( 
.A(n_4885),
.B(n_4863),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4892),
.B(n_4816),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4885),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4891),
.B(n_4823),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4891),
.B(n_4871),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4876),
.B(n_4858),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4906),
.Y(n_4921)
);

AOI211x1_ASAP7_75t_L g4922 ( 
.A1(n_4897),
.A2(n_4828),
.B(n_4827),
.C(n_4837),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4906),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4907),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4894),
.B(n_4865),
.Y(n_4925)
);

OR2x2_ASAP7_75t_L g4926 ( 
.A(n_4893),
.B(n_4858),
.Y(n_4926)
);

AND2x2_ASAP7_75t_L g4927 ( 
.A(n_4894),
.B(n_4871),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4895),
.B(n_4903),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4907),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4901),
.B(n_4872),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4901),
.Y(n_4931)
);

BUFx3_ASAP7_75t_L g4932 ( 
.A(n_4887),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4889),
.Y(n_4933)
);

AOI22xp33_ASAP7_75t_L g4934 ( 
.A1(n_4898),
.A2(n_4828),
.B1(n_4673),
.B2(n_4851),
.Y(n_4934)
);

AND2x2_ASAP7_75t_L g4935 ( 
.A(n_4895),
.B(n_4677),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4889),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4889),
.B(n_4772),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4874),
.B(n_4860),
.Y(n_4938)
);

INVxp67_ASAP7_75t_L g4939 ( 
.A(n_4911),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4933),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4936),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4910),
.B(n_4900),
.Y(n_4942)
);

NAND4xp25_ASAP7_75t_L g4943 ( 
.A(n_4934),
.B(n_4881),
.C(n_4830),
.D(n_4890),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4928),
.B(n_4900),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4916),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4909),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4932),
.Y(n_4947)
);

AOI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4934),
.A2(n_4903),
.B1(n_4702),
.B2(n_4898),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4912),
.B(n_4819),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4909),
.Y(n_4950)
);

NAND2x1p5_ASAP7_75t_L g4951 ( 
.A(n_4935),
.B(n_4904),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4914),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4914),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4937),
.Y(n_4954)
);

NAND2x1_ASAP7_75t_SL g4955 ( 
.A(n_4927),
.B(n_4904),
.Y(n_4955)
);

AND2x2_ASAP7_75t_L g4956 ( 
.A(n_4919),
.B(n_4877),
.Y(n_4956)
);

INVx2_ASAP7_75t_SL g4957 ( 
.A(n_4932),
.Y(n_4957)
);

NOR2x1_ASAP7_75t_L g4958 ( 
.A(n_4937),
.B(n_4887),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4918),
.Y(n_4959)
);

INVxp67_ASAP7_75t_L g4960 ( 
.A(n_4925),
.Y(n_4960)
);

OR3x2_ASAP7_75t_L g4961 ( 
.A(n_4938),
.B(n_4831),
.C(n_4836),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4957),
.B(n_4819),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4958),
.Y(n_4963)
);

INVx2_ASAP7_75t_L g4964 ( 
.A(n_4951),
.Y(n_4964)
);

INVx1_ASAP7_75t_SL g4965 ( 
.A(n_4955),
.Y(n_4965)
);

NAND2xp33_ASAP7_75t_R g4966 ( 
.A(n_4956),
.B(n_4868),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4944),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4942),
.Y(n_4968)
);

INVx4_ASAP7_75t_L g4969 ( 
.A(n_4947),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4945),
.B(n_4931),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4959),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4943),
.B(n_4939),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_4948),
.B(n_4877),
.Y(n_4973)
);

AND2x4_ASAP7_75t_L g4974 ( 
.A(n_4949),
.B(n_4921),
.Y(n_4974)
);

NAND2xp33_ASAP7_75t_SL g4975 ( 
.A(n_4940),
.B(n_4853),
.Y(n_4975)
);

AND2x4_ASAP7_75t_L g4976 ( 
.A(n_4941),
.B(n_4905),
.Y(n_4976)
);

CKINVDCx8_ASAP7_75t_R g4977 ( 
.A(n_4961),
.Y(n_4977)
);

OR2x2_ASAP7_75t_L g4978 ( 
.A(n_4960),
.B(n_4853),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4950),
.Y(n_4979)
);

OR2x2_ASAP7_75t_L g4980 ( 
.A(n_4965),
.B(n_4851),
.Y(n_4980)
);

OAI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4977),
.A2(n_4922),
.B1(n_4662),
.B2(n_4693),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4976),
.B(n_4819),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4976),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4970),
.B(n_4923),
.Y(n_4984)
);

NAND3xp33_ASAP7_75t_L g4985 ( 
.A(n_4963),
.B(n_4868),
.C(n_4905),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4964),
.Y(n_4986)
);

OR2x2_ASAP7_75t_L g4987 ( 
.A(n_4962),
.B(n_4772),
.Y(n_4987)
);

INVx2_ASAP7_75t_L g4988 ( 
.A(n_4969),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4973),
.B(n_4879),
.Y(n_4989)
);

OAI22xp5_ASAP7_75t_L g4990 ( 
.A1(n_4967),
.A2(n_4668),
.B1(n_4696),
.B2(n_4867),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4978),
.Y(n_4991)
);

NAND2x1_ASAP7_75t_L g4992 ( 
.A(n_4979),
.B(n_4883),
.Y(n_4992)
);

INVxp67_ASAP7_75t_SL g4993 ( 
.A(n_4966),
.Y(n_4993)
);

INVxp67_ASAP7_75t_SL g4994 ( 
.A(n_4982),
.Y(n_4994)
);

AOI22xp33_ASAP7_75t_L g4995 ( 
.A1(n_4986),
.A2(n_4924),
.B1(n_4929),
.B2(n_4862),
.Y(n_4995)
);

OAI211xp5_ASAP7_75t_SL g4996 ( 
.A1(n_4989),
.A2(n_4968),
.B(n_4920),
.C(n_4926),
.Y(n_4996)
);

OAI32xp33_ASAP7_75t_L g4997 ( 
.A1(n_4980),
.A2(n_4804),
.A3(n_4925),
.B1(n_4930),
.B2(n_4862),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4984),
.Y(n_4998)
);

OAI21xp33_ASAP7_75t_L g4999 ( 
.A1(n_4981),
.A2(n_4972),
.B(n_4809),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4983),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4993),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4992),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4990),
.B(n_4879),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4988),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4991),
.B(n_4875),
.Y(n_5005)
);

OA21x2_ASAP7_75t_L g5006 ( 
.A1(n_4985),
.A2(n_4913),
.B(n_4915),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4987),
.B(n_4974),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4984),
.Y(n_5008)
);

NOR2xp33_ASAP7_75t_L g5009 ( 
.A(n_4983),
.B(n_4930),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4984),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_5006),
.Y(n_5011)
);

OR2x2_ASAP7_75t_L g5012 ( 
.A(n_4998),
.B(n_4809),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_5006),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_5002),
.Y(n_5014)
);

OAI22xp33_ASAP7_75t_L g5015 ( 
.A1(n_5000),
.A2(n_4804),
.B1(n_4883),
.B2(n_4886),
.Y(n_5015)
);

INVxp67_ASAP7_75t_L g5016 ( 
.A(n_5009),
.Y(n_5016)
);

NAND3xp33_ASAP7_75t_L g5017 ( 
.A(n_4995),
.B(n_4975),
.C(n_4886),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_5008),
.Y(n_5018)
);

INVx2_ASAP7_75t_L g5019 ( 
.A(n_5010),
.Y(n_5019)
);

O2A1O1Ixp33_ASAP7_75t_L g5020 ( 
.A1(n_4997),
.A2(n_4915),
.B(n_4917),
.C(n_4954),
.Y(n_5020)
);

OAI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_5001),
.A2(n_4896),
.B(n_4888),
.Y(n_5021)
);

INVx1_ASAP7_75t_SL g5022 ( 
.A(n_5007),
.Y(n_5022)
);

NOR3xp33_ASAP7_75t_L g5023 ( 
.A(n_4996),
.B(n_4971),
.C(n_4952),
.Y(n_5023)
);

AOI21xp5_ASAP7_75t_L g5024 ( 
.A1(n_5005),
.A2(n_4950),
.B(n_4946),
.Y(n_5024)
);

XNOR2xp5_ASAP7_75t_L g5025 ( 
.A(n_5004),
.B(n_4899),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_5003),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4994),
.Y(n_5027)
);

OAI22xp33_ASAP7_75t_L g5028 ( 
.A1(n_4999),
.A2(n_4793),
.B1(n_4789),
.B2(n_4781),
.Y(n_5028)
);

OAI21xp33_ASAP7_75t_L g5029 ( 
.A1(n_4999),
.A2(n_4793),
.B(n_4789),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_5006),
.Y(n_5030)
);

AOI22xp33_ASAP7_75t_L g5031 ( 
.A1(n_4998),
.A2(n_4745),
.B1(n_4762),
.B2(n_4747),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_5009),
.A2(n_4882),
.B(n_4878),
.Y(n_5032)
);

INVx2_ASAP7_75t_L g5033 ( 
.A(n_5006),
.Y(n_5033)
);

AOI32xp33_ASAP7_75t_L g5034 ( 
.A1(n_4996),
.A2(n_4800),
.A3(n_4818),
.B1(n_4820),
.B2(n_4797),
.Y(n_5034)
);

CKINVDCx20_ASAP7_75t_R g5035 ( 
.A(n_4998),
.Y(n_5035)
);

OR2x2_ASAP7_75t_L g5036 ( 
.A(n_4998),
.B(n_4756),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_5012),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_5034),
.B(n_4884),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_5028),
.B(n_4873),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_5015),
.B(n_4902),
.Y(n_5040)
);

AOI22xp5_ASAP7_75t_L g5041 ( 
.A1(n_5035),
.A2(n_5022),
.B1(n_5023),
.B2(n_5019),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_5036),
.Y(n_5042)
);

OR2x2_ASAP7_75t_L g5043 ( 
.A(n_5017),
.B(n_4797),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_5031),
.B(n_4908),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_5018),
.B(n_4767),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_SL g5046 ( 
.A(n_5029),
.B(n_4798),
.Y(n_5046)
);

NOR2xp33_ASAP7_75t_L g5047 ( 
.A(n_5014),
.B(n_4953),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_5025),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_5021),
.B(n_4798),
.Y(n_5049)
);

NOR2x1_ASAP7_75t_L g5050 ( 
.A(n_5011),
.B(n_4852),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_5024),
.B(n_4800),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_5032),
.B(n_4818),
.Y(n_5052)
);

NOR2x1_ASAP7_75t_L g5053 ( 
.A(n_5013),
.B(n_4852),
.Y(n_5053)
);

NOR2xp33_ASAP7_75t_L g5054 ( 
.A(n_5016),
.B(n_4820),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_5020),
.B(n_4805),
.Y(n_5055)
);

AND2x4_ASAP7_75t_L g5056 ( 
.A(n_5027),
.B(n_4854),
.Y(n_5056)
);

NOR2xp33_ASAP7_75t_L g5057 ( 
.A(n_5026),
.B(n_5030),
.Y(n_5057)
);

NAND3x1_ASAP7_75t_L g5058 ( 
.A(n_5033),
.B(n_4784),
.C(n_4777),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_5034),
.B(n_4805),
.Y(n_5059)
);

AOI22xp33_ASAP7_75t_L g5060 ( 
.A1(n_5023),
.A2(n_4715),
.B1(n_4707),
.B2(n_4742),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_5034),
.B(n_4807),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5034),
.B(n_4807),
.Y(n_5062)
);

INVx1_ASAP7_75t_SL g5063 ( 
.A(n_5012),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_5034),
.B(n_4813),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_5012),
.Y(n_5065)
);

NOR3xp33_ASAP7_75t_SL g5066 ( 
.A(n_5040),
.B(n_4784),
.C(n_4777),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_5055),
.Y(n_5067)
);

XNOR2x2_ASAP7_75t_L g5068 ( 
.A(n_5050),
.B(n_5053),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_5056),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_5056),
.B(n_4813),
.Y(n_5070)
);

NAND2x1_ASAP7_75t_L g5071 ( 
.A(n_5052),
.B(n_4854),
.Y(n_5071)
);

AOI211xp5_ASAP7_75t_L g5072 ( 
.A1(n_5047),
.A2(n_4857),
.B(n_4825),
.C(n_4803),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5043),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5051),
.Y(n_5074)
);

INVx1_ASAP7_75t_SL g5075 ( 
.A(n_5063),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_5049),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_5060),
.B(n_4825),
.Y(n_5077)
);

NAND3xp33_ASAP7_75t_SL g5078 ( 
.A(n_5041),
.B(n_4857),
.C(n_4803),
.Y(n_5078)
);

INVx2_ASAP7_75t_SL g5079 ( 
.A(n_5045),
.Y(n_5079)
);

XNOR2xp5_ASAP7_75t_L g5080 ( 
.A(n_5048),
.B(n_4677),
.Y(n_5080)
);

NAND2xp33_ASAP7_75t_R g5081 ( 
.A(n_5037),
.B(n_4791),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_5059),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5061),
.Y(n_5083)
);

NOR4xp25_ASAP7_75t_SL g5084 ( 
.A(n_5046),
.B(n_4791),
.C(n_4733),
.D(n_4736),
.Y(n_5084)
);

INVxp67_ASAP7_75t_L g5085 ( 
.A(n_5054),
.Y(n_5085)
);

AND2x2_ASAP7_75t_L g5086 ( 
.A(n_5065),
.B(n_4734),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_5042),
.B(n_4669),
.Y(n_5087)
);

OR2x2_ASAP7_75t_L g5088 ( 
.A(n_5038),
.B(n_5044),
.Y(n_5088)
);

AOI21xp33_ASAP7_75t_L g5089 ( 
.A1(n_5057),
.A2(n_4779),
.B(n_4710),
.Y(n_5089)
);

XNOR2xp5_ASAP7_75t_L g5090 ( 
.A(n_5058),
.B(n_4666),
.Y(n_5090)
);

OAI21xp33_ASAP7_75t_L g5091 ( 
.A1(n_5039),
.A2(n_4779),
.B(n_4721),
.Y(n_5091)
);

BUFx6f_ASAP7_75t_L g5092 ( 
.A(n_5069),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_5086),
.B(n_5062),
.Y(n_5093)
);

AOI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_5075),
.A2(n_5064),
.B1(n_4714),
.B2(n_4721),
.Y(n_5094)
);

AOI22xp5_ASAP7_75t_L g5095 ( 
.A1(n_5091),
.A2(n_4714),
.B1(n_4769),
.B2(n_4640),
.Y(n_5095)
);

OAI21xp33_ASAP7_75t_L g5096 ( 
.A1(n_5080),
.A2(n_4746),
.B(n_4640),
.Y(n_5096)
);

OAI21xp33_ASAP7_75t_SL g5097 ( 
.A1(n_5070),
.A2(n_4710),
.B(n_4746),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_5071),
.A2(n_4674),
.B(n_4637),
.Y(n_5098)
);

OA22x2_ASAP7_75t_L g5099 ( 
.A1(n_5090),
.A2(n_4769),
.B1(n_4608),
.B2(n_4610),
.Y(n_5099)
);

OAI21xp5_ASAP7_75t_L g5100 ( 
.A1(n_5085),
.A2(n_4618),
.B(n_4614),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_L g5101 ( 
.A(n_5072),
.B(n_4685),
.Y(n_5101)
);

NOR2x1_ASAP7_75t_L g5102 ( 
.A(n_5078),
.B(n_4696),
.Y(n_5102)
);

INVxp67_ASAP7_75t_SL g5103 ( 
.A(n_5081),
.Y(n_5103)
);

AND2x2_ASAP7_75t_L g5104 ( 
.A(n_5079),
.B(n_5077),
.Y(n_5104)
);

INVx1_ASAP7_75t_SL g5105 ( 
.A(n_5068),
.Y(n_5105)
);

NOR3xp33_ASAP7_75t_SL g5106 ( 
.A(n_5073),
.B(n_4695),
.C(n_4689),
.Y(n_5106)
);

AOI21xp5_ASAP7_75t_L g5107 ( 
.A1(n_5089),
.A2(n_4692),
.B(n_4697),
.Y(n_5107)
);

AOI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_5076),
.A2(n_4769),
.B1(n_4734),
.B2(n_4741),
.Y(n_5108)
);

INVx2_ASAP7_75t_SL g5109 ( 
.A(n_5087),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_5066),
.Y(n_5110)
);

INVx2_ASAP7_75t_L g5111 ( 
.A(n_5099),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_5108),
.Y(n_5112)
);

OAI31xp33_ASAP7_75t_L g5113 ( 
.A1(n_5105),
.A2(n_5067),
.A3(n_5083),
.B(n_5082),
.Y(n_5113)
);

NAND3xp33_ASAP7_75t_L g5114 ( 
.A(n_5092),
.B(n_5074),
.C(n_5088),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_5103),
.A2(n_5084),
.B(n_4692),
.Y(n_5115)
);

HB1xp67_ASAP7_75t_L g5116 ( 
.A(n_5102),
.Y(n_5116)
);

O2A1O1Ixp5_ASAP7_75t_L g5117 ( 
.A1(n_5101),
.A2(n_4744),
.B(n_4713),
.C(n_4724),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5094),
.Y(n_5118)
);

INVx1_ASAP7_75t_SL g5119 ( 
.A(n_5092),
.Y(n_5119)
);

AOI22xp5_ASAP7_75t_L g5120 ( 
.A1(n_5096),
.A2(n_4741),
.B1(n_4713),
.B2(n_4731),
.Y(n_5120)
);

AOI322xp5_ASAP7_75t_L g5121 ( 
.A1(n_5106),
.A2(n_4657),
.A3(n_4685),
.B1(n_4702),
.B2(n_4697),
.C1(n_4730),
.C2(n_4731),
.Y(n_5121)
);

AOI31xp33_ASAP7_75t_L g5122 ( 
.A1(n_5093),
.A2(n_4691),
.A3(n_4690),
.B(n_4657),
.Y(n_5122)
);

AOI221xp5_ASAP7_75t_L g5123 ( 
.A1(n_5098),
.A2(n_4636),
.B1(n_4647),
.B2(n_4641),
.C(n_4639),
.Y(n_5123)
);

OAI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_5107),
.A2(n_4730),
.B(n_4724),
.Y(n_5124)
);

XNOR2xp5_ASAP7_75t_L g5125 ( 
.A(n_5095),
.B(n_4690),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5097),
.Y(n_5126)
);

NOR3x1_ASAP7_75t_L g5127 ( 
.A(n_5114),
.B(n_5110),
.C(n_5109),
.Y(n_5127)
);

AOI31xp33_ASAP7_75t_L g5128 ( 
.A1(n_5119),
.A2(n_5104),
.A3(n_5100),
.B(n_4686),
.Y(n_5128)
);

AOI21xp33_ASAP7_75t_L g5129 ( 
.A1(n_5126),
.A2(n_4768),
.B(n_4654),
.Y(n_5129)
);

CKINVDCx20_ASAP7_75t_R g5130 ( 
.A(n_5125),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_R g5131 ( 
.A(n_5118),
.B(n_484),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_5117),
.Y(n_5132)
);

OAI211xp5_ASAP7_75t_SL g5133 ( 
.A1(n_5113),
.A2(n_4649),
.B(n_4633),
.C(n_4768),
.Y(n_5133)
);

NAND4xp25_ASAP7_75t_SL g5134 ( 
.A(n_5115),
.B(n_4722),
.C(n_4757),
.D(n_4753),
.Y(n_5134)
);

OAI221xp5_ASAP7_75t_L g5135 ( 
.A1(n_5124),
.A2(n_5120),
.B1(n_5112),
.B2(n_5116),
.C(n_5111),
.Y(n_5135)
);

AOI222xp33_ASAP7_75t_L g5136 ( 
.A1(n_5123),
.A2(n_4722),
.B1(n_4757),
.B2(n_4753),
.C1(n_4683),
.C2(n_4679),
.Y(n_5136)
);

OAI222xp33_ASAP7_75t_L g5137 ( 
.A1(n_5121),
.A2(n_4617),
.B1(n_4623),
.B2(n_4683),
.C1(n_4679),
.C2(n_4620),
.Y(n_5137)
);

AOI221x1_ASAP7_75t_L g5138 ( 
.A1(n_5122),
.A2(n_4617),
.B1(n_4623),
.B2(n_4652),
.C(n_4620),
.Y(n_5138)
);

INVxp67_ASAP7_75t_SL g5139 ( 
.A(n_5115),
.Y(n_5139)
);

AOI22xp5_ASAP7_75t_L g5140 ( 
.A1(n_5119),
.A2(n_4652),
.B1(n_4701),
.B2(n_4705),
.Y(n_5140)
);

O2A1O1Ixp33_ASAP7_75t_L g5141 ( 
.A1(n_5116),
.A2(n_4701),
.B(n_4565),
.C(n_4705),
.Y(n_5141)
);

OAI211xp5_ASAP7_75t_L g5142 ( 
.A1(n_5113),
.A2(n_4656),
.B(n_4488),
.C(n_4489),
.Y(n_5142)
);

NOR2xp33_ASAP7_75t_L g5143 ( 
.A(n_5125),
.B(n_4659),
.Y(n_5143)
);

AOI221x1_ASAP7_75t_L g5144 ( 
.A1(n_5114),
.A2(n_4703),
.B1(n_4694),
.B2(n_4665),
.C(n_4661),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_SL g5145 ( 
.A(n_5131),
.B(n_4656),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_L g5146 ( 
.A(n_5140),
.B(n_5142),
.Y(n_5146)
);

NAND2xp33_ASAP7_75t_L g5147 ( 
.A(n_5132),
.B(n_4661),
.Y(n_5147)
);

NOR2xp33_ASAP7_75t_L g5148 ( 
.A(n_5128),
.B(n_4659),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_5143),
.B(n_4665),
.Y(n_5149)
);

OAI22xp5_ASAP7_75t_L g5150 ( 
.A1(n_5130),
.A2(n_5135),
.B1(n_5139),
.B2(n_5141),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5133),
.Y(n_5151)
);

NOR3xp33_ASAP7_75t_L g5152 ( 
.A(n_5129),
.B(n_4492),
.C(n_4597),
.Y(n_5152)
);

INVxp67_ASAP7_75t_L g5153 ( 
.A(n_5134),
.Y(n_5153)
);

NOR3xp33_ASAP7_75t_L g5154 ( 
.A(n_5127),
.B(n_4518),
.C(n_4573),
.Y(n_5154)
);

NOR2xp67_ASAP7_75t_L g5155 ( 
.A(n_5144),
.B(n_486),
.Y(n_5155)
);

NAND4xp75_ASAP7_75t_L g5156 ( 
.A(n_5138),
.B(n_4571),
.C(n_4694),
.D(n_4703),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_SL g5157 ( 
.A(n_5136),
.B(n_4671),
.Y(n_5157)
);

NOR2xp33_ASAP7_75t_L g5158 ( 
.A(n_5137),
.B(n_4671),
.Y(n_5158)
);

OAI21xp5_ASAP7_75t_L g5159 ( 
.A1(n_5128),
.A2(n_4558),
.B(n_4560),
.Y(n_5159)
);

NAND3xp33_ASAP7_75t_L g5160 ( 
.A(n_5132),
.B(n_4567),
.C(n_4495),
.Y(n_5160)
);

NOR3x2_ASAP7_75t_L g5161 ( 
.A(n_5127),
.B(n_487),
.C(n_488),
.Y(n_5161)
);

NAND4xp25_ASAP7_75t_L g5162 ( 
.A(n_5146),
.B(n_4549),
.C(n_4570),
.D(n_4532),
.Y(n_5162)
);

NAND4xp25_ASAP7_75t_L g5163 ( 
.A(n_5148),
.B(n_4582),
.C(n_4587),
.D(n_4496),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_5154),
.B(n_4454),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5149),
.B(n_4399),
.Y(n_5165)
);

OR2x2_ASAP7_75t_L g5166 ( 
.A(n_5160),
.B(n_4404),
.Y(n_5166)
);

INVxp67_ASAP7_75t_L g5167 ( 
.A(n_5147),
.Y(n_5167)
);

NOR3xp33_ASAP7_75t_L g5168 ( 
.A(n_5150),
.B(n_489),
.C(n_490),
.Y(n_5168)
);

OA211x2_ASAP7_75t_L g5169 ( 
.A1(n_5153),
.A2(n_489),
.B(n_491),
.C(n_492),
.Y(n_5169)
);

NOR2xp67_ASAP7_75t_L g5170 ( 
.A(n_5145),
.B(n_491),
.Y(n_5170)
);

OAI211xp5_ASAP7_75t_SL g5171 ( 
.A1(n_5151),
.A2(n_492),
.B(n_494),
.C(n_495),
.Y(n_5171)
);

NOR4xp25_ASAP7_75t_L g5172 ( 
.A(n_5157),
.B(n_4355),
.C(n_4354),
.D(n_4348),
.Y(n_5172)
);

AOI22xp5_ASAP7_75t_L g5173 ( 
.A1(n_5168),
.A2(n_5158),
.B1(n_5155),
.B2(n_5156),
.Y(n_5173)
);

INVxp67_ASAP7_75t_L g5174 ( 
.A(n_5170),
.Y(n_5174)
);

XNOR2xp5_ASAP7_75t_L g5175 ( 
.A(n_5169),
.B(n_5161),
.Y(n_5175)
);

NOR2x1_ASAP7_75t_L g5176 ( 
.A(n_5171),
.B(n_5166),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5165),
.Y(n_5177)
);

INVx2_ASAP7_75t_L g5178 ( 
.A(n_5164),
.Y(n_5178)
);

NOR2x2_ASAP7_75t_L g5179 ( 
.A(n_5178),
.B(n_5167),
.Y(n_5179)
);

NOR3xp33_ASAP7_75t_L g5180 ( 
.A(n_5174),
.B(n_5159),
.C(n_5162),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5175),
.B(n_5172),
.Y(n_5181)
);

AND2x2_ASAP7_75t_SL g5182 ( 
.A(n_5180),
.B(n_5177),
.Y(n_5182)
);

OAI22xp5_ASAP7_75t_SL g5183 ( 
.A1(n_5181),
.A2(n_5173),
.B1(n_5176),
.B2(n_5152),
.Y(n_5183)
);

A2O1A1Ixp33_ASAP7_75t_L g5184 ( 
.A1(n_5182),
.A2(n_5179),
.B(n_5163),
.C(n_496),
.Y(n_5184)
);

AOI22xp5_ASAP7_75t_L g5185 ( 
.A1(n_5184),
.A2(n_5183),
.B1(n_4404),
.B2(n_4347),
.Y(n_5185)
);

AOI22xp5_ASAP7_75t_L g5186 ( 
.A1(n_5185),
.A2(n_4404),
.B1(n_4369),
.B2(n_496),
.Y(n_5186)
);

HB1xp67_ASAP7_75t_L g5187 ( 
.A(n_5186),
.Y(n_5187)
);

INVx3_ASAP7_75t_L g5188 ( 
.A(n_5187),
.Y(n_5188)
);

OR2x2_ASAP7_75t_L g5189 ( 
.A(n_5188),
.B(n_494),
.Y(n_5189)
);

AOI22xp5_ASAP7_75t_L g5190 ( 
.A1(n_5189),
.A2(n_495),
.B1(n_497),
.B2(n_498),
.Y(n_5190)
);

AOI22xp5_ASAP7_75t_L g5191 ( 
.A1(n_5190),
.A2(n_497),
.B1(n_499),
.B2(n_500),
.Y(n_5191)
);

OAI22xp33_ASAP7_75t_L g5192 ( 
.A1(n_5191),
.A2(n_502),
.B1(n_503),
.B2(n_505),
.Y(n_5192)
);

OAI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_5192),
.A2(n_502),
.B1(n_503),
.B2(n_505),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5193),
.Y(n_5194)
);

AOI21xp5_ASAP7_75t_L g5195 ( 
.A1(n_5194),
.A2(n_506),
.B(n_507),
.Y(n_5195)
);

AOI221xp5_ASAP7_75t_L g5196 ( 
.A1(n_5195),
.A2(n_506),
.B1(n_507),
.B2(n_508),
.C(n_509),
.Y(n_5196)
);

OAI221xp5_ASAP7_75t_L g5197 ( 
.A1(n_5195),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.C(n_511),
.Y(n_5197)
);

AOI22xp5_ASAP7_75t_L g5198 ( 
.A1(n_5197),
.A2(n_5196),
.B1(n_511),
.B2(n_512),
.Y(n_5198)
);

AOI211xp5_ASAP7_75t_L g5199 ( 
.A1(n_5198),
.A2(n_510),
.B(n_513),
.C(n_514),
.Y(n_5199)
);


endmodule