module fake_jpeg_19641_n_378 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_52),
.Y(n_82)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_0),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_60),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_33),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_90),
.B1(n_104),
.B2(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_26),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_92),
.B(n_28),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_38),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_46),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_93),
.B1(n_97),
.B2(n_57),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_20),
.B1(n_27),
.B2(n_51),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_99),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_56),
.Y(n_142)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_58),
.C(n_60),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_121),
.C(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_117),
.Y(n_166)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_111),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_94),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_130),
.B1(n_69),
.B2(n_67),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_16),
.B1(n_28),
.B2(n_29),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_64),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_143),
.B1(n_85),
.B2(n_69),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_65),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_28),
.C(n_26),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_42),
.B1(n_47),
.B2(n_44),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_141),
.B1(n_86),
.B2(n_79),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_57),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_47),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_28),
.B1(n_29),
.B2(n_13),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_76),
.B(n_12),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_135),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_91),
.B(n_11),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_138),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_93),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_79),
.B(n_11),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_59),
.B1(n_34),
.B2(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_85),
.Y(n_152)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_75),
.B(n_10),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_146),
.A2(n_151),
.B1(n_169),
.B2(n_171),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_57),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_153),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_106),
.B1(n_143),
.B2(n_122),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_168),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_103),
.B(n_3),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_124),
.B(n_105),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_94),
.B1(n_77),
.B2(n_34),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_110),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_112),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_117),
.A2(n_77),
.B1(n_88),
.B2(n_56),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_1),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_172),
.B(n_176),
.CI(n_145),
.CON(n_183),
.SN(n_183)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_109),
.A2(n_141),
.B1(n_124),
.B2(n_106),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_9),
.B1(n_10),
.B2(n_6),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_15),
.C(n_14),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_118),
.A3(n_111),
.B1(n_108),
.B2(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_182),
.A2(n_189),
.B(n_193),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_184),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_191),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_217),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_107),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_192),
.B(n_205),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_107),
.B(n_105),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_122),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_144),
.B(n_3),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_206),
.B1(n_209),
.B2(n_171),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_129),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_129),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_158),
.C(n_175),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_1),
.B(n_4),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_112),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_150),
.A2(n_137),
.B1(n_133),
.B2(n_5),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_14),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_14),
.Y(n_208)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_151),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_11),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_214),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_155),
.B1(n_159),
.B2(n_181),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_4),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_164),
.A2(n_148),
.B1(n_146),
.B2(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_223),
.C(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_146),
.B1(n_169),
.B2(n_177),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_239),
.B1(n_251),
.B2(n_184),
.Y(n_265)
);

AO21x2_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_153),
.B(n_177),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_170),
.C(n_172),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_248),
.C(n_183),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_247),
.B1(n_187),
.B2(n_202),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_172),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_238),
.Y(n_270)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_176),
.A3(n_155),
.B1(n_156),
.B2(n_159),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_193),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_176),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_156),
.B1(n_159),
.B2(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_210),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_181),
.B1(n_163),
.B2(n_179),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_5),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_203),
.A2(n_179),
.B1(n_7),
.B2(n_8),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_255),
.A2(n_266),
.B(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_220),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_262),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_189),
.B1(n_193),
.B2(n_212),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_265),
.B1(n_235),
.B2(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_231),
.B(n_188),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_183),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_192),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_185),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_273),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_277),
.B1(n_255),
.B2(n_245),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_223),
.B(n_197),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_230),
.C(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_279),
.C(n_280),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_191),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_213),
.B(n_215),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_276),
.B(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_278),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_215),
.B1(n_182),
.B2(n_187),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_228),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_223),
.C(n_226),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_288),
.B1(n_295),
.B2(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_226),
.C(n_236),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_215),
.B(n_208),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_248),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_292),
.B1(n_265),
.B2(n_199),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_232),
.C(n_205),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_276),
.B1(n_269),
.B2(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_232),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_294),
.B1(n_271),
.B2(n_257),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_237),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g298 ( 
.A1(n_260),
.A2(n_251),
.B(n_239),
.C(n_225),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_298),
.A2(n_254),
.B(n_253),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_228),
.B1(n_227),
.B2(n_207),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_240),
.C(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_267),
.B1(n_277),
.B2(n_257),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_314),
.B1(n_317),
.B2(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_274),
.C(n_211),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_275),
.B1(n_261),
.B2(n_254),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_244),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_316),
.Y(n_330)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_281),
.B(n_214),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_320),
.B(n_295),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_253),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_299),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_206),
.B1(n_219),
.B2(n_216),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_218),
.B1(n_219),
.B2(n_183),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_294),
.B1(n_293),
.B2(n_296),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_285),
.C(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_328),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_285),
.C(n_287),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_331),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_291),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_296),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_336),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_303),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_340),
.B(n_344),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_320),
.B1(n_313),
.B2(n_317),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_343),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_314),
.B1(n_304),
.B2(n_319),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_342),
.A2(n_348),
.B1(n_327),
.B2(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_329),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_307),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_316),
.B(n_289),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_335),
.B(n_337),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_336),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_325),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_351),
.B(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_358),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_354),
.A2(n_359),
.B(n_350),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_328),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_359),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_349),
.B(n_5),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_357),
.B(n_338),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_186),
.C(n_7),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_186),
.C(n_8),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_SL g360 ( 
.A(n_352),
.B(n_348),
.C(n_342),
.Y(n_360)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_360),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_338),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_366),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_362),
.B(n_358),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_368),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_355),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_365),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_373),
.B(n_370),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_372),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_376),
.B(n_369),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_351),
.Y(n_378)
);


endmodule