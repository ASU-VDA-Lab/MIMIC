module fake_jpeg_19940_n_325 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_20),
.B1(n_15),
.B2(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_44),
.B1(n_30),
.B2(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_20),
.B1(n_15),
.B2(n_16),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_22),
.B(n_26),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_22),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_57),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_67),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_80),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_66),
.B1(n_46),
.B2(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_20),
.B1(n_15),
.B2(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_83),
.B1(n_48),
.B2(n_46),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_29),
.B1(n_38),
.B2(n_26),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_49),
.B1(n_51),
.B2(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_50),
.B1(n_54),
.B2(n_59),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_89),
.B1(n_34),
.B2(n_52),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_59),
.B1(n_63),
.B2(n_53),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_75),
.B(n_77),
.Y(n_114)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_105),
.B1(n_40),
.B2(n_35),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_62),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_41),
.B(n_29),
.C(n_38),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_87),
.B1(n_95),
.B2(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_78),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_38),
.B(n_17),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_81),
.B(n_74),
.Y(n_106)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_116),
.B(n_26),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_108),
.B1(n_35),
.B2(n_40),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_66),
.B1(n_97),
.B2(n_85),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_69),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_21),
.B(n_18),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_72),
.B(n_77),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_93),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_79),
.B(n_83),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_102),
.B(n_84),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_70),
.B1(n_46),
.B2(n_40),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_132),
.B1(n_135),
.B2(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_78),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_36),
.CI(n_27),
.CON(n_131),
.SN(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_143),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_162),
.B1(n_163),
.B2(n_133),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_101),
.C(n_86),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_108),
.C(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_100),
.B1(n_105),
.B2(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_151),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_145),
.A2(n_154),
.B(n_155),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_29),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_117),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_19),
.B1(n_12),
.B2(n_13),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_160),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_8),
.B(n_10),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_31),
.C(n_32),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_171),
.B(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_12),
.B1(n_23),
.B2(n_34),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_40),
.B1(n_35),
.B2(n_12),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_167),
.B1(n_132),
.B2(n_135),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_106),
.A2(n_21),
.B(n_18),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_21),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_35),
.B1(n_23),
.B2(n_45),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_45),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_21),
.B(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_180),
.C(n_181),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_187),
.B(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_131),
.C(n_121),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_131),
.C(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_131),
.B1(n_129),
.B2(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_195),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_112),
.B(n_10),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_45),
.B1(n_25),
.B2(n_24),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_25),
.C(n_24),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_191),
.C(n_76),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_24),
.C(n_45),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_9),
.B(n_10),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_32),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_140),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_144),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_213),
.B(n_225),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_175),
.A2(n_159),
.B1(n_156),
.B2(n_171),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_179),
.B1(n_187),
.B2(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_158),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_152),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_219),
.Y(n_231)
);

AOI21x1_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_152),
.B(n_154),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_194),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_222),
.B1(n_149),
.B2(n_150),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_169),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_150),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_181),
.C(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_237),
.C(n_208),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_233),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_197),
.B(n_183),
.C(n_177),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_204),
.B1(n_219),
.B2(n_210),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_184),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_170),
.C(n_149),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_192),
.B1(n_177),
.B2(n_172),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_208),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_243),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_221),
.A2(n_192),
.B1(n_191),
.B2(n_189),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_222),
.B1(n_216),
.B2(n_207),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_199),
.B1(n_188),
.B2(n_164),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_220),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_157),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_203),
.B(n_211),
.Y(n_247)
);

XOR2x2_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_218),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_265),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_226),
.B(n_241),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_247),
.B(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_257),
.B1(n_260),
.B2(n_234),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_201),
.B1(n_223),
.B2(n_210),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_232),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_210),
.B1(n_163),
.B2(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_220),
.C(n_164),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_32),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_76),
.C(n_14),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_32),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_244),
.B1(n_228),
.B2(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_279),
.B1(n_280),
.B2(n_2),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_269),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_248),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_234),
.C(n_76),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_248),
.C(n_14),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_14),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_0),
.B(n_1),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_255),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_10),
.B1(n_9),
.B2(n_23),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_249),
.B1(n_255),
.B2(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_290),
.B1(n_271),
.B2(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_263),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_287),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_7),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_14),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_0),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_272),
.B(n_277),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_2),
.B(n_3),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_31),
.B(n_14),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_11),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_282),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_270),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

OAI221xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_31),
.B1(n_11),
.B2(n_4),
.C(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_302),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_SL g313 ( 
.A(n_299),
.B(n_301),
.C(n_3),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_11),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_305),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_3),
.C(n_4),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_7),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_311),
.B(n_307),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_294),
.C(n_298),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_3),
.CI(n_4),
.CON(n_312),
.SN(n_312)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_4),
.B(n_5),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_6),
.B(n_7),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_6),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_312),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_309),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_319),
.B(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_306),
.C(n_300),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_314),
.C(n_6),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B1(n_7),
.B2(n_211),
.Y(n_325)
);


endmodule