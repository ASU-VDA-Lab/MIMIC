module fake_ariane_195_n_1754 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1754);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1754;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_75),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_54),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_72),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_19),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_88),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_38),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_94),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_12),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_96),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_137),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_37),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_60),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_27),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_64),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_61),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_54),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_98),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_57),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_66),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_33),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_156),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_83),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_121),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_2),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_140),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_44),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_39),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_51),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_105),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_99),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_89),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_45),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_153),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_31),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_116),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_168),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_166),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_55),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_71),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_76),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_162),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_26),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_126),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_82),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_112),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_15),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_68),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_90),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_17),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_113),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_111),
.Y(n_291)
);

INVxp33_ASAP7_75t_R g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_32),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_158),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_50),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_61),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_142),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_18),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_56),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_131),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_49),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_109),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_13),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_49),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_23),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_40),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_24),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_128),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_167),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_81),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_110),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_115),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_107),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_95),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_7),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_51),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_165),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_77),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_48),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_40),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_143),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_21),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_11),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_85),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_58),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_41),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_55),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_100),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_4),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_28),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_62),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_172),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_336),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_229),
.B(n_1),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_174),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_171),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_182),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_181),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_219),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_175),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_201),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_262),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_180),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_266),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_214),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_229),
.B(n_4),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_183),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_183),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_184),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_219),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_258),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_186),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_186),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_181),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_192),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_204),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_200),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_193),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_271),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_197),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_271),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_223),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_223),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_198),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_205),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_230),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_230),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_195),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_251),
.B(n_6),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_212),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_206),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_176),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_202),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_251),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_271),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_252),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_202),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_252),
.B(n_7),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_249),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_195),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_285),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_207),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_176),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_267),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_249),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_267),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_285),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_268),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_268),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_275),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_209),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_178),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_210),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_275),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_277),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_212),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_216),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_277),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_212),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_218),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_224),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_281),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_281),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_226),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_289),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_231),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_359),
.B(n_227),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_289),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_342),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_354),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_332),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_353),
.B(n_296),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_353),
.B(n_296),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_352),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_362),
.B(n_332),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_364),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_364),
.B(n_314),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_369),
.B(n_314),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_350),
.B(n_317),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_423),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_381),
.B(n_384),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_381),
.B(n_247),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_428),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_343),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_365),
.A2(n_196),
.B1(n_339),
.B2(n_221),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_366),
.A2(n_340),
.B1(n_244),
.B2(n_245),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_408),
.A2(n_318),
.B(n_317),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_410),
.B(n_318),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_357),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_344),
.B(n_215),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_412),
.B(n_177),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_416),
.B(n_247),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_367),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_371),
.Y(n_510)
);

INVx4_ASAP7_75t_SL g511 ( 
.A(n_503),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_358),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_452),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_432),
.A2(n_372),
.B1(n_378),
.B2(n_373),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_452),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_417),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_386),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_452),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_195),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_438),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

AOI22x1_ASAP7_75t_L g528 ( 
.A1(n_437),
.A2(n_462),
.B1(n_486),
.B2(n_447),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

XOR2x2_ASAP7_75t_L g530 ( 
.A(n_482),
.B(n_368),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_453),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_502),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_453),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_417),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_503),
.B(n_195),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_454),
.B(n_346),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_482),
.C(n_393),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_473),
.B(n_505),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_442),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_491),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_503),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_441),
.B(n_387),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_473),
.B(n_374),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_420),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_424),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_465),
.B(n_413),
.C(n_404),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_500),
.B(n_348),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_494),
.A2(n_400),
.B1(n_391),
.B2(n_405),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_461),
.B(n_415),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_457),
.B(n_392),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_480),
.A2(n_414),
.B1(n_394),
.B2(n_419),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_479),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_479),
.B(n_401),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_446),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_479),
.B(n_407),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_424),
.Y(n_568)
);

AND2x2_ASAP7_75t_SL g569 ( 
.A(n_494),
.B(n_305),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_473),
.B(n_399),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_375),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_493),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_461),
.B(n_379),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_461),
.B(n_399),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_461),
.B(n_425),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_437),
.B(n_425),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_472),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_451),
.B(n_383),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_472),
.B(n_178),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_437),
.B(n_427),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_238),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_505),
.B(n_376),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_505),
.B(n_443),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_491),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_458),
.B(n_397),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_451),
.B(n_427),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_493),
.B(n_418),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_492),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_460),
.B(n_403),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_437),
.B(n_321),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_443),
.B(n_179),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_492),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_458),
.B(n_246),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_492),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_460),
.B(n_421),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_503),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_494),
.A2(n_309),
.B1(n_305),
.B2(n_327),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_492),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_468),
.A2(n_321),
.B(n_217),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_437),
.B(n_211),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_496),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_496),
.Y(n_612)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_468),
.A2(n_471),
.B(n_470),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_468),
.B(n_355),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_443),
.B(n_179),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_476),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

BUFx8_ASAP7_75t_SL g621 ( 
.A(n_454),
.Y(n_621)
);

AND3x2_ASAP7_75t_L g622 ( 
.A(n_454),
.B(n_292),
.C(n_196),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_496),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_496),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_496),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_496),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_474),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_471),
.B(n_211),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_447),
.B(n_237),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_458),
.B(n_436),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_474),
.B(n_253),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_458),
.B(n_189),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_475),
.B(n_177),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_494),
.A2(n_327),
.B1(n_309),
.B2(n_339),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_480),
.B(n_300),
.C(n_221),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_503),
.B(n_238),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_475),
.B(n_237),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_475),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_501),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_474),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_447),
.B(n_259),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_447),
.B(n_259),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_260),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_501),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_494),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_447),
.B(n_170),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_501),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_543),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_545),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_507),
.B(n_518),
.Y(n_653)
);

AO221x1_ASAP7_75t_L g654 ( 
.A1(n_649),
.A2(n_477),
.B1(n_177),
.B2(n_334),
.C(n_238),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_534),
.A2(n_494),
.B1(n_503),
.B2(n_439),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_540),
.B(n_447),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_580),
.B(n_576),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_581),
.B(n_462),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_631),
.B(n_462),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_534),
.A2(n_503),
.B1(n_504),
.B2(n_469),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_525),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_550),
.B(n_501),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_563),
.Y(n_664)
);

NAND2x1_ASAP7_75t_L g665 ( 
.A(n_602),
.B(n_503),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_565),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_631),
.B(n_462),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_521),
.B(n_462),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_574),
.B(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_462),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_550),
.B(n_501),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_550),
.B(n_501),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_486),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_510),
.B(n_486),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_556),
.B(n_575),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_569),
.A2(n_504),
.B1(n_439),
.B2(n_499),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_602),
.B(n_501),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_510),
.B(n_486),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_510),
.B(n_486),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_608),
.A2(n_486),
.B(n_483),
.C(n_484),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_558),
.B(n_481),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_566),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_520),
.A2(n_481),
.B(n_483),
.C(n_484),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_571),
.B(n_483),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_591),
.B(n_484),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_574),
.B(n_485),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_537),
.A2(n_485),
.B1(n_487),
.B2(n_488),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_547),
.B(n_485),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_601),
.B(n_487),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_587),
.B(n_488),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_569),
.A2(n_504),
.B1(n_439),
.B2(n_499),
.Y(n_691)
);

BUFx8_ASAP7_75t_L g692 ( 
.A(n_649),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_609),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_629),
.A2(n_489),
.B1(n_495),
.B2(n_498),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_587),
.B(n_489),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_542),
.B(n_489),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_639),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_542),
.B(n_495),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_545),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_552),
.B(n_495),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_552),
.B(n_498),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_594),
.B(n_498),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_615),
.B(n_436),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_535),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_613),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_596),
.B(n_439),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_613),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_512),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_512),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_596),
.B(n_444),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_545),
.B(n_448),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_561),
.B(n_448),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_577),
.A2(n_554),
.B(n_568),
.C(n_553),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_555),
.B(n_449),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_586),
.B(n_444),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_617),
.B(n_444),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_617),
.B(n_633),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_578),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_633),
.B(n_583),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_586),
.B(n_449),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_584),
.B(n_444),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_570),
.B(n_445),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_586),
.B(n_463),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_586),
.B(n_463),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_564),
.B(n_464),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_619),
.B(n_464),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_555),
.B(n_497),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_599),
.B(n_497),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_595),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_570),
.B(n_445),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_628),
.B(n_445),
.Y(n_733)
);

OR2x6_ASAP7_75t_L g734 ( 
.A(n_567),
.B(n_450),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_519),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_562),
.B(n_501),
.C(n_455),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_610),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_646),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_522),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_638),
.B(n_450),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_555),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_522),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_636),
.A2(n_466),
.B1(n_499),
.B2(n_490),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_635),
.A2(n_466),
.B1(n_490),
.B2(n_478),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_616),
.B(n_501),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_646),
.B(n_450),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_529),
.B(n_450),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_604),
.A2(n_490),
.B1(n_478),
.B2(n_469),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_551),
.A2(n_478),
.B1(n_469),
.B2(n_466),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_529),
.B(n_455),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_630),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_523),
.B(n_215),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_523),
.B(n_337),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_529),
.B(n_455),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_514),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_560),
.B(n_456),
.C(n_455),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_529),
.B(n_456),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_642),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_529),
.B(n_456),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_511),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_590),
.B(n_456),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_531),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_634),
.B(n_459),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_634),
.A2(n_490),
.B1(n_478),
.B2(n_469),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_533),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_533),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_511),
.B(n_459),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_511),
.B(n_459),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_634),
.B(n_459),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_647),
.B(n_466),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_528),
.A2(n_279),
.B1(n_288),
.B2(n_335),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_634),
.A2(n_236),
.B1(n_189),
.B2(n_232),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_627),
.A2(n_236),
.B1(n_240),
.B2(n_256),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_557),
.B(n_232),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_506),
.B(n_261),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_634),
.B(n_433),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_506),
.B(n_269),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_634),
.B(n_433),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_506),
.B(n_433),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_627),
.B(n_256),
.C(n_240),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_621),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_592),
.Y(n_783)
);

BUFx5_ASAP7_75t_L g784 ( 
.A(n_513),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_509),
.B(n_524),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_509),
.B(n_433),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_509),
.B(n_433),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_524),
.B(n_433),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_641),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_528),
.A2(n_284),
.B1(n_294),
.B2(n_301),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_524),
.B(n_435),
.Y(n_791)
);

NOR2xp67_ASAP7_75t_L g792 ( 
.A(n_515),
.B(n_435),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_511),
.B(n_282),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_513),
.A2(n_242),
.B1(n_241),
.B2(n_239),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_532),
.B(n_435),
.Y(n_795)
);

AO22x2_ASAP7_75t_L g796 ( 
.A1(n_632),
.A2(n_322),
.B1(n_270),
.B2(n_274),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_532),
.B(n_435),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_532),
.B(n_435),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_546),
.B(n_283),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_514),
.B(n_337),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_538),
.A2(n_265),
.B1(n_310),
.B2(n_297),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_622),
.B(n_265),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_546),
.B(n_287),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_546),
.B(n_435),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_549),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_514),
.B(n_194),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_746),
.A2(n_517),
.B(n_516),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_656),
.A2(n_517),
.B(n_516),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_656),
.A2(n_527),
.B(n_526),
.Y(n_809)
);

NOR2x1_ASAP7_75t_L g810 ( 
.A(n_699),
.B(n_538),
.Y(n_810)
);

OAI21xp33_ASAP7_75t_L g811 ( 
.A1(n_684),
.A2(n_293),
.B(n_290),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_653),
.B(n_614),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_760),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_684),
.B(n_614),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_677),
.A2(n_527),
.B(n_526),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_693),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_722),
.B(n_614),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_760),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_710),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_703),
.B(n_623),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_785),
.A2(n_541),
.B(n_536),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_668),
.A2(n_541),
.B(n_536),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_726),
.B(n_514),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_670),
.A2(n_579),
.B(n_548),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_708),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_726),
.B(n_623),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_657),
.A2(n_579),
.B(n_548),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_709),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_738),
.A2(n_589),
.B(n_588),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_710),
.B(n_514),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_699),
.B(n_572),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_673),
.A2(n_589),
.B(n_588),
.Y(n_832)
);

AOI21xp33_ASAP7_75t_L g833 ( 
.A1(n_675),
.A2(n_539),
.B(n_632),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_728),
.B(n_572),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_685),
.A2(n_597),
.B(n_593),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_651),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_688),
.A2(n_597),
.B(n_593),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_771),
.A2(n_600),
.B(n_598),
.Y(n_838)
);

NOR2x1_ASAP7_75t_L g839 ( 
.A(n_741),
.B(n_585),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_730),
.B(n_573),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_730),
.B(n_573),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_700),
.B(n_582),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_701),
.B(n_582),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_692),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_675),
.A2(n_603),
.B(n_606),
.C(n_640),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_771),
.A2(n_600),
.B(n_598),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_677),
.A2(n_745),
.B(n_702),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_755),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_669),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_716),
.B(n_741),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_725),
.A2(n_530),
.B1(n_645),
.B2(n_648),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_716),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_725),
.A2(n_530),
.B1(n_645),
.B2(n_648),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_745),
.A2(n_607),
.B(n_605),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_719),
.B(n_724),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_662),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_710),
.B(n_544),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_733),
.A2(n_640),
.B(n_603),
.C(n_606),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_666),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_723),
.A2(n_607),
.B(n_605),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_732),
.B(n_612),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_696),
.B(n_612),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_663),
.A2(n_620),
.B(n_611),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_789),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_663),
.A2(n_620),
.B(n_611),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_717),
.B(n_539),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_664),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_674),
.A2(n_626),
.B1(n_625),
.B2(n_624),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_792),
.B(n_618),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_735),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_698),
.B(n_618),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_665),
.B(n_544),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_678),
.A2(n_679),
.B1(n_660),
.B2(n_667),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_682),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_689),
.B(n_625),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_782),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_690),
.B(n_624),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_695),
.B(n_626),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_720),
.B(n_544),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_739),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_706),
.A2(n_544),
.B1(n_329),
.B2(n_328),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_671),
.A2(n_637),
.B(n_585),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_671),
.A2(n_637),
.B(n_220),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_731),
.B(n_270),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_676),
.A2(n_429),
.B(n_434),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_761),
.B(n_274),
.Y(n_887)
);

AO21x1_ASAP7_75t_L g888 ( 
.A1(n_681),
.A2(n_434),
.B(n_429),
.Y(n_888)
);

AOI21xp33_ASAP7_75t_L g889 ( 
.A1(n_761),
.A2(n_721),
.B(n_756),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_737),
.B(n_297),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_672),
.A2(n_203),
.B(n_286),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_751),
.B(n_758),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_676),
.A2(n_429),
.B(n_434),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_762),
.A2(n_312),
.B(n_322),
.C(n_323),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_711),
.B(n_310),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_727),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_755),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_755),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_727),
.B(n_621),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_683),
.A2(n_323),
.B(n_312),
.C(n_331),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_742),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_718),
.A2(n_311),
.B1(n_313),
.B2(n_326),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_774),
.A2(n_331),
.B(n_430),
.C(n_320),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_672),
.A2(n_257),
.B(n_185),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_734),
.B(n_430),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_713),
.B(n_430),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_691),
.A2(n_680),
.B(n_705),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_707),
.A2(n_263),
.B(n_190),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_686),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_650),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_784),
.B(n_238),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_734),
.B(n_431),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_704),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_784),
.B(n_661),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_697),
.B(n_715),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_763),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_780),
.A2(n_264),
.B(n_191),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_784),
.B(n_238),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_729),
.B(n_334),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_659),
.B(n_334),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_712),
.B(n_334),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_786),
.A2(n_788),
.B(n_787),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_791),
.A2(n_272),
.B(n_333),
.Y(n_923)
);

NOR2x1_ASAP7_75t_R g924 ( 
.A(n_652),
.B(n_173),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_692),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_691),
.A2(n_714),
.B(n_766),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_783),
.B(n_431),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_795),
.A2(n_255),
.B(n_330),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_767),
.A2(n_254),
.B(n_325),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_784),
.B(n_661),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_797),
.A2(n_250),
.B(n_324),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_798),
.A2(n_248),
.B(n_319),
.Y(n_932)
);

AO21x1_ASAP7_75t_L g933 ( 
.A1(n_740),
.A2(n_431),
.B(n_316),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_784),
.B(n_199),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_781),
.B(n_208),
.C(n_213),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_804),
.A2(n_276),
.B(n_222),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_734),
.A2(n_278),
.B1(n_225),
.B2(n_315),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_800),
.A2(n_431),
.B(n_316),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_658),
.B(n_8),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_772),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_773),
.B(n_228),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_782),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_796),
.B(n_431),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_790),
.A2(n_694),
.B(n_776),
.C(n_799),
.Y(n_944)
);

AOI21xp33_ASAP7_75t_L g945 ( 
.A1(n_736),
.A2(n_291),
.B(n_235),
.Y(n_945)
);

O2A1O1Ixp5_ASAP7_75t_L g946 ( 
.A1(n_800),
.A2(n_431),
.B(n_19),
.C(n_21),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_782),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_805),
.A2(n_295),
.B(n_243),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_749),
.B(n_18),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_770),
.A2(n_298),
.B(n_273),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_776),
.A2(n_302),
.B(n_306),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_796),
.B(n_431),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_773),
.B(n_308),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_743),
.B(n_27),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_752),
.A2(n_431),
.B(n_316),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_764),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_687),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_778),
.A2(n_316),
.B(n_280),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_796),
.B(n_431),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_778),
.A2(n_316),
.B(n_280),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_799),
.A2(n_234),
.B(n_233),
.C(n_194),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_803),
.A2(n_280),
.B(n_234),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_775),
.B(n_28),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_752),
.B(n_280),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_803),
.B(n_29),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_747),
.A2(n_280),
.B(n_234),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_775),
.B(n_30),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_768),
.B(n_30),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_768),
.B(n_32),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_769),
.B(n_34),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_743),
.A2(n_36),
.B(n_41),
.C(n_42),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_747),
.A2(n_234),
.B(n_233),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_753),
.B(n_36),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_753),
.B(n_744),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_744),
.B(n_42),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_802),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_765),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_748),
.B(n_45),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_777),
.B(n_101),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_655),
.A2(n_748),
.B(n_779),
.C(n_801),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_801),
.A2(n_233),
.B1(n_194),
.B2(n_50),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_913),
.B(n_794),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_913),
.B(n_802),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_816),
.B(n_769),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_965),
.A2(n_655),
.B(n_759),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_865),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_814),
.A2(n_793),
.B(n_806),
.Y(n_987)
);

INVxp33_ASAP7_75t_L g988 ( 
.A(n_867),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_965),
.A2(n_759),
.B(n_757),
.C(n_754),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_944),
.A2(n_806),
.B(n_757),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_820),
.A2(n_654),
.B(n_754),
.C(n_750),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_856),
.B(n_46),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_957),
.B(n_46),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_850),
.B(n_47),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_971),
.A2(n_52),
.B(n_53),
.C(n_57),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_874),
.A2(n_233),
.B1(n_194),
.B2(n_59),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_833),
.B(n_53),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_916),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_819),
.B(n_194),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_852),
.B(n_854),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_836),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_853),
.B(n_60),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_868),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_877),
.Y(n_1004)
);

BUFx8_ASAP7_75t_L g1005 ( 
.A(n_925),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_947),
.B(n_118),
.Y(n_1006)
);

BUFx12f_ASAP7_75t_L g1007 ( 
.A(n_877),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_845),
.B(n_127),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_949),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_R g1010 ( 
.A(n_963),
.B(n_976),
.Y(n_1010)
);

OA22x2_ASAP7_75t_L g1011 ( 
.A1(n_896),
.A2(n_63),
.B1(n_161),
.B2(n_74),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_853),
.B(n_69),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_892),
.B(n_79),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_899),
.Y(n_1014)
);

AND2x6_ASAP7_75t_SL g1015 ( 
.A(n_967),
.B(n_84),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_813),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_817),
.A2(n_87),
.B1(n_91),
.B2(n_102),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_831),
.Y(n_1018)
);

NAND2x1p5_ASAP7_75t_L g1019 ( 
.A(n_813),
.B(n_108),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_820),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_826),
.A2(n_150),
.B1(n_154),
.B2(n_157),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_875),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_819),
.B(n_813),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_811),
.A2(n_940),
.B(n_935),
.C(n_894),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_857),
.A2(n_860),
.B1(n_981),
.B2(n_834),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_851),
.B(n_813),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_934),
.A2(n_848),
.B(n_922),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_825),
.Y(n_1028)
);

AOI22x1_ASAP7_75t_L g1029 ( 
.A1(n_835),
.A2(n_824),
.B1(n_822),
.B2(n_832),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_926),
.A2(n_812),
.B(n_914),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_915),
.B(n_910),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_828),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_914),
.A2(n_930),
.B(n_807),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_967),
.B(n_943),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_819),
.B(n_818),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_844),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_819),
.B(n_935),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_930),
.A2(n_907),
.B(n_838),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_981),
.A2(n_974),
.B1(n_949),
.B2(n_879),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_952),
.B(n_959),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_847),
.A2(n_872),
.B(n_863),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_937),
.B(n_844),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_954),
.A2(n_980),
.B1(n_880),
.B2(n_977),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_885),
.B(n_890),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_910),
.B(n_924),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_844),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_887),
.B(n_895),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_973),
.A2(n_968),
.B1(n_969),
.B2(n_970),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_878),
.A2(n_862),
.B(n_843),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_844),
.B(n_849),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_900),
.A2(n_909),
.B(n_889),
.C(n_978),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_905),
.B(n_912),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_876),
.A2(n_975),
.B1(n_812),
.B2(n_842),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_840),
.B(n_841),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_827),
.A2(n_861),
.B(n_837),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_902),
.B(n_956),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_870),
.A2(n_871),
.B1(n_901),
.B2(n_881),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_927),
.B(n_939),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_849),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_968),
.A2(n_970),
.B1(n_969),
.B2(n_939),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_870),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_911),
.A2(n_918),
.B(n_960),
.C(n_958),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_849),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_903),
.A2(n_882),
.B(n_929),
.C(n_846),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_876),
.A2(n_955),
.B(n_883),
.C(n_808),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_821),
.A2(n_809),
.B(n_864),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_941),
.A2(n_953),
.B1(n_956),
.B2(n_964),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_859),
.A2(n_918),
.B(n_911),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_912),
.B(n_898),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_921),
.B(n_919),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_897),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_810),
.B(n_898),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_869),
.A2(n_946),
.B(n_823),
.C(n_951),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_R g1075 ( 
.A(n_897),
.B(n_898),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_906),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_873),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_SL g1078 ( 
.A1(n_815),
.A2(n_830),
.B(n_839),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_830),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_920),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_886),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_979),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_SL g1083 ( 
.A(n_979),
.B(n_858),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_893),
.B(n_950),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_948),
.B(n_904),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_946),
.A2(n_945),
.B1(n_891),
.B2(n_884),
.C(n_961),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_873),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_859),
.A2(n_855),
.B(n_829),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_962),
.A2(n_908),
.B(n_932),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_917),
.B(n_936),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_923),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_866),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_931),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_966),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_972),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_933),
.A2(n_866),
.B(n_859),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_938),
.B(n_850),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_967),
.A2(n_632),
.B1(n_500),
.B2(n_347),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_856),
.A2(n_684),
.B1(n_657),
.B2(n_965),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_850),
.B(n_507),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_942),
.B(n_652),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_913),
.B(n_354),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_SL g1104 ( 
.A1(n_965),
.A2(n_684),
.B(n_771),
.C(n_559),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_836),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_850),
.B(n_467),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_856),
.B(n_728),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_865),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_818),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_965),
.A2(n_507),
.B(n_684),
.C(n_675),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_850),
.B(n_507),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_965),
.A2(n_684),
.B(n_771),
.C(n_559),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_856),
.B(n_728),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_856),
.A2(n_684),
.B1(n_657),
.B2(n_965),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_816),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_814),
.A2(n_684),
.B(n_944),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_965),
.A2(n_703),
.B(n_684),
.C(n_653),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1061),
.C(n_1099),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1119),
.A2(n_1106),
.B(n_1102),
.Y(n_1126)
);

AO32x2_ASAP7_75t_L g1127 ( 
.A1(n_1049),
.A2(n_1044),
.A3(n_1054),
.B1(n_1040),
.B2(n_996),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1124),
.A2(n_1106),
.B(n_1102),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1024),
.A2(n_1000),
.B(n_1052),
.C(n_982),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1001),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1048),
.B(n_1108),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_986),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1113),
.A2(n_1117),
.B(n_1115),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_1101),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_997),
.A2(n_995),
.B1(n_1116),
.B2(n_1103),
.C(n_1098),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1113),
.A2(n_1117),
.B(n_1115),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_1109),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1004),
.B(n_1006),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1104),
.A2(n_1114),
.B(n_1009),
.C(n_992),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1081),
.A2(n_1122),
.B1(n_1121),
.B2(n_1118),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1120),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1055),
.B(n_1118),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1046),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1014),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1052),
.A2(n_1065),
.B(n_985),
.C(n_1045),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1034),
.B(n_988),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_1070),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1121),
.A2(n_1123),
.B1(n_1122),
.B2(n_993),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1123),
.A2(n_1042),
.B(n_1084),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1107),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_SL g1152 ( 
.A1(n_1095),
.A2(n_1085),
.B(n_1092),
.C(n_1043),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1042),
.A2(n_1050),
.B(n_1066),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1039),
.A2(n_1033),
.B(n_990),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1067),
.A2(n_1069),
.B(n_1088),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1059),
.B(n_1076),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1067),
.A2(n_1069),
.B(n_1090),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1075),
.B(n_1082),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1105),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1093),
.A2(n_990),
.B(n_1089),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_995),
.A2(n_1057),
.B(n_1074),
.C(n_989),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1025),
.B(n_1031),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1063),
.A2(n_987),
.B(n_1094),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1060),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_983),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1100),
.A2(n_1112),
.B1(n_984),
.B2(n_1011),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_994),
.B(n_1036),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1013),
.A2(n_1083),
.B(n_1086),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_991),
.A2(n_1002),
.B(n_1038),
.C(n_1078),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_1091),
.B(n_1068),
.C(n_1017),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_989),
.A2(n_1020),
.B(n_1051),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1080),
.A2(n_1079),
.B(n_1097),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1015),
.B(n_1053),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1005),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1053),
.B(n_1022),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1005),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1019),
.A2(n_1012),
.B(n_999),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_1008),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1021),
.A2(n_1087),
.B(n_1047),
.C(n_1035),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1023),
.A2(n_1072),
.B(n_1073),
.Y(n_1182)
);

OAI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1018),
.A2(n_1026),
.B1(n_1073),
.B2(n_1032),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1028),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1071),
.A2(n_1058),
.B(n_1026),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1041),
.B(n_1062),
.Y(n_1186)
);

AO32x2_ASAP7_75t_L g1187 ( 
.A1(n_1047),
.A2(n_1087),
.A3(n_1041),
.B1(n_1016),
.B2(n_1072),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1072),
.B(n_1077),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_SL g1189 ( 
.A(n_1037),
.Y(n_1189)
);

BUFx4_ASAP7_75t_R g1190 ( 
.A(n_1037),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_SL g1191 ( 
.A1(n_1110),
.A2(n_1111),
.B(n_1124),
.C(n_1119),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1064),
.A2(n_1111),
.B(n_1099),
.Y(n_1192)
);

AOI221x1_ASAP7_75t_L g1193 ( 
.A1(n_1064),
.A2(n_1111),
.B1(n_1049),
.B2(n_1119),
.C(n_1099),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1109),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1001),
.Y(n_1197)
);

INVx8_ASAP7_75t_L g1198 ( 
.A(n_1007),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1096),
.A2(n_1027),
.B(n_1056),
.Y(n_1199)
);

AOI221x1_ASAP7_75t_L g1200 ( 
.A1(n_1111),
.A2(n_1049),
.B1(n_1119),
.B2(n_1099),
.C(n_965),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1030),
.A2(n_933),
.A3(n_888),
.B(n_1033),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1099),
.C(n_1119),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1119),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1111),
.A2(n_1119),
.B(n_1099),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1001),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1069),
.A2(n_933),
.B(n_1056),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1001),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1103),
.B(n_500),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1061),
.C(n_1119),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1111),
.B(n_1061),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1016),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1109),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1049),
.A2(n_507),
.B1(n_432),
.B2(n_627),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1034),
.B(n_867),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1109),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1219)
);

AOI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_1111),
.A2(n_997),
.B1(n_1119),
.B2(n_1099),
.C(n_774),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1111),
.A2(n_1119),
.B(n_1099),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1111),
.B(n_1061),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1103),
.B(n_500),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1049),
.A2(n_507),
.B1(n_432),
.B2(n_627),
.Y(n_1227)
);

AOI221x1_ASAP7_75t_L g1228 ( 
.A1(n_1111),
.A2(n_1049),
.B1(n_1119),
.B2(n_1099),
.C(n_965),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1103),
.B(n_500),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1061),
.C(n_1119),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_986),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1107),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1109),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1030),
.A2(n_933),
.A3(n_888),
.B(n_1033),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1053),
.B(n_853),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1069),
.A2(n_933),
.B(n_1056),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_986),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1030),
.A2(n_933),
.A3(n_888),
.B(n_1033),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1030),
.A2(n_933),
.A3(n_888),
.B(n_1033),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1003),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1049),
.A2(n_507),
.B1(n_432),
.B2(n_627),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1111),
.A2(n_1119),
.B(n_1099),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1061),
.C(n_1119),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1003),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1016),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1248)
);

AOI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1102),
.A2(n_1113),
.B(n_1106),
.Y(n_1249)
);

AOI221xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1111),
.A2(n_995),
.B1(n_1124),
.B2(n_1024),
.C(n_811),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1061),
.C(n_1119),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1005),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1056),
.A2(n_1029),
.B(n_1027),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1030),
.A2(n_933),
.A3(n_888),
.B(n_1033),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1102),
.A2(n_1113),
.B(n_1106),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_986),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1119),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1111),
.B(n_500),
.C(n_440),
.Y(n_1259)
);

AOI221x1_ASAP7_75t_L g1260 ( 
.A1(n_1111),
.A2(n_1049),
.B1(n_1119),
.B2(n_1099),
.C(n_965),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1261)
);

AO32x2_ASAP7_75t_L g1262 ( 
.A1(n_1049),
.A2(n_1044),
.A3(n_1054),
.B1(n_1040),
.B2(n_996),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_SL g1263 ( 
.A1(n_1194),
.A2(n_1248),
.B1(n_1261),
.B2(n_1206),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1136),
.A2(n_1220),
.B1(n_1212),
.B2(n_1223),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1190),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1135),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1166),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1159),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1194),
.A2(n_1222),
.B1(n_1261),
.B2(n_1225),
.Y(n_1269)
);

BUFx8_ASAP7_75t_L g1270 ( 
.A(n_1175),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1197),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1145),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1207),
.Y(n_1273)
);

BUFx8_ASAP7_75t_L g1274 ( 
.A(n_1133),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1136),
.A2(n_1220),
.B1(n_1227),
.B2(n_1215),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1257),
.Y(n_1276)
);

INVx4_ASAP7_75t_SL g1277 ( 
.A(n_1189),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1138),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1242),
.A2(n_1203),
.B1(n_1252),
.B2(n_1225),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1231),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1209),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1198),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1198),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1222),
.A2(n_1205),
.B1(n_1217),
.B2(n_1204),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1145),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1238),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1200),
.A2(n_1260),
.B1(n_1228),
.B2(n_1193),
.Y(n_1287)
);

BUFx10_ASAP7_75t_L g1288 ( 
.A(n_1210),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_L g1289 ( 
.A1(n_1125),
.A2(n_1245),
.B(n_1230),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1205),
.A2(n_1258),
.B1(n_1204),
.B2(n_1171),
.Y(n_1290)
);

INVx8_ASAP7_75t_L g1291 ( 
.A(n_1198),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1221),
.A2(n_1243),
.B1(n_1258),
.B2(n_1167),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1144),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1211),
.A2(n_1251),
.B(n_1229),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1162),
.A2(n_1131),
.B1(n_1156),
.B2(n_1163),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1176),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1144),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1224),
.A2(n_1259),
.B(n_1161),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1174),
.A2(n_1162),
.B1(n_1131),
.B2(n_1180),
.Y(n_1299)
);

INVx3_ASAP7_75t_SL g1300 ( 
.A(n_1234),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1146),
.A2(n_1192),
.B1(n_1126),
.B2(n_1128),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1128),
.A2(n_1141),
.B1(n_1149),
.B2(n_1143),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_1156),
.B1(n_1246),
.B2(n_1241),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1213),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1202),
.A2(n_1169),
.B(n_1134),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1166),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1178),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1234),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1151),
.A2(n_1232),
.B1(n_1149),
.B2(n_1168),
.Y(n_1309)
);

BUFx2_ASAP7_75t_SL g1310 ( 
.A(n_1196),
.Y(n_1310)
);

BUFx2_ASAP7_75t_SL g1311 ( 
.A(n_1214),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1218),
.B(n_1148),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1213),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

OAI21xp33_ASAP7_75t_L g1315 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1141),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1184),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1187),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1142),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1148),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1143),
.A2(n_1137),
.B1(n_1169),
.B2(n_1154),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1250),
.A2(n_1191),
.B(n_1170),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1139),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1154),
.A2(n_1155),
.B1(n_1153),
.B2(n_1256),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1186),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1187),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1247),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1127),
.A2(n_1262),
.B1(n_1188),
.B2(n_1183),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1185),
.A2(n_1127),
.B1(n_1262),
.B2(n_1158),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1249),
.A2(n_1150),
.B1(n_1157),
.B2(n_1160),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1182),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1173),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1140),
.Y(n_1332)
);

BUFx2_ASAP7_75t_SL g1333 ( 
.A(n_1172),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1173),
.A2(n_1150),
.B1(n_1237),
.B2(n_1208),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1208),
.A2(n_1237),
.B1(n_1179),
.B2(n_1199),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1164),
.A2(n_1132),
.B1(n_1254),
.B2(n_1244),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1195),
.A2(n_1219),
.B1(n_1233),
.B2(n_1226),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1201),
.B(n_1235),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1181),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1216),
.A2(n_1201),
.B1(n_1235),
.B2(n_1239),
.Y(n_1340)
);

OAI21xp33_ASAP7_75t_L g1341 ( 
.A1(n_1152),
.A2(n_1235),
.B(n_1239),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1255),
.A2(n_1111),
.B1(n_1203),
.B2(n_1194),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1255),
.A2(n_1000),
.B1(n_796),
.B2(n_1136),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1255),
.A2(n_1000),
.B1(n_796),
.B2(n_1136),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1138),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1194),
.A2(n_1000),
.B1(n_796),
.B2(n_1049),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1145),
.Y(n_1348)
);

CKINVDCx6p67_ASAP7_75t_R g1349 ( 
.A(n_1253),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1194),
.B(n_1061),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1130),
.Y(n_1351)
);

CKINVDCx6p67_ASAP7_75t_R g1352 ( 
.A(n_1253),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1166),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1131),
.B(n_1129),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1190),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1215),
.A2(n_1242),
.B1(n_1227),
.B2(n_1228),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1177),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1198),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1215),
.A2(n_1242),
.B1(n_1227),
.B2(n_1228),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1215),
.A2(n_1242),
.B1(n_1227),
.B2(n_1228),
.Y(n_1360)
);

AND2x4_ASAP7_75t_SL g1361 ( 
.A(n_1144),
.B(n_1236),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1136),
.A2(n_1000),
.B1(n_796),
.B2(n_833),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1130),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1136),
.A2(n_1000),
.B1(n_796),
.B2(n_833),
.Y(n_1364)
);

INVxp33_ASAP7_75t_L g1365 ( 
.A(n_1280),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1320),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1315),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1323),
.A2(n_1337),
.B(n_1305),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1318),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1362),
.A2(n_1364),
.B1(n_1347),
.B2(n_1345),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1338),
.B(n_1268),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1271),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1273),
.B(n_1281),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1276),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1341),
.A2(n_1337),
.B(n_1334),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1278),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1351),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1317),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1363),
.B(n_1328),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1342),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1301),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1328),
.B(n_1263),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1362),
.A2(n_1364),
.B1(n_1347),
.B2(n_1344),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1343),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1339),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1339),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1317),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1310),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1267),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1317),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1325),
.B(n_1265),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1357),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1325),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1327),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1350),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1265),
.B(n_1355),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1334),
.A2(n_1335),
.B(n_1336),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1319),
.Y(n_1400)
);

INVx11_ASAP7_75t_L g1401 ( 
.A(n_1270),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1335),
.A2(n_1321),
.B(n_1290),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1331),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1339),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1350),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1263),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1294),
.A2(n_1264),
.B(n_1290),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1269),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1269),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1332),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1311),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1279),
.B(n_1284),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1354),
.B(n_1279),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1329),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1329),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1284),
.A2(n_1289),
.B(n_1264),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1340),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1340),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1275),
.A2(n_1309),
.B(n_1303),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1292),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1326),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1344),
.A2(n_1345),
.B1(n_1355),
.B2(n_1275),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1300),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1306),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1309),
.B(n_1296),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1295),
.B(n_1287),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1307),
.A2(n_1316),
.B(n_1333),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1295),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1353),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1298),
.A2(n_1287),
.B(n_1326),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1300),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1356),
.A2(n_1360),
.B(n_1359),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1296),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1330),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1356),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1308),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1414),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1407),
.A2(n_1360),
.B1(n_1359),
.B2(n_1299),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1407),
.A2(n_1299),
.B1(n_1322),
.B2(n_1353),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1368),
.B(n_1288),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1370),
.B(n_1286),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1393),
.B(n_1285),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1368),
.B(n_1288),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1432),
.A2(n_1348),
.B1(n_1272),
.B2(n_1285),
.C(n_1297),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1378),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1367),
.B(n_1313),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1432),
.A2(n_1272),
.B(n_1358),
.C(n_1322),
.Y(n_1447)
);

AO21x1_ASAP7_75t_L g1448 ( 
.A1(n_1426),
.A2(n_1361),
.B(n_1304),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1426),
.A2(n_1314),
.B(n_1324),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1423),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1410),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1367),
.B(n_1366),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1394),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1366),
.B(n_1274),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1434),
.B(n_1431),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1434),
.B(n_1283),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1376),
.B(n_1283),
.Y(n_1457)
);

AO32x1_ASAP7_75t_L g1458 ( 
.A1(n_1387),
.A2(n_1282),
.A3(n_1274),
.B1(n_1293),
.B2(n_1346),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1375),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1375),
.B(n_1349),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1369),
.A2(n_1277),
.B(n_1291),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1369),
.A2(n_1277),
.B(n_1291),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1374),
.B(n_1352),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1383),
.A2(n_1415),
.B(n_1414),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.B(n_1266),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1412),
.A2(n_1413),
.B(n_1398),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1397),
.B(n_1405),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1405),
.B(n_1413),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_SL g1469 ( 
.A1(n_1410),
.A2(n_1436),
.B(n_1390),
.C(n_1401),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1391),
.A2(n_1400),
.A3(n_1372),
.B1(n_1396),
.B2(n_1381),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1393),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1365),
.B(n_1372),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_L g1473 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1433),
.B(n_1404),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1386),
.B(n_1420),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1412),
.A2(n_1385),
.B1(n_1371),
.B2(n_1406),
.C(n_1408),
.Y(n_1476)
);

AO32x2_ASAP7_75t_L g1477 ( 
.A1(n_1391),
.A2(n_1381),
.A3(n_1417),
.B1(n_1418),
.B2(n_1380),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1416),
.A2(n_1402),
.B(n_1430),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1380),
.B(n_1388),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1416),
.A2(n_1402),
.B(n_1430),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1427),
.A2(n_1415),
.B(n_1428),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1419),
.A2(n_1408),
.B(n_1406),
.C(n_1409),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1422),
.A2(n_1409),
.B1(n_1420),
.B2(n_1435),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1389),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1410),
.B(n_1401),
.Y(n_1485)
);

AOI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1424),
.A2(n_1429),
.B(n_1428),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1461),
.B(n_1421),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1399),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1481),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1468),
.B(n_1386),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1468),
.B(n_1392),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1439),
.A2(n_1384),
.B1(n_1419),
.B2(n_1377),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1398),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1438),
.A2(n_1377),
.B1(n_1403),
.B2(n_1399),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1470),
.B(n_1399),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1470),
.B(n_1399),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1464),
.B(n_1382),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1472),
.B(n_1377),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1467),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1459),
.B(n_1377),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1450),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1437),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1437),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1464),
.B(n_1382),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1395),
.Y(n_1506)
);

AND2x6_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1421),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1475),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1452),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1484),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1440),
.B(n_1373),
.C(n_1379),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1442),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1493),
.B(n_1444),
.C(n_1440),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1493),
.A2(n_1483),
.B1(n_1476),
.B2(n_1449),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1488),
.A2(n_1483),
.B1(n_1476),
.B2(n_1482),
.C(n_1444),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1511),
.B(n_1443),
.C(n_1480),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1511),
.B(n_1443),
.C(n_1480),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1503),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1501),
.B(n_1455),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1502),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1502),
.B(n_1454),
.C(n_1446),
.D(n_1469),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1489),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1503),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1501),
.B(n_1465),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1504),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1492),
.B(n_1462),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1453),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1507),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1491),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_SL g1533 ( 
.A(n_1507),
.B(n_1447),
.Y(n_1533)
);

AO21x2_ASAP7_75t_L g1534 ( 
.A1(n_1489),
.A2(n_1478),
.B(n_1486),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1501),
.B(n_1499),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_1466),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1507),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1488),
.B(n_1478),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_SL g1539 ( 
.A(n_1496),
.B(n_1447),
.C(n_1448),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1441),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1512),
.B(n_1471),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1495),
.A2(n_1505),
.B(n_1498),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1512),
.B(n_1474),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1535),
.B(n_1496),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1529),
.B(n_1508),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1535),
.B(n_1525),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1518),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1524),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1525),
.B(n_1496),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1523),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1516),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1531),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1534),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1524),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1531),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1532),
.B(n_1490),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1497),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1537),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1526),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1539),
.B(n_1517),
.C(n_1516),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1534),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1537),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1520),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1521),
.B(n_1508),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1538),
.B(n_1506),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.B(n_1506),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1487),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1542),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1553),
.A2(n_1514),
.B1(n_1515),
.B2(n_1536),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1548),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1574),
.B(n_1542),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1544),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1548),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1574),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1558),
.B(n_1532),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1549),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1556),
.B(n_1567),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1567),
.B(n_1513),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1546),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1547),
.B(n_1544),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1571),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1547),
.B(n_1543),
.Y(n_1596)
);

NAND2x1_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1536),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1550),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1550),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1552),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1543),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1550),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1513),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1558),
.B(n_1521),
.Y(n_1607)
);

OAI31xp67_ASAP7_75t_L g1608 ( 
.A1(n_1546),
.A2(n_1510),
.A3(n_1573),
.B(n_1572),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1560),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1560),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1571),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1551),
.B(n_1541),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1565),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1560),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1578),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1579),
.B(n_1571),
.Y(n_1622)
);

NAND2x1_ASAP7_75t_L g1623 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1579),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1625)
);

NOR2x2_ASAP7_75t_L g1626 ( 
.A(n_1608),
.B(n_1575),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1551),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1578),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1591),
.A2(n_1539),
.B(n_1515),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1545),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1583),
.B(n_1546),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1584),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1596),
.B(n_1545),
.Y(n_1633)
);

NAND2xp67_ASAP7_75t_L g1634 ( 
.A(n_1576),
.B(n_1572),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1590),
.B(n_1606),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1582),
.B(n_1556),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1577),
.A2(n_1590),
.B1(n_1585),
.B2(n_1536),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1596),
.B(n_1545),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1613),
.B(n_1566),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1588),
.B(n_1563),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1545),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1603),
.B(n_1563),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1563),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1584),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1597),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1613),
.B(n_1566),
.Y(n_1646)
);

XOR2x2_ASAP7_75t_L g1647 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1589),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1563),
.Y(n_1649)
);

AOI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1612),
.A2(n_1569),
.A3(n_1564),
.B(n_1485),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1587),
.B(n_1556),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1554),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1586),
.Y(n_1654)
);

INVx3_ASAP7_75t_SL g1655 ( 
.A(n_1586),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1635),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1655),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1636),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_SL g1660 ( 
.A1(n_1634),
.A2(n_1608),
.B(n_1617),
.C(n_1614),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1629),
.A2(n_1538),
.B1(n_1449),
.B2(n_1573),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1615),
.Y(n_1663)
);

OAI322xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1652),
.A2(n_1607),
.A3(n_1611),
.B1(n_1605),
.B2(n_1589),
.C1(n_1581),
.C2(n_1610),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

AOI31xp33_ASAP7_75t_L g1666 ( 
.A1(n_1654),
.A2(n_1595),
.A3(n_1564),
.B(n_1569),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1624),
.A2(n_1573),
.B(n_1572),
.C(n_1568),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1625),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1643),
.B(n_1554),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1650),
.A2(n_1569),
.B(n_1564),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1624),
.B(n_1605),
.C(n_1598),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1554),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1625),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1643),
.B(n_1555),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1623),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1640),
.B(n_1555),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1622),
.B(n_1599),
.C(n_1593),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1630),
.B(n_1633),
.Y(n_1679)
);

OAI322xp33_ASAP7_75t_L g1680 ( 
.A1(n_1622),
.A2(n_1616),
.A3(n_1559),
.B1(n_1568),
.B2(n_1618),
.C1(n_1609),
.C2(n_1600),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1657),
.B(n_1637),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1656),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1663),
.B(n_1630),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1668),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1665),
.A2(n_1538),
.B1(n_1647),
.B2(n_1559),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1633),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1663),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1679),
.B(n_1638),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1660),
.A2(n_1631),
.B(n_1623),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1679),
.B(n_1638),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1676),
.Y(n_1692)
);

OAI21xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1666),
.A2(n_1651),
.B(n_1631),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1676),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1658),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1665),
.A2(n_1538),
.B1(n_1647),
.B2(n_1568),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1662),
.A2(n_1651),
.B1(n_1559),
.B2(n_1538),
.C(n_1645),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1675),
.A2(n_1573),
.B1(n_1651),
.B2(n_1536),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1675),
.A2(n_1651),
.B1(n_1536),
.B2(n_1533),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1662),
.A2(n_1533),
.B1(n_1534),
.B2(n_1495),
.Y(n_1702)
);

XOR2xp5_ASAP7_75t_L g1703 ( 
.A(n_1688),
.B(n_1671),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_L g1704 ( 
.A(n_1683),
.B(n_1680),
.C(n_1671),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1687),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1689),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1684),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1685),
.Y(n_1708)
);

XNOR2xp5_ASAP7_75t_L g1709 ( 
.A(n_1686),
.B(n_1659),
.Y(n_1709)
);

AOI31xp33_ASAP7_75t_L g1710 ( 
.A1(n_1685),
.A2(n_1670),
.A3(n_1678),
.B(n_1681),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1694),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1702),
.A2(n_1698),
.B1(n_1682),
.B2(n_1693),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1707),
.Y(n_1714)
);

NAND2x1_ASAP7_75t_L g1715 ( 
.A(n_1710),
.B(n_1690),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1683),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1708),
.Y(n_1717)
);

NAND4xp25_ASAP7_75t_L g1718 ( 
.A(n_1704),
.B(n_1692),
.C(n_1695),
.D(n_1670),
.Y(n_1718)
);

AOI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1703),
.A2(n_1697),
.B(n_1696),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1704),
.B(n_1667),
.C(n_1699),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1705),
.B(n_1680),
.C(n_1661),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1712),
.C(n_1711),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1720),
.A2(n_1709),
.B1(n_1700),
.B2(n_1701),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1715),
.A2(n_1672),
.B1(n_1645),
.B2(n_1706),
.C(n_1681),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1721),
.A2(n_1664),
.B(n_1645),
.C(n_1646),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1716),
.Y(n_1726)
);

NAND4xp75_ASAP7_75t_L g1727 ( 
.A(n_1719),
.B(n_1669),
.C(n_1674),
.D(n_1649),
.Y(n_1727)
);

NAND4xp25_ASAP7_75t_L g1728 ( 
.A(n_1726),
.B(n_1722),
.C(n_1718),
.D(n_1714),
.Y(n_1728)
);

OAI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1725),
.A2(n_1717),
.B1(n_1639),
.B2(n_1646),
.C(n_1644),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1724),
.A2(n_1677),
.B(n_1639),
.C(n_1648),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_R g1731 ( 
.A(n_1727),
.B(n_1457),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1723),
.A2(n_1619),
.B1(n_1632),
.B2(n_1556),
.C(n_1674),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1726),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1733),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1669),
.Y(n_1735)
);

INVxp33_ASAP7_75t_SL g1736 ( 
.A(n_1731),
.Y(n_1736)
);

XOR2xp5_ASAP7_75t_L g1737 ( 
.A(n_1732),
.B(n_1463),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1729),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1738),
.C(n_1735),
.Y(n_1739)
);

NOR2x1p5_ASAP7_75t_L g1740 ( 
.A(n_1736),
.B(n_1730),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1737),
.B(n_1601),
.C(n_1587),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1740),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1742),
.Y(n_1743)
);

AND3x1_ASAP7_75t_L g1744 ( 
.A(n_1743),
.B(n_1739),
.C(n_1741),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1743),
.A2(n_1616),
.B1(n_1642),
.B2(n_1627),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1744),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1621),
.B1(n_1642),
.B2(n_1627),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1621),
.B1(n_1620),
.B2(n_1641),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1747),
.B(n_1601),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1602),
.B(n_1620),
.Y(n_1750)
);

OAI21xp33_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1748),
.B(n_1641),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1602),
.B1(n_1653),
.B2(n_1564),
.C(n_1569),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_R g1753 ( 
.A1(n_1752),
.A2(n_1653),
.B1(n_1458),
.B2(n_1561),
.C(n_1557),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1454),
.B(n_1460),
.C(n_1456),
.Y(n_1754)
);


endmodule