module real_aes_7917_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_792;
wire n_673;
wire n_503;
wire n_386;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_0), .A2(n_209), .B1(n_451), .B2(n_475), .Y(n_474) );
XOR2x2_ASAP7_75t_L g593 ( .A(n_1), .B(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_2), .A2(n_230), .B1(n_381), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_3), .A2(n_63), .B1(n_329), .B2(n_597), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_4), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_5), .A2(n_24), .B1(n_220), .B2(n_589), .C1(n_613), .C2(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_6), .A2(n_236), .B1(n_401), .B2(n_583), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_7), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_8), .A2(n_175), .B1(n_468), .B2(n_539), .Y(n_701) );
INVx1_ASAP7_75t_L g647 ( .A(n_9), .Y(n_647) );
OA22x2_ASAP7_75t_L g618 ( .A1(n_10), .A2(n_619), .B1(n_620), .B2(n_648), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_10), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_11), .A2(n_150), .B1(n_633), .B2(n_635), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_12), .A2(n_105), .B1(n_339), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_13), .A2(n_74), .B1(n_603), .B2(n_605), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_14), .A2(n_17), .B1(n_287), .B2(n_446), .C(n_448), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_15), .A2(n_64), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_16), .A2(n_223), .B1(n_675), .B2(n_676), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_18), .A2(n_266), .B1(n_338), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_19), .A2(n_76), .B1(n_287), .B2(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g769 ( .A(n_20), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_21), .A2(n_121), .B1(n_625), .B2(n_838), .Y(n_837) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_22), .A2(n_84), .B1(n_292), .B2(n_297), .Y(n_300) );
INVx1_ASAP7_75t_L g790 ( .A(n_22), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_23), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g588 ( .A1(n_25), .A2(n_103), .B1(n_126), .B2(n_421), .C1(n_513), .C2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_26), .A2(n_30), .B1(n_610), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_27), .A2(n_153), .B1(n_310), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_28), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_29), .A2(n_231), .B1(n_472), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g393 ( .A(n_31), .Y(n_393) );
AOI222xp33_ASAP7_75t_L g752 ( .A1(n_32), .A2(n_91), .B1(n_247), .B2(n_363), .C1(n_383), .C2(n_418), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_33), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_34), .A2(n_187), .B1(n_363), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_35), .A2(n_65), .B1(n_338), .B2(n_664), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_36), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_37), .A2(n_38), .B1(n_597), .B2(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g645 ( .A(n_39), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_40), .A2(n_208), .B1(n_355), .B2(n_539), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_41), .A2(n_159), .B1(n_346), .B2(n_559), .Y(n_575) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_42), .A2(n_87), .B1(n_292), .B2(n_293), .Y(n_302) );
INVx1_ASAP7_75t_L g791 ( .A(n_42), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_43), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_44), .A2(n_54), .B1(n_536), .B2(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_45), .A2(n_794), .B1(n_795), .B2(n_813), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_45), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_46), .A2(n_154), .B1(n_358), .B2(n_497), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_47), .A2(n_156), .B1(n_675), .B2(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_48), .Y(n_847) );
INVx1_ASAP7_75t_L g639 ( .A(n_49), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_50), .A2(n_268), .B1(n_303), .B2(n_437), .C(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g630 ( .A(n_51), .Y(n_630) );
INVx1_ASAP7_75t_L g638 ( .A(n_52), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_53), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_55), .A2(n_145), .B1(n_451), .B2(n_669), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_56), .B(n_597), .Y(n_692) );
INVx1_ASAP7_75t_L g567 ( .A(n_57), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_58), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_59), .B(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_SL g758 ( .A1(n_60), .A2(n_253), .B1(n_628), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_61), .Y(n_709) );
INVx1_ASAP7_75t_L g449 ( .A(n_62), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_66), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_67), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_68), .A2(n_251), .B1(n_525), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_69), .A2(n_206), .B1(n_468), .B2(n_561), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_70), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_71), .B(n_329), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_72), .A2(n_163), .B1(n_478), .B2(n_530), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_73), .A2(n_197), .B1(n_641), .B2(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_75), .A2(n_188), .B1(n_287), .B2(n_303), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_77), .A2(n_158), .B1(n_399), .B2(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_78), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_79), .A2(n_152), .B1(n_338), .B2(n_498), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_80), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_81), .A2(n_117), .B1(n_305), .B2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_82), .A2(n_252), .B1(n_381), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_83), .A2(n_258), .B1(n_324), .B2(n_331), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_85), .A2(n_144), .B1(n_317), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_86), .A2(n_88), .B1(n_339), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_89), .A2(n_213), .B1(n_310), .B2(n_609), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_90), .A2(n_255), .B1(n_305), .B2(n_699), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_92), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_93), .A2(n_205), .B1(n_303), .B2(n_475), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_94), .A2(n_224), .B1(n_333), .B2(n_383), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_95), .Y(n_829) );
INVx1_ASAP7_75t_L g278 ( .A(n_96), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_97), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_98), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_99), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_100), .A2(n_191), .B1(n_610), .B2(n_673), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_101), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g274 ( .A(n_102), .Y(n_274) );
INVx1_ASAP7_75t_L g772 ( .A(n_104), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_106), .A2(n_257), .B1(n_395), .B2(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_107), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_108), .A2(n_233), .B1(n_317), .B2(n_539), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_109), .A2(n_180), .B1(n_352), .B2(n_468), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_110), .A2(n_119), .B1(n_539), .B2(n_673), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_111), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_112), .Y(n_546) );
INVx1_ASAP7_75t_L g397 ( .A(n_113), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_114), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_115), .A2(n_168), .B1(n_363), .B2(n_401), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_116), .A2(n_132), .B1(n_218), .B2(n_733), .C1(n_735), .C2(n_736), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_118), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_120), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_122), .A2(n_129), .B1(n_401), .B2(n_583), .Y(n_599) );
INVx1_ASAP7_75t_L g386 ( .A(n_123), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_124), .A2(n_219), .B1(n_471), .B2(n_478), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_125), .A2(n_181), .B1(n_625), .B2(n_628), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_127), .A2(n_210), .B1(n_482), .B2(n_484), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_128), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_130), .A2(n_262), .B1(n_609), .B2(n_610), .Y(n_608) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_131), .A2(n_706), .B1(n_737), .B2(n_738), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_131), .Y(n_737) );
INVx1_ASAP7_75t_L g622 ( .A(n_133), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_134), .A2(n_137), .B1(n_287), .B2(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g391 ( .A(n_135), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_136), .A2(n_246), .B1(n_482), .B2(n_628), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_138), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g400 ( .A1(n_139), .A2(n_185), .B1(n_192), .B2(n_357), .C1(n_401), .C2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_140), .A2(n_171), .B1(n_309), .B2(n_316), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_141), .A2(n_269), .B1(n_323), .B2(n_666), .C(n_728), .Y(n_727) );
AOI222xp33_ASAP7_75t_L g356 ( .A1(n_142), .A2(n_176), .B1(n_212), .B2(n_357), .C1(n_358), .C2(n_362), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_143), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_146), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_147), .A2(n_190), .B1(n_454), .B2(n_475), .Y(n_540) );
AND2x2_ASAP7_75t_L g277 ( .A(n_148), .B(n_278), .Y(n_277) );
AO22x1_ASAP7_75t_L g404 ( .A1(n_149), .A2(n_405), .B1(n_455), .B2(n_456), .Y(n_404) );
INVx1_ASAP7_75t_L g455 ( .A(n_149), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_151), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_155), .A2(n_161), .B1(n_725), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_157), .A2(n_248), .B1(n_577), .B2(n_578), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_160), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_162), .A2(n_237), .B1(n_333), .B2(n_338), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_164), .A2(n_263), .B1(n_628), .B2(n_808), .Y(n_807) );
AND2x6_ASAP7_75t_L g273 ( .A(n_165), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_165), .Y(n_784) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_166), .A2(n_227), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_167), .A2(n_256), .B1(n_316), .B2(n_372), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_169), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_170), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_172), .A2(n_201), .B1(n_402), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_173), .A2(n_228), .B1(n_472), .B2(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_174), .B(n_324), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_177), .A2(n_250), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g703 ( .A(n_178), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_179), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_182), .A2(n_260), .B1(n_344), .B2(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g822 ( .A(n_183), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_183), .A2(n_822), .B1(n_824), .B2(n_851), .Y(n_823) );
INVx1_ASAP7_75t_L g375 ( .A(n_184), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_186), .Y(n_591) );
INVx1_ASAP7_75t_L g403 ( .A(n_189), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_193), .A2(n_221), .B1(n_603), .B2(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_194), .B(n_598), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_195), .B(n_362), .Y(n_423) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_196), .A2(n_238), .B1(n_292), .B2(n_297), .Y(n_296) );
XOR2x2_ASAP7_75t_L g283 ( .A(n_198), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g452 ( .A(n_199), .Y(n_452) );
INVx1_ASAP7_75t_L g644 ( .A(n_200), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_202), .A2(n_245), .B1(n_333), .B2(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g555 ( .A(n_203), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_204), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_207), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_211), .A2(n_271), .B(n_279), .C(n_792), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_214), .B(n_380), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_215), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_216), .A2(n_264), .B1(n_335), .B2(n_358), .Y(n_694) );
INVx1_ASAP7_75t_L g623 ( .A(n_217), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_222), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_225), .Y(n_480) );
XOR2x2_ASAP7_75t_L g508 ( .A(n_226), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_227), .B(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_229), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_232), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_234), .A2(n_241), .B1(n_350), .B2(n_353), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_235), .Y(n_729) );
INVx1_ASAP7_75t_L g787 ( .A(n_238), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_239), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_240), .A2(n_265), .B1(n_323), .B2(n_329), .Y(n_322) );
INVx1_ASAP7_75t_L g515 ( .A(n_242), .Y(n_515) );
OA22x2_ASAP7_75t_L g653 ( .A1(n_243), .A2(n_654), .B1(n_655), .B2(n_679), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_243), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_244), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_249), .Y(n_659) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
INVx1_ASAP7_75t_L g631 ( .A(n_259), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_261), .A2(n_464), .B1(n_503), .B2(n_504), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_261), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_267), .Y(n_548) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_274), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g820 ( .A1(n_275), .A2(n_782), .B(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_650), .B1(n_777), .B2(n_778), .C(n_779), .Y(n_279) );
INVxp67_ASAP7_75t_L g777 ( .A(n_280), .Y(n_777) );
XOR2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_459), .Y(n_280) );
OAI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_404), .B1(n_457), .B2(n_458), .Y(n_281) );
INVx1_ASAP7_75t_L g457 ( .A(n_282), .Y(n_457) );
XOR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_366), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_283), .A2(n_652), .B1(n_653), .B2(n_680), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_283), .Y(n_652) );
NAND4xp75_ASAP7_75t_L g284 ( .A(n_285), .B(n_321), .C(n_342), .D(n_356), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_308), .Y(n_285) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_288), .Y(n_468) );
BUFx2_ASAP7_75t_SL g586 ( .A(n_288), .Y(n_586) );
INVx2_ASAP7_75t_L g710 ( .A(n_288), .Y(n_710) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_298), .Y(n_288) );
AND2x6_ASAP7_75t_L g352 ( .A(n_289), .B(n_327), .Y(n_352) );
AND2x4_ASAP7_75t_L g355 ( .A(n_289), .B(n_315), .Y(n_355) );
AND2x6_ASAP7_75t_L g357 ( .A(n_289), .B(n_341), .Y(n_357) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_290), .B(n_296), .Y(n_307) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g313 ( .A(n_291), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_291), .B(n_296), .Y(n_320) );
AND2x2_ASAP7_75t_L g337 ( .A(n_291), .B(n_300), .Y(n_337) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g314 ( .A(n_296), .Y(n_314) );
INVx1_ASAP7_75t_L g361 ( .A(n_296), .Y(n_361) );
AND2x4_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g345 ( .A(n_298), .B(n_313), .Y(n_345) );
AND2x4_ASAP7_75t_L g347 ( .A(n_298), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_298), .B(n_313), .Y(n_389) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g315 ( .A(n_299), .B(n_302), .Y(n_315) );
OR2x2_ASAP7_75t_L g328 ( .A(n_299), .B(n_302), .Y(n_328) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g341 ( .A(n_300), .B(n_302), .Y(n_341) );
AND2x2_ASAP7_75t_L g360 ( .A(n_301), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g429 ( .A(n_301), .Y(n_429) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
INVx4_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_304), .A2(n_467), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_621) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g472 ( .A(n_306), .Y(n_472) );
INVx2_ASAP7_75t_L g604 ( .A(n_306), .Y(n_604) );
BUFx3_ASAP7_75t_L g678 ( .A(n_306), .Y(n_678) );
AND2x4_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
AND2x6_ASAP7_75t_L g331 ( .A(n_307), .B(n_315), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_307), .B(n_315), .Y(n_378) );
INVx1_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g532 ( .A(n_310), .Y(n_532) );
INVx5_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g373 ( .A(n_311), .Y(n_373) );
INVx1_ASAP7_75t_L g483 ( .A(n_311), .Y(n_483) );
INVx2_ASAP7_75t_L g561 ( .A(n_311), .Y(n_561) );
INVx3_ASAP7_75t_L g577 ( .A(n_311), .Y(n_577) );
INVx4_ASAP7_75t_L g627 ( .A(n_311), .Y(n_627) );
INVx8_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_313), .B(n_315), .Y(n_441) );
INVx1_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx4f_ASAP7_75t_SL g444 ( .A(n_317), .Y(n_444) );
BUFx2_ASAP7_75t_L g533 ( .A(n_317), .Y(n_533) );
BUFx2_ASAP7_75t_L g578 ( .A(n_317), .Y(n_578) );
BUFx2_ASAP7_75t_L g628 ( .A(n_317), .Y(n_628) );
INVx6_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g484 ( .A(n_318), .Y(n_484) );
INVx1_ASAP7_75t_SL g838 ( .A(n_318), .Y(n_838) );
OR2x6_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
INVx1_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_322), .B(n_332), .Y(n_321) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g381 ( .A(n_325), .Y(n_381) );
INVx2_ASAP7_75t_L g523 ( .A(n_325), .Y(n_523) );
INVx2_ASAP7_75t_L g597 ( .A(n_325), .Y(n_597) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g411 ( .A(n_328), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g804 ( .A(n_330), .Y(n_804) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
BUFx4f_ASAP7_75t_L g598 ( .A(n_331), .Y(n_598) );
BUFx2_ASAP7_75t_L g666 ( .A(n_331), .Y(n_666) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g641 ( .A(n_334), .Y(n_641) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g525 ( .A(n_335), .Y(n_525) );
BUFx3_ASAP7_75t_L g583 ( .A(n_335), .Y(n_583) );
BUFx2_ASAP7_75t_L g664 ( .A(n_335), .Y(n_664) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x4_ASAP7_75t_L g359 ( .A(n_337), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g364 ( .A(n_337), .B(n_365), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_337), .B(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
BUFx2_ASAP7_75t_SL g614 ( .A(n_339), .Y(n_614) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_339), .Y(n_767) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g435 ( .A(n_340), .Y(n_435) );
INVx1_ASAP7_75t_L g434 ( .A(n_341), .Y(n_434) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_349), .Y(n_342) );
INVx1_ASAP7_75t_L g447 ( .A(n_344), .Y(n_447) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g539 ( .A(n_345), .Y(n_539) );
BUFx3_ASAP7_75t_L g559 ( .A(n_345), .Y(n_559) );
BUFx3_ASAP7_75t_L g634 ( .A(n_345), .Y(n_634) );
INVxp67_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g437 ( .A(n_347), .Y(n_437) );
BUFx2_ASAP7_75t_SL g475 ( .A(n_347), .Y(n_475) );
BUFx2_ASAP7_75t_L g566 ( .A(n_347), .Y(n_566) );
INVx1_ASAP7_75t_L g606 ( .A(n_347), .Y(n_606) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_347), .Y(n_635) );
BUFx3_ASAP7_75t_L g673 ( .A(n_347), .Y(n_673) );
BUFx3_ASAP7_75t_L g726 ( .A(n_347), .Y(n_726) );
AND2x2_ASAP7_75t_L g699 ( .A(n_348), .B(n_429), .Y(n_699) );
INVx2_ASAP7_75t_L g827 ( .A(n_350), .Y(n_827) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_SL g530 ( .A(n_351), .Y(n_530) );
INVx4_ASAP7_75t_L g564 ( .A(n_351), .Y(n_564) );
INVx2_ASAP7_75t_L g762 ( .A(n_351), .Y(n_762) );
INVx11_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx11_ASAP7_75t_L g396 ( .A(n_352), .Y(n_396) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_L g454 ( .A(n_354), .Y(n_454) );
INVx6_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g478 ( .A(n_355), .Y(n_478) );
BUFx3_ASAP7_75t_L g610 ( .A(n_355), .Y(n_610) );
BUFx3_ASAP7_75t_L g744 ( .A(n_355), .Y(n_744) );
BUFx3_ASAP7_75t_L g418 ( .A(n_357), .Y(n_418) );
INVx2_ASAP7_75t_SL g492 ( .A(n_357), .Y(n_492) );
INVx4_ASAP7_75t_L g514 ( .A(n_357), .Y(n_514) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_357), .Y(n_613) );
INVx2_ASAP7_75t_L g688 ( .A(n_357), .Y(n_688) );
INVx1_ASAP7_75t_L g494 ( .A(n_358), .Y(n_494) );
BUFx4f_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_359), .Y(n_401) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_359), .Y(n_519) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_359), .Y(n_735) );
BUFx2_ASAP7_75t_L g771 ( .A(n_359), .Y(n_771) );
INVx1_ASAP7_75t_L g365 ( .A(n_361), .Y(n_365) );
INVx1_ASAP7_75t_L g646 ( .A(n_362), .Y(n_646) );
BUFx4f_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g590 ( .A(n_363), .Y(n_590) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_364), .Y(n_498) );
XOR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_403), .Y(n_366) );
NAND4xp75_ASAP7_75t_L g367 ( .A(n_368), .B(n_374), .C(n_384), .D(n_400), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OA211x2_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_379), .C(n_382), .Y(n_374) );
OA211x2_ASAP7_75t_L g579 ( .A1(n_376), .A2(n_580), .B(n_581), .C(n_582), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g840 ( .A1(n_376), .A2(n_488), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_840) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_392), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_390), .B2(n_391), .Y(n_385) );
OAI221xp5_ASAP7_75t_SL g476 ( .A1(n_387), .A2(n_477), .B1(n_479), .B2(n_480), .C(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g722 ( .A(n_388), .Y(n_722) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_397), .B2(n_398), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx4_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
INVx4_ASAP7_75t_L g609 ( .A(n_396), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_396), .A2(n_453), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_396), .A2(n_477), .B1(n_718), .B2(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
INVx1_ASAP7_75t_L g660 ( .A(n_402), .Y(n_660) );
INVx2_ASAP7_75t_L g458 ( .A(n_404), .Y(n_458) );
INVx1_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
AND3x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_436), .C(n_445), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_416), .C(n_424), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_413), .B2(n_414), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
INVx2_ASAP7_75t_L g637 ( .A(n_410), .Y(n_637) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g547 ( .A(n_411), .Y(n_547) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_417), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g798 ( .A1(n_417), .A2(n_799), .B(n_800), .Y(n_798) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_430), .B2(n_431), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_426), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g554 ( .A(n_428), .Y(n_554) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g502 ( .A(n_432), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_433), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
BUFx2_ASAP7_75t_L g731 ( .A(n_433), .Y(n_731) );
OR2x6_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_442), .B2(n_443), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_440), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
BUFx2_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_617), .B1(n_618), .B2(n_649), .Y(n_459) );
INVx1_ASAP7_75t_L g649 ( .A(n_460), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_505), .B2(n_616), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_465), .B(n_485), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
OAI221xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_469), .B1(n_470), .B2(n_473), .C(n_474), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
BUFx3_ASAP7_75t_L g675 ( .A(n_468), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_470), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
OAI221xp5_ASAP7_75t_SL g833 ( .A1(n_470), .A2(n_834), .B1(n_835), .B2(n_836), .C(n_837), .Y(n_833) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g835 ( .A(n_475), .Y(n_835) );
OAI221xp5_ASAP7_75t_SL g826 ( .A1(n_477), .A2(n_827), .B1(n_828), .B2(n_829), .C(n_830), .Y(n_826) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_491), .C(n_499), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_490), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_490), .A2(n_637), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B1(n_494), .B2(n_495), .C(n_496), .Y(n_491) );
OAI222xp33_ASAP7_75t_L g846 ( .A1(n_492), .A2(n_494), .B1(n_847), .B2(n_848), .C1(n_849), .C2(n_850), .Y(n_846) );
OAI222xp33_ASAP7_75t_L g657 ( .A1(n_494), .A2(n_512), .B1(n_658), .B2(n_659), .C1(n_660), .C2(n_661), .Y(n_657) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g736 ( .A(n_498), .Y(n_736) );
INVx2_ASAP7_75t_L g849 ( .A(n_498), .Y(n_849) );
INVx1_ASAP7_75t_L g616 ( .A(n_505), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_569), .B2(n_570), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_541), .B1(n_542), .B2(n_568), .Y(n_507) );
INVx2_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
NAND3x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_526), .C(n_534), .Y(n_509) );
NOR2x1_ASAP7_75t_SL g510 ( .A(n_511), .B(n_520), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_515), .B(n_516), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI222xp33_ASAP7_75t_L g642 ( .A1(n_514), .A2(n_643), .B1(n_644), .B2(n_645), .C1(n_646), .C2(n_647), .Y(n_642) );
BUFx2_ASAP7_75t_L g734 ( .A(n_514), .Y(n_734) );
INVx1_ASAP7_75t_L g643 ( .A(n_517), .Y(n_643) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .C(n_524), .Y(n_520) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_567), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_556), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .C(n_552), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_554), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
BUFx3_ASAP7_75t_L g669 ( .A(n_559), .Y(n_669) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_561), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_572), .B1(n_592), .B2(n_615), .Y(n_570) );
INVx3_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_591), .Y(n_572) );
NAND4xp75_ASAP7_75t_L g573 ( .A(n_574), .B(n_579), .C(n_584), .D(n_588), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g615 ( .A(n_593), .Y(n_615) );
NAND4xp75_ASAP7_75t_L g594 ( .A(n_595), .B(n_600), .C(n_607), .D(n_612), .Y(n_594) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_596), .B(n_599), .Y(n_595) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g648 ( .A(n_620), .Y(n_648) );
OR4x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_629), .C(n_636), .D(n_642), .Y(n_620) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_627), .Y(n_759) );
INVxp67_ASAP7_75t_L g715 ( .A(n_628), .Y(n_715) );
BUFx4f_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g832 ( .A(n_634), .Y(n_832) );
INVx1_ASAP7_75t_L g778 ( .A(n_650), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_681), .B1(n_775), .B2(n_776), .Y(n_650) );
INVx1_ASAP7_75t_L g775 ( .A(n_651), .Y(n_775) );
INVx1_ASAP7_75t_L g680 ( .A(n_653), .Y(n_680) );
INVx2_ASAP7_75t_L g679 ( .A(n_655), .Y(n_679) );
NAND3x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_667), .C(n_671), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_662), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g776 ( .A(n_681), .Y(n_776) );
XOR2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_704), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_703), .Y(n_684) );
NAND2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_695), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_691), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B(n_690), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .C(n_694), .Y(n_691) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_739), .B1(n_773), .B2(n_774), .Y(n_704) );
INVx1_ASAP7_75t_L g773 ( .A(n_705), .Y(n_773) );
INVx1_ASAP7_75t_L g738 ( .A(n_706), .Y(n_738) );
AND4x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_716), .C(n_727), .D(n_732), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_712), .Y(n_707) );
INVx3_ASAP7_75t_L g812 ( .A(n_710), .Y(n_812) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_717), .B(n_720), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g768 ( .A1(n_734), .A2(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g774 ( .A(n_739), .Y(n_774) );
XNOR2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_754), .Y(n_739) );
XOR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_753), .Y(n_740) );
NAND4xp75_ASAP7_75t_L g741 ( .A(n_742), .B(n_746), .C(n_749), .D(n_752), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
XOR2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_772), .Y(n_754) );
NOR4xp75_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .C(n_764), .D(n_768), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_SL g845 ( .A(n_767), .Y(n_845) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
NOR2x1_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .Y(n_780) );
OR2x2_ASAP7_75t_SL g854 ( .A(n_781), .B(n_786), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_783), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_783), .B(n_818), .Y(n_821) );
CKINVDCx16_ASAP7_75t_R g818 ( .A(n_784), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
OAI322xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_814), .A3(n_815), .B1(n_819), .B2(n_822), .C1(n_823), .C2(n_852), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND3x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_805), .C(n_809), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g851 ( .A(n_824), .Y(n_851) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_839), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_833), .Y(n_825) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_SL g839 ( .A(n_840), .B(n_846), .Y(n_839) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_854), .Y(n_853) );
endmodule