module fake_ibex_1040_n_3542 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_568, n_52, n_448, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3542);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3542;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_2498;
wire n_2235;
wire n_1802;
wire n_1944;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2897;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_667;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_2837;
wire n_1840;
wire n_671;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_641;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_2707;
wire n_1929;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_2663;
wire n_1960;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2451;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3510;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_606;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2697;
wire n_2224;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2599;
wire n_974;
wire n_1036;
wire n_2076;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2829;
wire n_1255;
wire n_2036;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_3357;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_594;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_847;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1599;
wire n_712;
wire n_1539;
wire n_1400;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2612;
wire n_2193;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_2716;
wire n_3495;
wire n_863;
wire n_597;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_2439;
wire n_1925;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2985;
wire n_2045;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_634;
wire n_991;
wire n_961;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2920;
wire n_2087;
wire n_3290;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_648;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_722;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_1871;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2348;
wire n_2093;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_2867;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_2433;
wire n_2816;
wire n_1931;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_599;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2790;
wire n_1693;
wire n_698;
wire n_2034;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_632;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3380;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2618;
wire n_2357;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2302;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_3482;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_172),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_468),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_577),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_497),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_578),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_529),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_164),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_5),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_4),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_396),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_357),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_189),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_499),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_84),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_266),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_338),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_264),
.Y(n_610)
);

INVxp33_ASAP7_75t_R g611 ( 
.A(n_559),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_466),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_28),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_192),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_54),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_519),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_567),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_186),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_354),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_266),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_558),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_358),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_306),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_371),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_180),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_258),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_452),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_388),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_32),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_299),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_547),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_259),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_431),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_22),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_498),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_590),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_84),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_534),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_435),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_509),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_201),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_210),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_221),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_310),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_141),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_580),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_29),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_517),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_530),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_299),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_442),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_259),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_334),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_61),
.Y(n_656)
);

CKINVDCx14_ASAP7_75t_R g657 ( 
.A(n_355),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_188),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_575),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_569),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_478),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_232),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_560),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_122),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_119),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_524),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_23),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_545),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_231),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_592),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_206),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_279),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_323),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_97),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_168),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_114),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_165),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_143),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_471),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_337),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_400),
.Y(n_684)
);

BUFx5_ASAP7_75t_L g685 ( 
.A(n_460),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_555),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_331),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_446),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_447),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_238),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_233),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_413),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_582),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_187),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_488),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_294),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_510),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_327),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_42),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_428),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_528),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_61),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_97),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_539),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_106),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_24),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_194),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_485),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_472),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_220),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_156),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_4),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_249),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_591),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_167),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_451),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_490),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_81),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_293),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_109),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_564),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_277),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_500),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_96),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_221),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_436),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_307),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_269),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_276),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_132),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_332),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_99),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_520),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_208),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_50),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_562),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_197),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_508),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_34),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_533),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_412),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_116),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_210),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_411),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_568),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_583),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_104),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_571),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_95),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_134),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_525),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_141),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_133),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_60),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_65),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_224),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_220),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_344),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_83),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_502),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_231),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_44),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_255),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_255),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_418),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_314),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_553),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_226),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_153),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_208),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_109),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_169),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_101),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_280),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_258),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_275),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_36),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_586),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_434),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_356),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_395),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_43),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_275),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_304),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_170),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_543),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_554),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_351),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_546),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_518),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_484),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_303),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_563),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_93),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_492),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_41),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_40),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_336),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_556),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_182),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_250),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_503),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_223),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_286),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_382),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_257),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_302),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_190),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_354),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_198),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_527),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_189),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_566),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_359),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_87),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_576),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_387),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_286),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_536),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_102),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_78),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_15),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_362),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_475),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_433),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_516),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_108),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_104),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_62),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_565),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_235),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_409),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_70),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_496),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_342),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_514),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_473),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_63),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_60),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_470),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_115),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_459),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_391),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_116),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_522),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_235),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_103),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_493),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_147),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_437),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_48),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_20),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_389),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_504),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_374),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_55),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_507),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_32),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_424),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_372),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_550),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_584),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_242),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_241),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_146),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_217),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_52),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_444),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_119),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_479),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_66),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_276),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_513),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_64),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_587),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_300),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_323),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_238),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_541),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_535),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_398),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_262),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_340),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_247),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_146),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_538),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_570),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_511),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_343),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_588),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_557),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_28),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_183),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_456),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_273),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_133),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_14),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_251),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_40),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_350),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_260),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_245),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_405),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_22),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_369),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_573),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_106),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_390),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_526),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_150),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_406),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_303),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_37),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_117),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_122),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_126),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_325),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_46),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_523),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_549),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_361),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_333),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_289),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_489),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_544),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_531),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_155),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_271),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_13),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_506),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_296),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_295),
.Y(n_932)
);

BUFx2_ASAP7_75t_SL g933 ( 
.A(n_164),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_385),
.Y(n_934)
);

BUFx10_ASAP7_75t_L g935 ( 
.A(n_144),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_140),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_415),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_103),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_401),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_57),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_51),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_81),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_343),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_551),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_458),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_206),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_12),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_35),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_175),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_383),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_574),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_540),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_19),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_178),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_0),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_123),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_548),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_194),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_288),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_120),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_197),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_101),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_312),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_552),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_137),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_218),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_227),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_71),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_281),
.Y(n_969)
);

BUFx10_ASAP7_75t_L g970 ( 
.A(n_215),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_183),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_16),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_10),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_12),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_272),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_31),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_572),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_71),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_370),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_118),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_234),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_213),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_11),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_162),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_512),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_505),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_329),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_515),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_521),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_95),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_561),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_198),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_142),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_86),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_241),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_244),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_256),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_137),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_161),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_426),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_425),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_796),
.B(n_0),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_693),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_802),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_847),
.B(n_1),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_802),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_847),
.B(n_1),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_639),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_837),
.B(n_2),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_639),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_807),
.B(n_2),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_639),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_802),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_729),
.B(n_3),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_867),
.B(n_3),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_867),
.B(n_5),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_607),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_893),
.B(n_6),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_893),
.B(n_6),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_802),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_607),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_605),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_894),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_894),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_657),
.B(n_7),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_759),
.B(n_7),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_999),
.B(n_8),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_820),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_894),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_605),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_837),
.B(n_8),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_894),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_939),
.B(n_9),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_675),
.B(n_9),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_897),
.B(n_10),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_945),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_897),
.B(n_613),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_647),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_613),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_673),
.Y(n_1041)
);

INVx5_ASAP7_75t_L g1042 ( 
.A(n_945),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_945),
.Y(n_1043)
);

CKINVDCx11_ASAP7_75t_R g1044 ( 
.A(n_644),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_647),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_939),
.B(n_11),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_626),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_703),
.B(n_13),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_673),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_766),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_671),
.Y(n_1051)
);

INVx5_ASAP7_75t_L g1052 ( 
.A(n_693),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_693),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_703),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_767),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_626),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_626),
.Y(n_1057)
);

AND2x6_ASAP7_75t_L g1058 ( 
.A(n_597),
.B(n_363),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_767),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_626),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_766),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_917),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_703),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_735),
.B(n_14),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_710),
.B(n_15),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_594),
.B(n_16),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_594),
.B(n_17),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_917),
.B(n_17),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_671),
.Y(n_1069)
);

AND2x6_ASAP7_75t_L g1070 ( 
.A(n_597),
.B(n_593),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_683),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_735),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_928),
.B(n_18),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_735),
.B(n_18),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_928),
.B(n_987),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_624),
.B(n_19),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_767),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_596),
.B(n_20),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_898),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_658),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_683),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_624),
.B(n_21),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_898),
.B(n_21),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_745),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_627),
.B(n_23),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_694),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_616),
.B(n_24),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_799),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_935),
.B(n_25),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_658),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_658),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_635),
.B(n_25),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_799),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_857),
.B(n_364),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_935),
.B(n_26),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_987),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_627),
.B(n_26),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_799),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_805),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_685),
.B(n_621),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_630),
.B(n_27),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_685),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_630),
.B(n_27),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_658),
.Y(n_1105)
);

BUFx12f_ASAP7_75t_L g1106 ( 
.A(n_935),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_732),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_685),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_631),
.B(n_29),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_955),
.B(n_30),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_631),
.B(n_30),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_955),
.B(n_31),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_732),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_732),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_642),
.B(n_648),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_732),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_633),
.B(n_33),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_782),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_650),
.B(n_33),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_685),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_782),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_694),
.B(n_34),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_719),
.Y(n_1123)
);

BUFx8_ASAP7_75t_L g1124 ( 
.A(n_719),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_663),
.B(n_35),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_955),
.B(n_36),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_782),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_595),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1034),
.A2(n_798),
.B1(n_633),
.B2(n_714),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1005),
.A2(n_798),
.B1(n_714),
.B2(n_700),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_855),
.B1(n_861),
.B2(n_700),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1012),
.A2(n_665),
.B1(n_677),
.B2(n_644),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1028),
.B(n_970),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1007),
.A2(n_861),
.B1(n_888),
.B2(n_855),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1041),
.B(n_970),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1049),
.B(n_970),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1013),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1015),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1022),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1002),
.A2(n_994),
.B1(n_677),
.B2(n_690),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1010),
.B(n_628),
.Y(n_1142)
);

AO22x2_ASAP7_75t_L g1143 ( 
.A1(n_1014),
.A2(n_1015),
.B1(n_1018),
.B2(n_1016),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1030),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_SL g1145 ( 
.A1(n_1066),
.A2(n_601),
.B1(n_602),
.B2(n_600),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1016),
.A2(n_920),
.B1(n_888),
.B2(n_608),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1010),
.B(n_628),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1054),
.B(n_629),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1018),
.A2(n_920),
.B1(n_610),
.B2(n_614),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1011),
.A2(n_690),
.B1(n_691),
.B2(n_665),
.Y(n_1150)
);

OAI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1026),
.A2(n_994),
.B1(n_706),
.B2(n_722),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1019),
.A2(n_611),
.B1(n_933),
.B2(n_715),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1027),
.A2(n_706),
.B1(n_722),
.B2(n_691),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1054),
.B(n_629),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1040),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1019),
.A2(n_618),
.B1(n_619),
.B2(n_604),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1067),
.A2(n_756),
.B1(n_757),
.B2(n_730),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1035),
.A2(n_620),
.B1(n_649),
.B2(n_643),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1076),
.A2(n_655),
.B1(n_656),
.B2(n_654),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1035),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_1083),
.A2(n_1086),
.B1(n_1102),
.B2(n_1098),
.Y(n_1161)
);

XOR2xp5_ASAP7_75t_L g1162 ( 
.A(n_1085),
.B(n_730),
.Y(n_1162)
);

OAI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1104),
.A2(n_666),
.B1(n_676),
.B2(n_662),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1068),
.A2(n_680),
.B1(n_681),
.B2(n_678),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1068),
.A2(n_698),
.B1(n_699),
.B2(n_696),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1073),
.A2(n_615),
.B1(n_764),
.B2(n_752),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1109),
.A2(n_757),
.B1(n_761),
.B2(n_756),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1072),
.B(n_725),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1072),
.B(n_632),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1080),
.B(n_632),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1111),
.A2(n_769),
.B1(n_794),
.B2(n_761),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1050),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1061),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_1037),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1063),
.A2(n_794),
.B1(n_810),
.B2(n_769),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1013),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1080),
.B(n_725),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1122),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1008),
.A2(n_705),
.B1(n_711),
.B2(n_702),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1073),
.A2(n_713),
.B1(n_718),
.B2(n_712),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1182)
);

OAI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1117),
.A2(n_827),
.B1(n_974),
.B2(n_810),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1079),
.A2(n_727),
.B1(n_728),
.B2(n_724),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1128),
.B(n_991),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1003),
.B(n_634),
.Y(n_1186)
);

AO22x2_ASAP7_75t_L g1187 ( 
.A1(n_1122),
.A2(n_815),
.B1(n_849),
.B2(n_788),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1106),
.A2(n_737),
.B1(n_739),
.B2(n_734),
.Y(n_1188)
);

NAND3x1_ASAP7_75t_L g1189 ( 
.A(n_1048),
.B(n_974),
.C(n_827),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1064),
.A2(n_996),
.B1(n_918),
.B2(n_995),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1044),
.A2(n_747),
.B1(n_750),
.B2(n_742),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1192)
);

AO22x2_ASAP7_75t_L g1193 ( 
.A1(n_1074),
.A2(n_623),
.B1(n_636),
.B2(n_609),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1095),
.A2(n_646),
.B1(n_652),
.B2(n_645),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1065),
.A2(n_754),
.B1(n_755),
.B2(n_753),
.Y(n_1195)
);

CKINVDCx11_ASAP7_75t_R g1196 ( 
.A(n_1075),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1025),
.A2(n_763),
.B1(n_770),
.B2(n_758),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1084),
.A2(n_773),
.B1(n_775),
.B2(n_771),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1199)
);

OR2x6_ASAP7_75t_L g1200 ( 
.A(n_1090),
.B(n_789),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1128),
.B(n_634),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1075),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1096),
.A2(n_674),
.B1(n_679),
.B2(n_669),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1110),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1055),
.A2(n_777),
.B1(n_780),
.B2(n_776),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1112),
.A2(n_784),
.B1(n_785),
.B2(n_783),
.Y(n_1206)
);

AO22x2_ASAP7_75t_L g1207 ( 
.A1(n_1126),
.A2(n_993),
.B1(n_997),
.B2(n_992),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1055),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1062),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1115),
.A2(n_1124),
.B1(n_1031),
.B2(n_1033),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1078),
.A2(n_797),
.B1(n_800),
.B2(n_792),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1097),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1124),
.A2(n_804),
.B1(n_809),
.B2(n_801),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1055),
.A2(n_814),
.B1(n_821),
.B2(n_812),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1059),
.B(n_842),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1009),
.A2(n_831),
.B1(n_835),
.B2(n_828),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1100),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1059),
.B(n_842),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1017),
.A2(n_998),
.B1(n_990),
.B2(n_707),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1059),
.A2(n_720),
.B1(n_731),
.B2(n_687),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1077),
.B(n_991),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1114),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_1094),
.B1(n_1099),
.B2(n_1089),
.Y(n_1223)
);

OA22x2_ASAP7_75t_L g1224 ( 
.A1(n_1017),
.A2(n_916),
.B1(n_927),
.B2(n_900),
.Y(n_1224)
);

AO22x2_ASAP7_75t_L g1225 ( 
.A1(n_1021),
.A2(n_980),
.B1(n_978),
.B2(n_749),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1077),
.B(n_1089),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1021),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1089),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1094),
.A2(n_762),
.B1(n_768),
.B2(n_743),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_SL g1230 ( 
.A(n_1039),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1046),
.A2(n_839),
.B1(n_841),
.B2(n_838),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1114),
.Y(n_1232)
);

AO22x2_ASAP7_75t_L g1233 ( 
.A1(n_1039),
.A2(n_774),
.B1(n_803),
.B2(n_772),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1114),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1088),
.A2(n_852),
.B1(n_856),
.B2(n_846),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1094),
.A2(n_806),
.B1(n_818),
.B2(n_808),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1116),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1116),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1116),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_822),
.B1(n_833),
.B2(n_829),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1099),
.A2(n_865),
.B1(n_872),
.B2(n_864),
.Y(n_1241)
);

AND2x2_ASAP7_75t_SL g1242 ( 
.A(n_1093),
.B(n_959),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1119),
.A2(n_1125),
.B1(n_1070),
.B2(n_1058),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1058),
.A2(n_876),
.B1(n_877),
.B2(n_874),
.Y(n_1244)
);

AO22x2_ASAP7_75t_L g1245 ( 
.A1(n_1045),
.A2(n_851),
.B1(n_858),
.B2(n_844),
.Y(n_1245)
);

AO22x2_ASAP7_75t_L g1246 ( 
.A1(n_1045),
.A2(n_866),
.B1(n_869),
.B2(n_863),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1058),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1051),
.B(n_1000),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1051),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1069),
.Y(n_1251)
);

AND2x2_ASAP7_75t_SL g1252 ( 
.A(n_1069),
.B(n_959),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1121),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1071),
.A2(n_882),
.B1(n_892),
.B2(n_878),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1071),
.B(n_1000),
.Y(n_1255)
);

AO22x2_ASAP7_75t_L g1256 ( 
.A1(n_1082),
.A2(n_883),
.B1(n_884),
.B2(n_871),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1058),
.A2(n_907),
.B1(n_914),
.B2(n_902),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1082),
.A2(n_922),
.B1(n_931),
.B2(n_915),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1121),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1127),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1070),
.A2(n_938),
.B1(n_941),
.B2(n_932),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1087),
.B(n_968),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1087),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1070),
.A2(n_943),
.B1(n_947),
.B2(n_942),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1123),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_R g1266 ( 
.A1(n_1123),
.A2(n_895),
.B1(n_896),
.B2(n_885),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1070),
.A2(n_953),
.B1(n_954),
.B2(n_949),
.Y(n_1267)
);

NAND2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1101),
.B(n_956),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1103),
.B(n_968),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1108),
.B(n_668),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1120),
.B(n_973),
.Y(n_1271)
);

NAND3x1_ASAP7_75t_L g1272 ( 
.A(n_1127),
.B(n_901),
.C(n_899),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1127),
.A2(n_961),
.B1(n_962),
.B2(n_958),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1004),
.Y(n_1274)
);

INVx8_ASAP7_75t_L g1275 ( 
.A(n_1004),
.Y(n_1275)
);

AO22x2_ASAP7_75t_L g1276 ( 
.A1(n_1004),
.A2(n_910),
.B1(n_912),
.B2(n_904),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1006),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1006),
.A2(n_965),
.B1(n_966),
.B2(n_963),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1047),
.A2(n_971),
.B1(n_975),
.B2(n_967),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1006),
.Y(n_1280)
);

AND2x2_ASAP7_75t_SL g1281 ( 
.A(n_1047),
.B(n_913),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1029),
.B(n_976),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1029),
.B(n_981),
.Y(n_1283)
);

OAI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1029),
.A2(n_936),
.B1(n_940),
.B2(n_923),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_982),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1038),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1038),
.B(n_983),
.Y(n_1287)
);

OA22x2_ASAP7_75t_L g1288 ( 
.A1(n_1042),
.A2(n_984),
.B1(n_946),
.B2(n_969),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1042),
.Y(n_1289)
);

AO22x2_ASAP7_75t_L g1290 ( 
.A1(n_1042),
.A2(n_972),
.B1(n_948),
.B2(n_670),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1043),
.A2(n_682),
.B1(n_697),
.B2(n_688),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1043),
.A2(n_790),
.B1(n_723),
.B2(n_726),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1043),
.A2(n_960),
.B1(n_889),
.B2(n_929),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1047),
.A2(n_740),
.B1(n_760),
.B2(n_721),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1056),
.A2(n_782),
.B1(n_929),
.B2(n_889),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_1056),
.A2(n_786),
.B1(n_793),
.B2(n_781),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1056),
.Y(n_1297)
);

AO22x2_ASAP7_75t_L g1298 ( 
.A1(n_1057),
.A2(n_823),
.B1(n_834),
.B2(n_813),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1057),
.B(n_889),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1057),
.B(n_843),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1060),
.A2(n_929),
.B1(n_960),
.B2(n_889),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1060),
.A2(n_960),
.B1(n_929),
.B2(n_868),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1060),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1081),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1081),
.A2(n_960),
.B1(n_870),
.B2(n_879),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1081),
.A2(n_880),
.B1(n_881),
.B2(n_854),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1091),
.B(n_805),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1091),
.A2(n_903),
.B1(n_908),
.B2(n_890),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1091),
.Y(n_1309)
);

NAND3x1_ASAP7_75t_L g1310 ( 
.A(n_1092),
.B(n_911),
.C(n_909),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1092),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1092),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1105),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1105),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1105),
.A2(n_952),
.B1(n_957),
.B2(n_924),
.Y(n_1315)
);

OA22x2_ASAP7_75t_L g1316 ( 
.A1(n_1107),
.A2(n_1001),
.B1(n_625),
.B2(n_716),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1107),
.Y(n_1317)
);

AO22x2_ASAP7_75t_L g1318 ( 
.A1(n_1107),
.A2(n_692),
.B1(n_795),
.B2(n_621),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1113),
.A2(n_599),
.B1(n_603),
.B2(n_598),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1113),
.A2(n_612),
.B1(n_617),
.B2(n_606),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1113),
.A2(n_637),
.B1(n_638),
.B2(n_622),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1118),
.B(n_850),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1118),
.A2(n_692),
.B1(n_921),
.B2(n_795),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1118),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1013),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1020),
.A2(n_921),
.B1(n_850),
.B2(n_816),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1036),
.A2(n_641),
.B1(n_651),
.B2(n_640),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1020),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1020),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1023),
.A2(n_824),
.B1(n_830),
.B2(n_684),
.Y(n_1330)
);

AO22x2_ASAP7_75t_L g1331 ( 
.A1(n_1023),
.A2(n_950),
.B1(n_989),
.B2(n_930),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1023),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1024),
.A2(n_659),
.B1(n_660),
.B2(n_653),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1036),
.B(n_661),
.Y(n_1334)
);

INVx8_ASAP7_75t_L g1335 ( 
.A(n_1024),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1024),
.A2(n_667),
.B1(n_672),
.B2(n_664),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1032),
.A2(n_988),
.B1(n_686),
.B2(n_695),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1032),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1032),
.A2(n_689),
.B1(n_704),
.B2(n_701),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1036),
.B(n_708),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1022),
.Y(n_1341)
);

OA22x2_ASAP7_75t_L g1342 ( 
.A1(n_1008),
.A2(n_717),
.B1(n_733),
.B2(n_709),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1052),
.B(n_736),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1307),
.Y(n_1344)
);

INVxp33_ASAP7_75t_SL g1345 ( 
.A(n_1132),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1174),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1140),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1175),
.B(n_738),
.Y(n_1348)
);

AND2x2_ASAP7_75t_SL g1349 ( 
.A(n_1135),
.B(n_37),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1202),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1142),
.B(n_741),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_SL g1352 ( 
.A(n_1247),
.B(n_986),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1244),
.B(n_744),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1204),
.B(n_985),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1139),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1160),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1168),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1147),
.Y(n_1358)
);

XOR2xp5_ASAP7_75t_L g1359 ( 
.A(n_1162),
.B(n_1152),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1144),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1178),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1269),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1227),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1250),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1196),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1133),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1251),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1155),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1263),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1265),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1148),
.B(n_746),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1249),
.B(n_748),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1247),
.B(n_751),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1131),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1212),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1172),
.Y(n_1376)
);

XOR2x2_ASAP7_75t_L g1377 ( 
.A(n_1189),
.B(n_38),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1243),
.A2(n_778),
.B(n_765),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1186),
.B(n_779),
.Y(n_1379)
);

XOR2x2_ASAP7_75t_L g1380 ( 
.A(n_1176),
.B(n_38),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1173),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1209),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1341),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

AND2x6_ASAP7_75t_L g1385 ( 
.A(n_1257),
.B(n_685),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1219),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1219),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1154),
.B(n_787),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1217),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1225),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1270),
.A2(n_811),
.B(n_791),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1225),
.Y(n_1392)
);

XOR2xp5_ASAP7_75t_L g1393 ( 
.A(n_1152),
.B(n_39),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1169),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_1296),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1299),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1299),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1233),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1233),
.Y(n_1399)
);

XOR2xp5_ASAP7_75t_L g1400 ( 
.A(n_1130),
.B(n_39),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1245),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1245),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1129),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1331),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1246),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1261),
.B(n_817),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1255),
.B(n_819),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1246),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1264),
.B(n_825),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1222),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1170),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1256),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1256),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1143),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1143),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1179),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1193),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1275),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1146),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1185),
.B(n_826),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1191),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1193),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1232),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1203),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1200),
.B(n_41),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1203),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1207),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1207),
.Y(n_1428)
);

XOR2xp5_ASAP7_75t_L g1429 ( 
.A(n_1149),
.B(n_42),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1201),
.B(n_832),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1288),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1136),
.B(n_43),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1267),
.B(n_836),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1316),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1252),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1134),
.B(n_840),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1200),
.B(n_845),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1208),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1192),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_SL g1440 ( 
.A(n_1194),
.B(n_848),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1161),
.B(n_853),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1230),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1137),
.B(n_1210),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1199),
.Y(n_1444)
);

XNOR2x2_ASAP7_75t_L g1445 ( 
.A(n_1190),
.B(n_44),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1258),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1226),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1205),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1282),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1283),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1215),
.B(n_859),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1218),
.B(n_860),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1271),
.A2(n_873),
.B(n_862),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1234),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1237),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1285),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1151),
.B(n_45),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1224),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1296),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1214),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1221),
.B(n_875),
.Y(n_1461)
);

NOR2xp67_ASAP7_75t_L g1462 ( 
.A(n_1274),
.B(n_365),
.Y(n_1462)
);

XOR2xp5_ASAP7_75t_L g1463 ( 
.A(n_1157),
.B(n_1167),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1197),
.B(n_1198),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1228),
.B(n_886),
.Y(n_1465)
);

XNOR2xp5_ASAP7_75t_L g1466 ( 
.A(n_1171),
.B(n_45),
.Y(n_1466)
);

AND2x2_ASAP7_75t_SL g1467 ( 
.A(n_1281),
.B(n_46),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1298),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1206),
.B(n_887),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_R g1470 ( 
.A(n_1182),
.B(n_891),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1289),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1298),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1318),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1318),
.Y(n_1474)
);

XNOR2xp5_ASAP7_75t_L g1475 ( 
.A(n_1183),
.B(n_47),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1275),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1276),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1164),
.B(n_905),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1331),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1290),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1290),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1334),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1340),
.Y(n_1484)
);

XOR2xp5_ASAP7_75t_L g1485 ( 
.A(n_1153),
.B(n_47),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1242),
.B(n_906),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1180),
.B(n_919),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1238),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1300),
.Y(n_1489)
);

XOR2xp5_ASAP7_75t_L g1490 ( 
.A(n_1141),
.B(n_48),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1187),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1239),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1187),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1292),
.A2(n_926),
.B(n_925),
.Y(n_1494)
);

XNOR2xp5_ASAP7_75t_L g1495 ( 
.A(n_1150),
.B(n_49),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1306),
.Y(n_1496)
);

INVxp33_ASAP7_75t_L g1497 ( 
.A(n_1211),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1156),
.B(n_1158),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1287),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1184),
.B(n_979),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1284),
.Y(n_1501)
);

XOR2xp5_ASAP7_75t_L g1502 ( 
.A(n_1166),
.B(n_1188),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1190),
.B(n_934),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1286),
.B(n_366),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1165),
.B(n_1181),
.Y(n_1505)
);

NAND2xp33_ASAP7_75t_SL g1506 ( 
.A(n_1343),
.B(n_937),
.Y(n_1506)
);

INVx3_ASAP7_75t_R g1507 ( 
.A(n_1248),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1213),
.B(n_977),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1342),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1291),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1279),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1253),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1216),
.B(n_944),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1291),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1220),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1229),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1231),
.B(n_951),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1236),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1273),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1240),
.Y(n_1520)
);

XNOR2x2_ASAP7_75t_L g1521 ( 
.A(n_1166),
.B(n_49),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1259),
.B(n_1260),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1323),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1235),
.B(n_964),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1315),
.Y(n_1525)
);

NOR2xp67_ASAP7_75t_L g1526 ( 
.A(n_1277),
.B(n_367),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1310),
.A2(n_685),
.B(n_373),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1280),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1294),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1223),
.B(n_685),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1330),
.B(n_368),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1308),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1319),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1254),
.Y(n_1534)
);

INVxp33_ASAP7_75t_L g1535 ( 
.A(n_1320),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1241),
.B(n_375),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1305),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1327),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1333),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1278),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1195),
.B(n_376),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1326),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1321),
.B(n_50),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1335),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1322),
.Y(n_1545)
);

BUFx5_ASAP7_75t_L g1546 ( 
.A(n_1304),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1145),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1337),
.B(n_51),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1159),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_SL g1550 ( 
.A(n_1163),
.B(n_377),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1272),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1293),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1309),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1268),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1302),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1266),
.Y(n_1556)
);

XOR2xp5_ASAP7_75t_L g1557 ( 
.A(n_1339),
.B(n_52),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1295),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1314),
.B(n_53),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1335),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1325),
.B(n_53),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1312),
.B(n_54),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1301),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1336),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1317),
.Y(n_1565)
);

XOR2xp5_ASAP7_75t_L g1566 ( 
.A(n_1324),
.B(n_55),
.Y(n_1566)
);

XNOR2xp5_ASAP7_75t_L g1567 ( 
.A(n_1297),
.B(n_56),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1303),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1138),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1311),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1313),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1138),
.B(n_378),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1338),
.Y(n_1573)
);

XOR2xp5_ASAP7_75t_L g1574 ( 
.A(n_1177),
.B(n_56),
.Y(n_1574)
);

INVxp33_ASAP7_75t_L g1575 ( 
.A(n_1177),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1332),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1328),
.B(n_57),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1329),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1204),
.B(n_58),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1142),
.B(n_58),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1249),
.B(n_379),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1196),
.Y(n_1582)
);

INVx8_ASAP7_75t_L g1583 ( 
.A(n_1200),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1174),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1174),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1174),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1174),
.B(n_380),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1174),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1223),
.B(n_59),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1204),
.B(n_59),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1133),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1174),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1174),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1174),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1174),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1174),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1174),
.B(n_381),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1174),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1307),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1174),
.B(n_384),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1307),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1174),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1174),
.Y(n_1603)
);

AND2x6_ASAP7_75t_L g1604 ( 
.A(n_1243),
.B(n_386),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1174),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1204),
.B(n_62),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1174),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1174),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_SL g1609 ( 
.A(n_1200),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1174),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1247),
.B(n_392),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1174),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1174),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1174),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1174),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1133),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1204),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1174),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1174),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1307),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1174),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1174),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1307),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1243),
.A2(n_589),
.B(n_394),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1174),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1275),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1247),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1174),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1174),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1244),
.B(n_393),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1174),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1174),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1174),
.B(n_397),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1355),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1356),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1544),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1617),
.B(n_63),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1346),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1363),
.A2(n_402),
.B(n_399),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1365),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1544),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1617),
.B(n_64),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1463),
.B(n_1556),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1364),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1349),
.B(n_65),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1374),
.B(n_66),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1584),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1416),
.B(n_67),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1351),
.B(n_67),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1585),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1425),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1544),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1351),
.B(n_68),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1414),
.B(n_68),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1586),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1415),
.B(n_69),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1569),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1386),
.B(n_69),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1367),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1627),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1588),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1592),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1371),
.B(n_70),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1387),
.B(n_72),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1593),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1390),
.B(n_72),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1418),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1392),
.B(n_73),
.Y(n_1670)
);

BUFx4f_ASAP7_75t_SL g1671 ( 
.A(n_1418),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1371),
.B(n_73),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1398),
.B(n_74),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1418),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1425),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1476),
.B(n_74),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1624),
.A2(n_404),
.B(n_403),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1354),
.B(n_1503),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1524),
.B(n_75),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1524),
.B(n_75),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1399),
.B(n_76),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1443),
.B(n_76),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1478),
.B(n_77),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1562),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1369),
.Y(n_1685)
);

AND2x2_ASAP7_75t_SL g1686 ( 
.A(n_1467),
.B(n_77),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1478),
.B(n_78),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1425),
.B(n_79),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1401),
.B(n_79),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1594),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1562),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1358),
.B(n_80),
.Y(n_1692)
);

AND2x6_ASAP7_75t_L g1693 ( 
.A(n_1459),
.B(n_407),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1394),
.B(n_80),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1352),
.B(n_585),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1469),
.B(n_82),
.Y(n_1696)
);

OR2x2_ASAP7_75t_SL g1697 ( 
.A(n_1457),
.B(n_82),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1595),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1411),
.B(n_83),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1370),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1626),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1596),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1402),
.B(n_85),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1598),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1602),
.Y(n_1706)
);

AND2x6_ASAP7_75t_L g1707 ( 
.A(n_1468),
.B(n_408),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1505),
.B(n_85),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1441),
.B(n_1511),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1347),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1464),
.B(n_86),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1360),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1368),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1604),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1376),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1603),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1404),
.B(n_87),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1437),
.B(n_88),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1435),
.B(n_88),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1605),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1437),
.B(n_89),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1432),
.B(n_89),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1417),
.B(n_90),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1405),
.B(n_90),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1372),
.B(n_91),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1408),
.B(n_91),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1412),
.B(n_92),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1381),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1382),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1480),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1580),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1372),
.B(n_92),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1513),
.B(n_93),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1413),
.B(n_94),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1514),
.B(n_94),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1395),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1555),
.A2(n_414),
.B(n_410),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1407),
.B(n_96),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1442),
.B(n_98),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1383),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1580),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1742)
);

OR2x2_ASAP7_75t_SL g1743 ( 
.A(n_1359),
.B(n_98),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1426),
.B(n_99),
.Y(n_1744)
);

AND2x2_ASAP7_75t_SL g1745 ( 
.A(n_1611),
.B(n_100),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1560),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1607),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1352),
.B(n_416),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1427),
.B(n_100),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1579),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1608),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1428),
.B(n_102),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1407),
.B(n_105),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1373),
.B(n_1624),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1492),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1610),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1590),
.B(n_105),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1546),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1604),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1472),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1606),
.B(n_107),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1501),
.B(n_107),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1362),
.B(n_108),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1515),
.B(n_110),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1583),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1546),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1604),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1612),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1516),
.B(n_110),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1518),
.B(n_111),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1613),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1614),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1520),
.B(n_111),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1396),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1499),
.B(n_112),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1465),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1471),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1546),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1388),
.B(n_112),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1350),
.B(n_113),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1534),
.B(n_113),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1546),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1615),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1618),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1547),
.B(n_114),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1546),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1549),
.B(n_115),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1496),
.B(n_117),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1373),
.B(n_581),
.Y(n_1789)
);

BUFx5_ASAP7_75t_L g1790 ( 
.A(n_1604),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1513),
.B(n_118),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1583),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1473),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1471),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1583),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1397),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1465),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1535),
.B(n_120),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1410),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1619),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1500),
.B(n_1498),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1449),
.B(n_121),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1514),
.B(n_121),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1440),
.A2(n_1540),
.B1(n_1479),
.B2(n_1477),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1458),
.B(n_123),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1450),
.B(n_1456),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1621),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1622),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1508),
.B(n_1497),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1423),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1483),
.B(n_124),
.Y(n_1811)
);

AND2x2_ASAP7_75t_SL g1812 ( 
.A(n_1611),
.B(n_124),
.Y(n_1812)
);

AND2x2_ASAP7_75t_SL g1813 ( 
.A(n_1440),
.B(n_125),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1484),
.B(n_125),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1625),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1436),
.B(n_126),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1474),
.B(n_127),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1454),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1455),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1495),
.B(n_127),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1451),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1574),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1628),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1488),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1512),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1486),
.B(n_128),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1528),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1582),
.B(n_128),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1375),
.B(n_129),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1344),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1491),
.B(n_129),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1629),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1493),
.B(n_130),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1599),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1481),
.B(n_417),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1589),
.B(n_130),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1482),
.B(n_419),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1565),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1431),
.B(n_131),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1389),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1601),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1620),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1509),
.B(n_1554),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1553),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1577),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1525),
.B(n_131),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1623),
.Y(n_1847)
);

NAND2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1439),
.B(n_1444),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1558),
.A2(n_421),
.B(n_420),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1570),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1537),
.A2(n_423),
.B(n_422),
.Y(n_1851)
);

INVx4_ASAP7_75t_L g1852 ( 
.A(n_1385),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1466),
.B(n_132),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1568),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1475),
.B(n_134),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1447),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1438),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1451),
.B(n_135),
.Y(n_1858)
);

AND2x2_ASAP7_75t_SL g1859 ( 
.A(n_1550),
.B(n_135),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1564),
.B(n_136),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1571),
.Y(n_1861)
);

INVxp33_ASAP7_75t_L g1862 ( 
.A(n_1379),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1573),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1559),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1391),
.B(n_136),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1486),
.B(n_138),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1542),
.B(n_1631),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1391),
.B(n_138),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1632),
.B(n_139),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1561),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1581),
.A2(n_429),
.B(n_427),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1581),
.A2(n_432),
.B(n_430),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1385),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1494),
.B(n_139),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1487),
.B(n_140),
.Y(n_1875)
);

AND2x2_ASAP7_75t_SL g1876 ( 
.A(n_1550),
.B(n_142),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1494),
.B(n_143),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1384),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1545),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1420),
.B(n_144),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1576),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1578),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1434),
.B(n_145),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1563),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1551),
.B(n_145),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1357),
.Y(n_1886)
);

INVxp67_ASAP7_75t_SL g1887 ( 
.A(n_1403),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1538),
.B(n_147),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1517),
.B(n_148),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1552),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1529),
.B(n_438),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1385),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1353),
.B(n_148),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1539),
.B(n_149),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1523),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1489),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1361),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1543),
.B(n_149),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1609),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1385),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1430),
.B(n_150),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1532),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1630),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1406),
.B(n_151),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1409),
.B(n_151),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1548),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1522),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1348),
.B(n_152),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1522),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1490),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1531),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1485),
.B(n_152),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1530),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1541),
.B(n_153),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1400),
.Y(n_1915)
);

BUFx8_ASAP7_75t_L g1916 ( 
.A(n_1609),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1433),
.B(n_1452),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1429),
.B(n_154),
.Y(n_1918)
);

NOR2xp67_ASAP7_75t_L g1919 ( 
.A(n_1366),
.B(n_154),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1393),
.B(n_155),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1531),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1445),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1461),
.B(n_156),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1521),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1587),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1597),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1572),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1377),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1600),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1536),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1633),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1462),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1507),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1527),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1527),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1502),
.B(n_157),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1557),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1419),
.B(n_157),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1453),
.A2(n_440),
.B(n_439),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1462),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1504),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1519),
.B(n_158),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1504),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1526),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1566),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_SL g1946 ( 
.A(n_1421),
.B(n_1448),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1446),
.B(n_158),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1533),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1380),
.B(n_159),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1575),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1378),
.A2(n_443),
.B(n_441),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1567),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1460),
.B(n_159),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1526),
.B(n_160),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1506),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1470),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1345),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1591),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1616),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1374),
.B(n_160),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1617),
.B(n_161),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1617),
.B(n_162),
.Y(n_1962)
);

AND2x2_ASAP7_75t_SL g1963 ( 
.A(n_1467),
.B(n_163),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1374),
.B(n_163),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1363),
.A2(n_448),
.B(n_445),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1363),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1617),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1374),
.B(n_165),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1617),
.B(n_166),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1617),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1617),
.B(n_166),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1970),
.B(n_167),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1644),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1967),
.B(n_168),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1709),
.B(n_169),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1657),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1684),
.Y(n_1977)
);

OR2x6_ASAP7_75t_L g1978 ( 
.A(n_1765),
.B(n_170),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1636),
.Y(n_1979)
);

BUFx4f_ASAP7_75t_L g1980 ( 
.A(n_1686),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1644),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1709),
.B(n_171),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1660),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1906),
.B(n_171),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1660),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1682),
.B(n_1801),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1637),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1671),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1685),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1636),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1685),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1765),
.B(n_172),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1745),
.B(n_449),
.Y(n_1993)
);

AND2x6_ASAP7_75t_L g1994 ( 
.A(n_1714),
.B(n_1759),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1957),
.B(n_1862),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1682),
.B(n_173),
.Y(n_1996)
);

CKINVDCx6p67_ASAP7_75t_R g1997 ( 
.A(n_1701),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1765),
.B(n_1792),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1700),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1852),
.B(n_173),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1643),
.B(n_174),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1745),
.B(n_450),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1711),
.B(n_174),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1686),
.B(n_175),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1792),
.B(n_176),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1700),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1862),
.B(n_176),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1792),
.B(n_177),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1963),
.B(n_177),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1963),
.B(n_178),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1708),
.B(n_179),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1820),
.B(n_179),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1671),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1853),
.B(n_180),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_SL g2015 ( 
.A(n_1812),
.B(n_453),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1640),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1669),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1966),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1966),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1879),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1669),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1684),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1896),
.B(n_181),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1896),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1879),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1916),
.Y(n_2026)
);

BUFx3_ASAP7_75t_L g2027 ( 
.A(n_1916),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1855),
.B(n_181),
.Y(n_2028)
);

NAND2x1p5_ASAP7_75t_L g2029 ( 
.A(n_1795),
.B(n_1669),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1795),
.Y(n_2030)
);

NAND2x1p5_ASAP7_75t_L g2031 ( 
.A(n_1795),
.B(n_182),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1669),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_SL g2033 ( 
.A(n_1812),
.B(n_184),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1636),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1879),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1715),
.Y(n_2036)
);

AND2x6_ASAP7_75t_L g2037 ( 
.A(n_1714),
.B(n_184),
.Y(n_2037)
);

NAND2x1_ASAP7_75t_L g2038 ( 
.A(n_1636),
.B(n_454),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1742),
.B(n_185),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1652),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1715),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1763),
.B(n_185),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1916),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1728),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1728),
.Y(n_2045)
);

INVx5_ASAP7_75t_L g2046 ( 
.A(n_1652),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1742),
.B(n_186),
.Y(n_2047)
);

INVx4_ASAP7_75t_L g2048 ( 
.A(n_1652),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1912),
.B(n_187),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1763),
.B(n_188),
.Y(n_2050)
);

INVx5_ASAP7_75t_L g2051 ( 
.A(n_1658),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_SL g2052 ( 
.A(n_1859),
.B(n_1876),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1776),
.B(n_1797),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1637),
.Y(n_2054)
);

BUFx12f_ASAP7_75t_L g2055 ( 
.A(n_1640),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1641),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1912),
.B(n_190),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1731),
.B(n_191),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_1701),
.B(n_191),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1961),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1775),
.B(n_192),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1809),
.B(n_193),
.Y(n_2062)
);

AND2x2_ASAP7_75t_SL g2063 ( 
.A(n_1813),
.B(n_193),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_1971),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_1676),
.B(n_195),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1729),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1731),
.B(n_195),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_1856),
.B(n_196),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1856),
.B(n_196),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1729),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1740),
.Y(n_2071)
);

INVx2_ASAP7_75t_SL g2072 ( 
.A(n_1674),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1651),
.B(n_199),
.Y(n_2073)
);

NOR2xp67_ASAP7_75t_L g2074 ( 
.A(n_1714),
.B(n_455),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1658),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_1971),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_1821),
.B(n_199),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1675),
.B(n_200),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1821),
.B(n_200),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1775),
.B(n_201),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1741),
.B(n_1678),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1740),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1913),
.B(n_202),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1898),
.B(n_202),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1938),
.B(n_203),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1838),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1658),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_1658),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_1684),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1898),
.B(n_203),
.Y(n_2090)
);

BUFx12f_ASAP7_75t_L g2091 ( 
.A(n_1933),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_1887),
.B(n_204),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1942),
.B(n_204),
.Y(n_2093)
);

INVxp67_ASAP7_75t_L g2094 ( 
.A(n_1961),
.Y(n_2094)
);

NAND2x1p5_ASAP7_75t_L g2095 ( 
.A(n_1641),
.B(n_205),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1962),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1683),
.B(n_205),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1902),
.B(n_207),
.Y(n_2098)
);

BUFx4f_ASAP7_75t_SL g2099 ( 
.A(n_1933),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_1950),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1902),
.B(n_207),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1764),
.B(n_209),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1661),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_SL g2104 ( 
.A(n_1859),
.B(n_457),
.Y(n_2104)
);

INVx4_ASAP7_75t_L g2105 ( 
.A(n_1950),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1764),
.B(n_209),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1661),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1899),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_1945),
.B(n_211),
.Y(n_2109)
);

NAND2x1p5_ASAP7_75t_L g2110 ( 
.A(n_1674),
.B(n_211),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_1962),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1838),
.Y(n_2112)
);

BUFx2_ASAP7_75t_L g2113 ( 
.A(n_1969),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1843),
.B(n_212),
.Y(n_2114)
);

OR2x6_ASAP7_75t_L g2115 ( 
.A(n_1676),
.B(n_212),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1950),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1702),
.B(n_213),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1884),
.Y(n_2118)
);

CKINVDCx16_ASAP7_75t_R g2119 ( 
.A(n_1946),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1843),
.B(n_214),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1884),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_1950),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1661),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_1755),
.Y(n_2124)
);

BUFx4f_ASAP7_75t_L g2125 ( 
.A(n_1839),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_SL g2126 ( 
.A(n_1876),
.B(n_461),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_1969),
.Y(n_2127)
);

INVx6_ASAP7_75t_L g2128 ( 
.A(n_1933),
.Y(n_2128)
);

NAND2xp33_ASAP7_75t_L g2129 ( 
.A(n_1790),
.B(n_462),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1895),
.Y(n_2130)
);

BUFx3_ASAP7_75t_L g2131 ( 
.A(n_1755),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1895),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_1843),
.B(n_214),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1710),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_1948),
.Y(n_2135)
);

INVx3_ASAP7_75t_L g2136 ( 
.A(n_1661),
.Y(n_2136)
);

BUFx12f_ASAP7_75t_L g2137 ( 
.A(n_1828),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_SL g2138 ( 
.A(n_1813),
.B(n_463),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1665),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_1746),
.B(n_215),
.Y(n_2140)
);

INVx6_ASAP7_75t_L g2141 ( 
.A(n_1746),
.Y(n_2141)
);

BUFx4f_ASAP7_75t_L g2142 ( 
.A(n_1839),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1687),
.B(n_216),
.Y(n_2143)
);

NOR2x1p5_ASAP7_75t_L g2144 ( 
.A(n_1822),
.B(n_216),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1665),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1665),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1665),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1774),
.B(n_217),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1774),
.B(n_218),
.Y(n_2149)
);

NOR2xp67_ASAP7_75t_L g2150 ( 
.A(n_1714),
.B(n_464),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_SL g2151 ( 
.A(n_1717),
.B(n_219),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1958),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_1702),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1770),
.B(n_219),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1770),
.B(n_222),
.Y(n_2155)
);

OR2x6_ASAP7_75t_L g2156 ( 
.A(n_1885),
.B(n_222),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1773),
.B(n_223),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1773),
.B(n_224),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1696),
.B(n_225),
.Y(n_2159)
);

BUFx4f_ASAP7_75t_L g2160 ( 
.A(n_1839),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1889),
.B(n_225),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1890),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1890),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1702),
.B(n_226),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1889),
.B(n_227),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1710),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1806),
.B(n_228),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_1634),
.B(n_228),
.Y(n_2168)
);

INVx1_ASAP7_75t_SL g2169 ( 
.A(n_1642),
.Y(n_2169)
);

BUFx8_ASAP7_75t_SL g2170 ( 
.A(n_1688),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1702),
.B(n_229),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1635),
.B(n_229),
.Y(n_2172)
);

INVxp67_ASAP7_75t_SL g2173 ( 
.A(n_1684),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1865),
.B(n_230),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1712),
.Y(n_2175)
);

NAND2x1p5_ASAP7_75t_L g2176 ( 
.A(n_1744),
.B(n_230),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1777),
.Y(n_2177)
);

BUFx8_ASAP7_75t_L g2178 ( 
.A(n_1722),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1865),
.B(n_232),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_1885),
.B(n_233),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_1848),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_1638),
.B(n_234),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1777),
.Y(n_2183)
);

BUFx2_ASAP7_75t_L g2184 ( 
.A(n_1736),
.Y(n_2184)
);

INVx3_ASAP7_75t_L g2185 ( 
.A(n_1794),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1645),
.B(n_236),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_1730),
.Y(n_2187)
);

INVx3_ASAP7_75t_L g2188 ( 
.A(n_1794),
.Y(n_2188)
);

BUFx8_ASAP7_75t_SL g2189 ( 
.A(n_1956),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_1744),
.Y(n_2190)
);

OR2x6_ASAP7_75t_L g2191 ( 
.A(n_1885),
.B(n_236),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1868),
.B(n_237),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_1844),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1712),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_1937),
.B(n_237),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1868),
.B(n_239),
.Y(n_2196)
);

INVxp67_ASAP7_75t_SL g2197 ( 
.A(n_1691),
.Y(n_2197)
);

INVxp67_ASAP7_75t_L g2198 ( 
.A(n_1717),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_1744),
.B(n_239),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1826),
.B(n_1866),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1826),
.B(n_240),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1866),
.B(n_240),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1918),
.B(n_242),
.Y(n_2203)
);

BUFx2_ASAP7_75t_L g2204 ( 
.A(n_1749),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1713),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1733),
.B(n_243),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_1937),
.B(n_243),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1713),
.Y(n_2208)
);

BUFx3_ASAP7_75t_L g2209 ( 
.A(n_1848),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1647),
.B(n_244),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1810),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_1749),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1952),
.B(n_245),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1733),
.B(n_246),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1791),
.B(n_246),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1918),
.B(n_247),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_1650),
.B(n_1655),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1928),
.Y(n_2218)
);

AND2x2_ASAP7_75t_SL g2219 ( 
.A(n_1817),
.B(n_248),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_1844),
.Y(n_2220)
);

NOR2xp67_ASAP7_75t_L g2221 ( 
.A(n_1759),
.B(n_465),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1749),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1760),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1791),
.B(n_248),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1679),
.B(n_249),
.Y(n_2225)
);

CKINVDCx16_ASAP7_75t_R g2226 ( 
.A(n_1680),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1662),
.B(n_250),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1810),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1793),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_SL g2230 ( 
.A(n_1852),
.B(n_467),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1785),
.B(n_251),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1785),
.B(n_252),
.Y(n_2232)
);

NAND2x1_ASAP7_75t_L g2233 ( 
.A(n_1693),
.B(n_469),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1953),
.B(n_252),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1818),
.Y(n_2235)
);

INVx4_ASAP7_75t_L g2236 ( 
.A(n_1654),
.Y(n_2236)
);

BUFx4_ASAP7_75t_SL g2237 ( 
.A(n_1924),
.Y(n_2237)
);

OR2x6_ASAP7_75t_L g2238 ( 
.A(n_1836),
.B(n_253),
.Y(n_2238)
);

OR2x6_ASAP7_75t_L g2239 ( 
.A(n_1836),
.B(n_253),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1796),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1818),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1819),
.Y(n_2242)
);

INVx1_ASAP7_75t_SL g2243 ( 
.A(n_1718),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1953),
.B(n_254),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1819),
.Y(n_2245)
);

AND2x2_ASAP7_75t_SL g2246 ( 
.A(n_1817),
.B(n_254),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1663),
.B(n_256),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_SL g2248 ( 
.A(n_1852),
.B(n_474),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1824),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1796),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_1681),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1824),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1952),
.B(n_257),
.Y(n_2253)
);

OR2x6_ASAP7_75t_L g2254 ( 
.A(n_1654),
.B(n_260),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1667),
.B(n_261),
.Y(n_2255)
);

NOR2xp67_ASAP7_75t_SL g2256 ( 
.A(n_1759),
.B(n_261),
.Y(n_2256)
);

OR2x2_ASAP7_75t_L g2257 ( 
.A(n_1910),
.B(n_262),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1750),
.B(n_263),
.Y(n_2258)
);

INVxp67_ASAP7_75t_SL g2259 ( 
.A(n_1691),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1827),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1690),
.B(n_263),
.Y(n_2261)
);

BUFx12f_ASAP7_75t_L g2262 ( 
.A(n_1743),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1787),
.B(n_264),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_1915),
.B(n_265),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1827),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1787),
.B(n_265),
.Y(n_2266)
);

OR2x6_ASAP7_75t_L g2267 ( 
.A(n_1654),
.B(n_267),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_1698),
.B(n_267),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1854),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1703),
.B(n_1705),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1796),
.Y(n_2271)
);

OR2x6_ASAP7_75t_L g2272 ( 
.A(n_1656),
.B(n_1681),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_SL g2273 ( 
.A(n_1656),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1936),
.B(n_1920),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1721),
.B(n_268),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_1920),
.B(n_268),
.Y(n_2276)
);

AND2x2_ASAP7_75t_SL g2277 ( 
.A(n_1656),
.B(n_269),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_1706),
.B(n_270),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1781),
.B(n_270),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_1681),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1854),
.Y(n_2281)
);

NAND2x1p5_ASAP7_75t_L g2282 ( 
.A(n_1689),
.B(n_271),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_1689),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_1716),
.B(n_272),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_1697),
.B(n_273),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_1720),
.B(n_274),
.Y(n_2286)
);

NAND2x1p5_ASAP7_75t_L g2287 ( 
.A(n_1689),
.B(n_274),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_1747),
.B(n_277),
.Y(n_2288)
);

INVxp67_ASAP7_75t_L g2289 ( 
.A(n_1724),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_1844),
.Y(n_2290)
);

CKINVDCx8_ASAP7_75t_R g2291 ( 
.A(n_1759),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_SL g2292 ( 
.A(n_1900),
.B(n_476),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1867),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1781),
.B(n_278),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_1864),
.B(n_278),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1949),
.B(n_279),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1735),
.B(n_280),
.Y(n_2297)
);

NAND2x1p5_ASAP7_75t_L g2298 ( 
.A(n_1724),
.B(n_281),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_1724),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_1947),
.B(n_282),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1659),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1922),
.B(n_282),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1751),
.B(n_283),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_1756),
.B(n_1768),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_SL g2305 ( 
.A(n_1900),
.B(n_477),
.Y(n_2305)
);

NAND2x1_ASAP7_75t_L g2306 ( 
.A(n_1693),
.B(n_480),
.Y(n_2306)
);

INVxp67_ASAP7_75t_L g2307 ( 
.A(n_1757),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1845),
.B(n_283),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1659),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_1930),
.B(n_1649),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1861),
.Y(n_2311)
);

OR2x6_ASAP7_75t_L g2312 ( 
.A(n_1735),
.B(n_284),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_SL g2313 ( 
.A(n_1900),
.B(n_1790),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1845),
.B(n_284),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1861),
.Y(n_2315)
);

BUFx2_ASAP7_75t_L g2316 ( 
.A(n_1803),
.Y(n_2316)
);

CKINVDCx8_ASAP7_75t_R g2317 ( 
.A(n_1767),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_1757),
.Y(n_2318)
);

OR2x6_ASAP7_75t_L g2319 ( 
.A(n_1767),
.B(n_285),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_1761),
.Y(n_2320)
);

CKINVDCx8_ASAP7_75t_R g2321 ( 
.A(n_1767),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_1829),
.B(n_285),
.Y(n_2322)
);

AND2x6_ASAP7_75t_L g2323 ( 
.A(n_1767),
.B(n_287),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1771),
.B(n_287),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1878),
.B(n_288),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_1829),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1761),
.B(n_1959),
.Y(n_2327)
);

INVx6_ASAP7_75t_SL g2328 ( 
.A(n_1739),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_1772),
.B(n_289),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_SL g2330 ( 
.A(n_1790),
.B(n_290),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_1888),
.B(n_290),
.Y(n_2331)
);

INVx6_ASAP7_75t_L g2332 ( 
.A(n_1830),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_1691),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1863),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1798),
.B(n_291),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_1798),
.B(n_291),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1825),
.Y(n_2337)
);

BUFx8_ASAP7_75t_L g2338 ( 
.A(n_1874),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1956),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1666),
.Y(n_2340)
);

HB1xp67_ASAP7_75t_L g2341 ( 
.A(n_1803),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_1919),
.B(n_292),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_1783),
.B(n_292),
.Y(n_2343)
);

OR2x6_ASAP7_75t_L g2344 ( 
.A(n_1653),
.B(n_293),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1666),
.Y(n_2345)
);

NAND2x1p5_ASAP7_75t_L g2346 ( 
.A(n_1830),
.B(n_294),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1668),
.Y(n_2347)
);

CKINVDCx20_ASAP7_75t_R g2348 ( 
.A(n_1874),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_1825),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1668),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1863),
.Y(n_2351)
);

OR2x6_ASAP7_75t_L g2352 ( 
.A(n_1664),
.B(n_295),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_1784),
.B(n_1800),
.Y(n_2353)
);

NOR2x1_ASAP7_75t_L g2354 ( 
.A(n_1892),
.B(n_296),
.Y(n_2354)
);

BUFx2_ASAP7_75t_SL g2355 ( 
.A(n_1693),
.Y(n_2355)
);

AND2x6_ASAP7_75t_L g2356 ( 
.A(n_1892),
.B(n_297),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_1807),
.B(n_1808),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_1888),
.B(n_1894),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1857),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_1857),
.Y(n_2360)
);

OR2x6_ASAP7_75t_L g2361 ( 
.A(n_1672),
.B(n_297),
.Y(n_2361)
);

BUFx8_ASAP7_75t_SL g2362 ( 
.A(n_1930),
.Y(n_2362)
);

AND2x6_ASAP7_75t_L g2363 ( 
.A(n_1873),
.B(n_298),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_1857),
.Y(n_2364)
);

INVx4_ASAP7_75t_L g2365 ( 
.A(n_1693),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_1805),
.B(n_298),
.Y(n_2366)
);

INVx5_ASAP7_75t_L g2367 ( 
.A(n_1693),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1670),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_1877),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1894),
.B(n_300),
.Y(n_2370)
);

AND2x4_ASAP7_75t_L g2371 ( 
.A(n_1815),
.B(n_301),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_1825),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_1825),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_1877),
.B(n_301),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_1834),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1670),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1886),
.B(n_302),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1897),
.B(n_304),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1908),
.B(n_305),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1881),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_1799),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_1930),
.B(n_305),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1908),
.B(n_306),
.Y(n_2383)
);

BUFx12f_ASAP7_75t_L g2384 ( 
.A(n_1930),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_1752),
.B(n_307),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_1758),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_1911),
.B(n_308),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_1752),
.B(n_308),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1673),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_1762),
.B(n_309),
.Y(n_2390)
);

AND2x4_ASAP7_75t_L g2391 ( 
.A(n_1823),
.B(n_309),
.Y(n_2391)
);

NAND2x1_ASAP7_75t_L g2392 ( 
.A(n_1707),
.B(n_481),
.Y(n_2392)
);

AND2x2_ASAP7_75t_SL g2393 ( 
.A(n_1873),
.B(n_310),
.Y(n_2393)
);

INVx8_ASAP7_75t_L g2394 ( 
.A(n_1978),
.Y(n_2394)
);

CKINVDCx20_ASAP7_75t_R g2395 ( 
.A(n_2027),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2148),
.Y(n_2396)
);

BUFx2_ASAP7_75t_L g2397 ( 
.A(n_2272),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2293),
.B(n_1921),
.Y(n_2398)
);

INVx4_ASAP7_75t_L g2399 ( 
.A(n_1998),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2013),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2148),
.Y(n_2401)
);

BUFx2_ASAP7_75t_L g2402 ( 
.A(n_2272),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_1998),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2055),
.Y(n_2404)
);

NAND2x1p5_ASAP7_75t_L g2405 ( 
.A(n_2125),
.B(n_1758),
.Y(n_2405)
);

INVx8_ASAP7_75t_L g2406 ( 
.A(n_1978),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_1992),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2293),
.B(n_1921),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2149),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1981),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_1997),
.Y(n_2411)
);

INVx8_ASAP7_75t_L g2412 ( 
.A(n_1992),
.Y(n_2412)
);

BUFx3_ASAP7_75t_L g2413 ( 
.A(n_2026),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2046),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_1981),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_1985),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_SL g2417 ( 
.A(n_2065),
.Y(n_2417)
);

BUFx12f_ASAP7_75t_L g2418 ( 
.A(n_2043),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_1980),
.B(n_1834),
.Y(n_2419)
);

BUFx3_ASAP7_75t_L g2420 ( 
.A(n_2091),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1986),
.B(n_1804),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_1980),
.B(n_1841),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2149),
.Y(n_2423)
);

BUFx12f_ASAP7_75t_L g2424 ( 
.A(n_2016),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2075),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_2140),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2075),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2140),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_2135),
.Y(n_2429)
);

INVx4_ASAP7_75t_L g2430 ( 
.A(n_2125),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2254),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2039),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_1985),
.Y(n_2433)
);

CKINVDCx6p67_ASAP7_75t_R g2434 ( 
.A(n_2065),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2006),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2075),
.Y(n_2436)
);

INVx2_ASAP7_75t_SL g2437 ( 
.A(n_2141),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_2141),
.Y(n_2438)
);

BUFx12f_ASAP7_75t_L g2439 ( 
.A(n_1976),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2254),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2262),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2327),
.B(n_1841),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2301),
.B(n_2309),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_2267),
.Y(n_2444)
);

INVx3_ASAP7_75t_L g2445 ( 
.A(n_2046),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2039),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2123),
.Y(n_2447)
);

CKINVDCx11_ASAP7_75t_R g2448 ( 
.A(n_2115),
.Y(n_2448)
);

BUFx12f_ASAP7_75t_L g2449 ( 
.A(n_2108),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2047),
.Y(n_2450)
);

INVxp67_ASAP7_75t_L g2451 ( 
.A(n_2033),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2046),
.Y(n_2452)
);

BUFx2_ASAP7_75t_L g2453 ( 
.A(n_2142),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2047),
.Y(n_2454)
);

BUFx12f_ASAP7_75t_L g2455 ( 
.A(n_2152),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2006),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2142),
.A2(n_1934),
.B1(n_1935),
.B2(n_1911),
.Y(n_2457)
);

BUFx2_ASAP7_75t_SL g2458 ( 
.A(n_2273),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2291),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2223),
.Y(n_2460)
);

INVxp67_ASAP7_75t_SL g2461 ( 
.A(n_2052),
.Y(n_2461)
);

BUFx12f_ASAP7_75t_L g2462 ( 
.A(n_2115),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2223),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2317),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2068),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2229),
.Y(n_2466)
);

BUFx12f_ASAP7_75t_L g2467 ( 
.A(n_2178),
.Y(n_2467)
);

CKINVDCx16_ASAP7_75t_R g2468 ( 
.A(n_2119),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2099),
.Y(n_2469)
);

BUFx6f_ASAP7_75t_L g2470 ( 
.A(n_2123),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2070),
.Y(n_2471)
);

AO21x1_ASAP7_75t_L g2472 ( 
.A1(n_2052),
.A2(n_2126),
.B(n_2104),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2229),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_2321),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2160),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_2123),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2139),
.Y(n_2477)
);

INVx5_ASAP7_75t_L g2478 ( 
.A(n_2037),
.Y(n_2478)
);

INVx5_ASAP7_75t_SL g2479 ( 
.A(n_2319),
.Y(n_2479)
);

INVx5_ASAP7_75t_L g2480 ( 
.A(n_2037),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2124),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2024),
.Y(n_2482)
);

BUFx12f_ASAP7_75t_L g2483 ( 
.A(n_2178),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2024),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2070),
.Y(n_2485)
);

BUFx4_ASAP7_75t_SL g2486 ( 
.A(n_2181),
.Y(n_2486)
);

INVx8_ASAP7_75t_L g2487 ( 
.A(n_2273),
.Y(n_2487)
);

CKINVDCx6p67_ASAP7_75t_R g2488 ( 
.A(n_2119),
.Y(n_2488)
);

INVx2_ASAP7_75t_SL g2489 ( 
.A(n_2209),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2160),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2131),
.Y(n_2491)
);

NAND2x1p5_ASAP7_75t_L g2492 ( 
.A(n_2222),
.B(n_2236),
.Y(n_2492)
);

INVx6_ASAP7_75t_SL g2493 ( 
.A(n_2238),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2139),
.Y(n_2494)
);

NAND2x1p5_ASAP7_75t_L g2495 ( 
.A(n_2222),
.B(n_1766),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2139),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2365),
.B(n_1673),
.Y(n_2497)
);

INVx1_ASAP7_75t_SL g2498 ( 
.A(n_2068),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2308),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2267),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2145),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2348),
.A2(n_1914),
.B1(n_1893),
.B2(n_1904),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2219),
.A2(n_1914),
.B1(n_1816),
.B2(n_1904),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2029),
.Y(n_2504)
);

INVx1_ASAP7_75t_SL g2505 ( 
.A(n_2069),
.Y(n_2505)
);

CKINVDCx20_ASAP7_75t_R g2506 ( 
.A(n_2170),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2145),
.Y(n_2507)
);

BUFx3_ASAP7_75t_L g2508 ( 
.A(n_1988),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2301),
.B(n_1911),
.Y(n_2509)
);

BUFx8_ASAP7_75t_L g2510 ( 
.A(n_2005),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2314),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2069),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2237),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2338),
.Y(n_2514)
);

BUFx2_ASAP7_75t_L g2515 ( 
.A(n_2338),
.Y(n_2515)
);

BUFx3_ASAP7_75t_L g2516 ( 
.A(n_2362),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2384),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2077),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2071),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2077),
.Y(n_2520)
);

BUFx4f_ASAP7_75t_L g2521 ( 
.A(n_2156),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2145),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2079),
.Y(n_2523)
);

INVxp67_ASAP7_75t_L g2524 ( 
.A(n_2184),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2079),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2146),
.Y(n_2526)
);

NAND2x1p5_ASAP7_75t_L g2527 ( 
.A(n_2236),
.B(n_1766),
.Y(n_2527)
);

BUFx8_ASAP7_75t_L g2528 ( 
.A(n_2005),
.Y(n_2528)
);

BUFx8_ASAP7_75t_L g2529 ( 
.A(n_2008),
.Y(n_2529)
);

INVx5_ASAP7_75t_L g2530 ( 
.A(n_2037),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2168),
.Y(n_2531)
);

HB1xp67_ASAP7_75t_L g2532 ( 
.A(n_2283),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2189),
.Y(n_2533)
);

AND2x6_ASAP7_75t_L g2534 ( 
.A(n_2251),
.B(n_1873),
.Y(n_2534)
);

BUFx12f_ASAP7_75t_L g2535 ( 
.A(n_2218),
.Y(n_2535)
);

OR2x6_ASAP7_75t_L g2536 ( 
.A(n_2156),
.B(n_1873),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2137),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2168),
.Y(n_2538)
);

BUFx2_ASAP7_75t_SL g2539 ( 
.A(n_2008),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2071),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2128),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2251),
.Y(n_2542)
);

INVx5_ASAP7_75t_L g2543 ( 
.A(n_2037),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2082),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2172),
.Y(n_2545)
);

BUFx2_ASAP7_75t_SL g2546 ( 
.A(n_2323),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2309),
.B(n_1934),
.Y(n_2547)
);

BUFx2_ASAP7_75t_L g2548 ( 
.A(n_2319),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2100),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2082),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2340),
.B(n_1935),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2172),
.Y(n_2552)
);

BUFx3_ASAP7_75t_L g2553 ( 
.A(n_2122),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_1973),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2128),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2375),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2246),
.A2(n_1893),
.B1(n_1831),
.B2(n_1833),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2182),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2146),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_2187),
.Y(n_2560)
);

AO22x2_ASAP7_75t_L g2561 ( 
.A1(n_2355),
.A2(n_1754),
.B1(n_1833),
.B2(n_1831),
.Y(n_2561)
);

OR2x6_ASAP7_75t_L g2562 ( 
.A(n_2180),
.B(n_1704),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2182),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1983),
.Y(n_2564)
);

BUFx2_ASAP7_75t_SL g2565 ( 
.A(n_2323),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2210),
.Y(n_2566)
);

BUFx4_ASAP7_75t_SL g2567 ( 
.A(n_2180),
.Y(n_2567)
);

INVxp67_ASAP7_75t_SL g2568 ( 
.A(n_2251),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2283),
.Y(n_2569)
);

BUFx12f_ASAP7_75t_L g2570 ( 
.A(n_2144),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2332),
.Y(n_2571)
);

BUFx12f_ASAP7_75t_L g2572 ( 
.A(n_2144),
.Y(n_2572)
);

INVx3_ASAP7_75t_SL g2573 ( 
.A(n_2191),
.Y(n_2573)
);

INVx5_ASAP7_75t_L g2574 ( 
.A(n_2323),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2332),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2210),
.Y(n_2576)
);

OR2x6_ASAP7_75t_L g2577 ( 
.A(n_2191),
.B(n_1704),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2274),
.B(n_1811),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_1989),
.Y(n_2579)
);

BUFx12f_ASAP7_75t_L g2580 ( 
.A(n_2238),
.Y(n_2580)
);

INVx6_ASAP7_75t_SL g2581 ( 
.A(n_2239),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_1991),
.Y(n_2582)
);

INVx3_ASAP7_75t_SL g2583 ( 
.A(n_2277),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_1999),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2030),
.Y(n_2585)
);

INVx1_ASAP7_75t_SL g2586 ( 
.A(n_2299),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2227),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2018),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2056),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2227),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2019),
.Y(n_2591)
);

CKINVDCx16_ASAP7_75t_R g2592 ( 
.A(n_2151),
.Y(n_2592)
);

BUFx3_ASAP7_75t_L g2593 ( 
.A(n_2048),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2048),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2276),
.B(n_1842),
.Y(n_2595)
);

BUFx3_ASAP7_75t_L g2596 ( 
.A(n_2177),
.Y(n_2596)
);

CKINVDCx16_ASAP7_75t_R g2597 ( 
.A(n_2239),
.Y(n_2597)
);

INVx6_ASAP7_75t_L g2598 ( 
.A(n_2105),
.Y(n_2598)
);

CKINVDCx11_ASAP7_75t_R g2599 ( 
.A(n_2312),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2365),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_2342),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2177),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2086),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2051),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_2367),
.B(n_1778),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2146),
.Y(n_2606)
);

CKINVDCx16_ASAP7_75t_R g2607 ( 
.A(n_2226),
.Y(n_2607)
);

BUFx4f_ASAP7_75t_SL g2608 ( 
.A(n_2363),
.Y(n_2608)
);

NAND2x1p5_ASAP7_75t_L g2609 ( 
.A(n_2367),
.B(n_1778),
.Y(n_2609)
);

INVx5_ASAP7_75t_L g2610 ( 
.A(n_2323),
.Y(n_2610)
);

CKINVDCx20_ASAP7_75t_R g2611 ( 
.A(n_2226),
.Y(n_2611)
);

BUFx2_ASAP7_75t_SL g2612 ( 
.A(n_2363),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2342),
.Y(n_2613)
);

INVx5_ASAP7_75t_L g2614 ( 
.A(n_2363),
.Y(n_2614)
);

BUFx2_ASAP7_75t_L g2615 ( 
.A(n_2356),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2190),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2356),
.Y(n_2617)
);

BUFx4_ASAP7_75t_SL g2618 ( 
.A(n_2312),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_2105),
.Y(n_2619)
);

INVx3_ASAP7_75t_SL g2620 ( 
.A(n_2393),
.Y(n_2620)
);

INVx6_ASAP7_75t_L g2621 ( 
.A(n_2051),
.Y(n_2621)
);

INVx3_ASAP7_75t_L g2622 ( 
.A(n_2177),
.Y(n_2622)
);

INVx6_ASAP7_75t_L g2623 ( 
.A(n_2051),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2183),
.Y(n_2624)
);

INVx6_ASAP7_75t_L g2625 ( 
.A(n_2183),
.Y(n_2625)
);

INVx1_ASAP7_75t_SL g2626 ( 
.A(n_2204),
.Y(n_2626)
);

INVxp67_ASAP7_75t_SL g2627 ( 
.A(n_2212),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_1979),
.Y(n_2628)
);

INVx1_ASAP7_75t_SL g2629 ( 
.A(n_2280),
.Y(n_2629)
);

INVx1_ASAP7_75t_SL g2630 ( 
.A(n_2326),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2183),
.Y(n_2631)
);

BUFx3_ASAP7_75t_L g2632 ( 
.A(n_2040),
.Y(n_2632)
);

BUFx3_ASAP7_75t_L g2633 ( 
.A(n_2040),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_2031),
.Y(n_2634)
);

BUFx12f_ASAP7_75t_L g2635 ( 
.A(n_2059),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2333),
.Y(n_2636)
);

BUFx2_ASAP7_75t_L g2637 ( 
.A(n_2356),
.Y(n_2637)
);

INVx1_ASAP7_75t_SL g2638 ( 
.A(n_2175),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2175),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2114),
.Y(n_2640)
);

BUFx3_ASAP7_75t_L g2641 ( 
.A(n_2116),
.Y(n_2641)
);

NAND2x1p5_ASAP7_75t_L g2642 ( 
.A(n_2367),
.B(n_1782),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2247),
.Y(n_2643)
);

INVx4_ASAP7_75t_L g2644 ( 
.A(n_2356),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2114),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2340),
.B(n_1726),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_2095),
.Y(n_2647)
);

INVx3_ASAP7_75t_SL g2648 ( 
.A(n_2063),
.Y(n_2648)
);

BUFx3_ASAP7_75t_L g2649 ( 
.A(n_2247),
.Y(n_2649)
);

BUFx12f_ASAP7_75t_L g2650 ( 
.A(n_2264),
.Y(n_2650)
);

INVx4_ASAP7_75t_L g2651 ( 
.A(n_2363),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2328),
.Y(n_2652)
);

BUFx12f_ASAP7_75t_L g2653 ( 
.A(n_2109),
.Y(n_2653)
);

BUFx12f_ASAP7_75t_L g2654 ( 
.A(n_2257),
.Y(n_2654)
);

INVx6_ASAP7_75t_SL g2655 ( 
.A(n_2255),
.Y(n_2655)
);

BUFx2_ASAP7_75t_L g2656 ( 
.A(n_2176),
.Y(n_2656)
);

BUFx3_ASAP7_75t_L g2657 ( 
.A(n_2255),
.Y(n_2657)
);

INVxp33_ASAP7_75t_L g2658 ( 
.A(n_1995),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2333),
.Y(n_2659)
);

NAND2x1p5_ASAP7_75t_L g2660 ( 
.A(n_2120),
.B(n_1782),
.Y(n_2660)
);

NAND2x1p5_ASAP7_75t_L g2661 ( 
.A(n_2120),
.B(n_1786),
.Y(n_2661)
);

INVx5_ASAP7_75t_L g2662 ( 
.A(n_1979),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2112),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2049),
.B(n_1842),
.Y(n_2664)
);

INVx6_ASAP7_75t_L g2665 ( 
.A(n_2133),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2057),
.B(n_2203),
.Y(n_2666)
);

BUFx4f_ASAP7_75t_SL g2667 ( 
.A(n_2328),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2285),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2261),
.Y(n_2669)
);

BUFx3_ASAP7_75t_L g2670 ( 
.A(n_2261),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2198),
.B(n_1858),
.Y(n_2671)
);

INVx1_ASAP7_75t_SL g2672 ( 
.A(n_2205),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_1979),
.Y(n_2673)
);

INVx1_ASAP7_75t_SL g2674 ( 
.A(n_2205),
.Y(n_2674)
);

BUFx5_ASAP7_75t_L g2675 ( 
.A(n_1994),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2268),
.Y(n_2676)
);

BUFx12f_ASAP7_75t_L g2677 ( 
.A(n_2092),
.Y(n_2677)
);

INVx5_ASAP7_75t_L g2678 ( 
.A(n_1990),
.Y(n_2678)
);

BUFx12f_ASAP7_75t_L g2679 ( 
.A(n_2199),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2235),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2235),
.Y(n_2681)
);

INVx1_ASAP7_75t_SL g2682 ( 
.A(n_2241),
.Y(n_2682)
);

BUFx12f_ASAP7_75t_L g2683 ( 
.A(n_2282),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2345),
.B(n_1726),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2268),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2241),
.Y(n_2686)
);

INVx5_ASAP7_75t_L g2687 ( 
.A(n_1990),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2216),
.B(n_1847),
.Y(n_2688)
);

BUFx12f_ASAP7_75t_L g2689 ( 
.A(n_2287),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2242),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2278),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2278),
.Y(n_2692)
);

OR2x6_ASAP7_75t_L g2693 ( 
.A(n_2298),
.B(n_1727),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_1990),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2359),
.Y(n_2695)
);

INVx5_ASAP7_75t_L g2696 ( 
.A(n_1994),
.Y(n_2696)
);

BUFx2_ASAP7_75t_SL g2697 ( 
.A(n_2133),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2242),
.Y(n_2698)
);

BUFx2_ASAP7_75t_R g2699 ( 
.A(n_2297),
.Y(n_2699)
);

BUFx4_ASAP7_75t_SL g2700 ( 
.A(n_2344),
.Y(n_2700)
);

CKINVDCx16_ASAP7_75t_R g2701 ( 
.A(n_2004),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2339),
.Y(n_2702)
);

BUFx4_ASAP7_75t_SL g2703 ( 
.A(n_2344),
.Y(n_2703)
);

INVx5_ASAP7_75t_L g2704 ( 
.A(n_1994),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2284),
.Y(n_2705)
);

BUFx3_ASAP7_75t_L g2706 ( 
.A(n_2284),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2286),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2337),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2286),
.Y(n_2709)
);

BUFx3_ASAP7_75t_L g2710 ( 
.A(n_2288),
.Y(n_2710)
);

BUFx12f_ASAP7_75t_L g2711 ( 
.A(n_2346),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2243),
.B(n_1814),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2245),
.Y(n_2713)
);

INVx5_ASAP7_75t_L g2714 ( 
.A(n_1994),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2288),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2080),
.Y(n_2716)
);

INVx3_ASAP7_75t_SL g2717 ( 
.A(n_2303),
.Y(n_2717)
);

NAND2x1p5_ASAP7_75t_L g2718 ( 
.A(n_2080),
.B(n_1786),
.Y(n_2718)
);

INVx5_ASAP7_75t_L g2719 ( 
.A(n_2017),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2303),
.Y(n_2720)
);

CKINVDCx14_ASAP7_75t_R g2721 ( 
.A(n_2009),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2104),
.B(n_1790),
.Y(n_2722)
);

BUFx12f_ASAP7_75t_L g2723 ( 
.A(n_2324),
.Y(n_2723)
);

INVx4_ASAP7_75t_L g2724 ( 
.A(n_2324),
.Y(n_2724)
);

BUFx3_ASAP7_75t_L g2725 ( 
.A(n_2329),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2329),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2343),
.Y(n_2727)
);

BUFx2_ASAP7_75t_L g2728 ( 
.A(n_2058),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2126),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2296),
.B(n_1847),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2359),
.Y(n_2731)
);

INVx4_ASAP7_75t_L g2732 ( 
.A(n_2343),
.Y(n_2732)
);

BUFx3_ASAP7_75t_L g2733 ( 
.A(n_2371),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_2517),
.Y(n_2734)
);

BUFx12f_ASAP7_75t_L g2735 ( 
.A(n_2448),
.Y(n_2735)
);

AOI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2648),
.A2(n_2010),
.B1(n_2369),
.B2(n_2200),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2638),
.Y(n_2737)
);

OAI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2583),
.A2(n_1993),
.B1(n_2015),
.B2(n_2002),
.Y(n_2738)
);

BUFx2_ASAP7_75t_SL g2739 ( 
.A(n_2478),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2486),
.Y(n_2740)
);

BUFx2_ASAP7_75t_L g2741 ( 
.A(n_2510),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2648),
.A2(n_2583),
.B1(n_2521),
.B2(n_2417),
.Y(n_2742)
);

OAI22x1_ASAP7_75t_L g2743 ( 
.A1(n_2620),
.A2(n_2371),
.B1(n_2391),
.B2(n_2110),
.Y(n_2743)
);

INVx6_ASAP7_75t_L g2744 ( 
.A(n_2467),
.Y(n_2744)
);

BUFx2_ASAP7_75t_L g2745 ( 
.A(n_2510),
.Y(n_2745)
);

CKINVDCx20_ASAP7_75t_R g2746 ( 
.A(n_2469),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2521),
.A2(n_2001),
.B1(n_2062),
.B2(n_2007),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2460),
.Y(n_2748)
);

AOI22xp33_ASAP7_75t_SL g2749 ( 
.A1(n_2697),
.A2(n_2138),
.B1(n_2002),
.B2(n_2015),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_SL g2750 ( 
.A1(n_2394),
.A2(n_2138),
.B1(n_1993),
.B2(n_2330),
.Y(n_2750)
);

AOI22xp5_ASAP7_75t_L g2751 ( 
.A1(n_2417),
.A2(n_2081),
.B1(n_2244),
.B2(n_2234),
.Y(n_2751)
);

INVx8_ASAP7_75t_L g2752 ( 
.A(n_2483),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2638),
.Y(n_2753)
);

INVx2_ASAP7_75t_SL g2754 ( 
.A(n_2486),
.Y(n_2754)
);

BUFx2_ASAP7_75t_R g2755 ( 
.A(n_2429),
.Y(n_2755)
);

BUFx10_ASAP7_75t_L g2756 ( 
.A(n_2404),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2620),
.A2(n_2352),
.B1(n_2361),
.B2(n_2316),
.Y(n_2757)
);

INVx2_ASAP7_75t_SL g2758 ( 
.A(n_2487),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2463),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2448),
.A2(n_2361),
.B1(n_2352),
.B2(n_2253),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2466),
.Y(n_2761)
);

CKINVDCx11_ASAP7_75t_R g2762 ( 
.A(n_2395),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2639),
.Y(n_2763)
);

CKINVDCx6p67_ASAP7_75t_R g2764 ( 
.A(n_2599),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2639),
.Y(n_2765)
);

BUFx2_ASAP7_75t_SL g2766 ( 
.A(n_2478),
.Y(n_2766)
);

BUFx2_ASAP7_75t_L g2767 ( 
.A(n_2528),
.Y(n_2767)
);

BUFx10_ASAP7_75t_L g2768 ( 
.A(n_2513),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2473),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2698),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2666),
.B(n_2085),
.Y(n_2771)
);

OAI22xp5_ASAP7_75t_SL g2772 ( 
.A1(n_2597),
.A2(n_2391),
.B1(n_2078),
.B2(n_2073),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2599),
.A2(n_2503),
.B1(n_2406),
.B2(n_2412),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2672),
.Y(n_2774)
);

BUFx8_ASAP7_75t_L g2775 ( 
.A(n_2462),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2503),
.A2(n_2213),
.B1(n_2300),
.B2(n_2093),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2698),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2644),
.Y(n_2778)
);

INVx6_ASAP7_75t_L g2779 ( 
.A(n_2528),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2399),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2672),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2482),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_SL g2783 ( 
.A1(n_2394),
.A2(n_2248),
.B1(n_2292),
.B2(n_2230),
.Y(n_2783)
);

INVx6_ASAP7_75t_L g2784 ( 
.A(n_2529),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2394),
.A2(n_2113),
.B1(n_2096),
.B2(n_2067),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2406),
.A2(n_2412),
.B1(n_2572),
.B2(n_2570),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2674),
.Y(n_2787)
);

BUFx2_ASAP7_75t_SL g2788 ( 
.A(n_2478),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_SL g2789 ( 
.A1(n_2406),
.A2(n_2412),
.B1(n_2592),
.B2(n_2539),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2442),
.B(n_2012),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_SL g2791 ( 
.A1(n_2721),
.A2(n_2529),
.B1(n_2431),
.B2(n_2444),
.Y(n_2791)
);

CKINVDCx6p67_ASAP7_75t_R g2792 ( 
.A(n_2580),
.Y(n_2792)
);

OAI21xp5_ASAP7_75t_SL g2793 ( 
.A1(n_2721),
.A2(n_2067),
.B(n_2058),
.Y(n_2793)
);

CKINVDCx16_ASAP7_75t_R g2794 ( 
.A(n_2506),
.Y(n_2794)
);

BUFx12f_ASAP7_75t_L g2795 ( 
.A(n_2424),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2484),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_SL g2797 ( 
.A1(n_2431),
.A2(n_2248),
.B1(n_2292),
.B2(n_2230),
.Y(n_2797)
);

INVx6_ASAP7_75t_L g2798 ( 
.A(n_2399),
.Y(n_2798)
);

BUFx4f_ASAP7_75t_L g2799 ( 
.A(n_2434),
.Y(n_2799)
);

AOI22xp33_ASAP7_75t_L g2800 ( 
.A1(n_2493),
.A2(n_2014),
.B1(n_2028),
.B2(n_2186),
.Y(n_2800)
);

CKINVDCx20_ASAP7_75t_R g2801 ( 
.A(n_2395),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2717),
.B(n_1974),
.Y(n_2802)
);

AOI22xp33_ASAP7_75t_L g2803 ( 
.A1(n_2493),
.A2(n_2275),
.B1(n_2358),
.B2(n_2341),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_2619),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2502),
.A2(n_2169),
.B1(n_2127),
.B2(n_2053),
.Y(n_2805)
);

CKINVDCx20_ASAP7_75t_R g2806 ( 
.A(n_2516),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2410),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2660),
.A2(n_2289),
.B1(n_2318),
.B2(n_2307),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2581),
.A2(n_2295),
.B1(n_1996),
.B2(n_2258),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2674),
.Y(n_2810)
);

BUFx12f_ASAP7_75t_L g2811 ( 
.A(n_2418),
.Y(n_2811)
);

CKINVDCx20_ASAP7_75t_R g2812 ( 
.A(n_2560),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2593),
.Y(n_2813)
);

BUFx3_ASAP7_75t_L g2814 ( 
.A(n_2411),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2581),
.A2(n_1975),
.B1(n_1982),
.B2(n_2331),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2562),
.A2(n_2336),
.B1(n_2335),
.B2(n_2374),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_SL g2817 ( 
.A1(n_2440),
.A2(n_2305),
.B1(n_1790),
.B2(n_1707),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2594),
.Y(n_2818)
);

OAI21xp33_ASAP7_75t_L g2819 ( 
.A1(n_2502),
.A2(n_1875),
.B(n_2161),
.Y(n_2819)
);

INVx1_ASAP7_75t_SL g2820 ( 
.A(n_2700),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2415),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2421),
.B(n_2345),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2416),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2562),
.A2(n_2577),
.B1(n_2573),
.B2(n_2557),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2433),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2435),
.Y(n_2826)
);

OAI22xp5_ASAP7_75t_SL g2827 ( 
.A1(n_2573),
.A2(n_2306),
.B1(n_2392),
.B2(n_2233),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2562),
.A2(n_2165),
.B1(n_2064),
.B2(n_2076),
.Y(n_2828)
);

BUFx8_ASAP7_75t_L g2829 ( 
.A(n_2514),
.Y(n_2829)
);

BUFx3_ASAP7_75t_L g2830 ( 
.A(n_2413),
.Y(n_2830)
);

BUFx4_ASAP7_75t_R g2831 ( 
.A(n_2567),
.Y(n_2831)
);

INVx6_ASAP7_75t_L g2832 ( 
.A(n_2455),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2722),
.A2(n_1754),
.B(n_2729),
.Y(n_2833)
);

BUFx4f_ASAP7_75t_SL g2834 ( 
.A(n_2449),
.Y(n_2834)
);

AOI22xp5_ASAP7_75t_L g2835 ( 
.A1(n_2668),
.A2(n_2320),
.B1(n_1987),
.B2(n_2094),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2577),
.A2(n_2054),
.B1(n_2382),
.B2(n_2143),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2660),
.A2(n_2661),
.B1(n_2577),
.B2(n_2717),
.Y(n_2837)
);

INVx6_ASAP7_75t_L g2838 ( 
.A(n_2487),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2456),
.Y(n_2839)
);

BUFx3_ASAP7_75t_L g2840 ( 
.A(n_2481),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2557),
.A2(n_2225),
.B1(n_2097),
.B2(n_1790),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2425),
.Y(n_2842)
);

OAI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2661),
.A2(n_2111),
.B1(n_2060),
.B2(n_2174),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2682),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2471),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2701),
.A2(n_2322),
.B1(n_2350),
.B2(n_2347),
.Y(n_2846)
);

AOI22xp33_ASAP7_75t_L g2847 ( 
.A1(n_2440),
.A2(n_2444),
.B1(n_2500),
.B2(n_2407),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2718),
.A2(n_2192),
.B1(n_2196),
.B2(n_2179),
.Y(n_2848)
);

CKINVDCx8_ASAP7_75t_R g2849 ( 
.A(n_2458),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2682),
.Y(n_2850)
);

AOI22xp33_ASAP7_75t_SL g2851 ( 
.A1(n_2665),
.A2(n_2305),
.B1(n_1790),
.B2(n_1707),
.Y(n_2851)
);

CKINVDCx11_ASAP7_75t_R g2852 ( 
.A(n_2535),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2686),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2611),
.A2(n_1984),
.B1(n_2366),
.B2(n_2207),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2630),
.B(n_2302),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2686),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2718),
.A2(n_2084),
.B1(n_2090),
.B2(n_2379),
.Y(n_2857)
);

INVx4_ASAP7_75t_L g2858 ( 
.A(n_2608),
.Y(n_2858)
);

CKINVDCx20_ASAP7_75t_R g2859 ( 
.A(n_2611),
.Y(n_2859)
);

OAI22x1_ASAP7_75t_L g2860 ( 
.A1(n_2601),
.A2(n_2613),
.B1(n_2451),
.B2(n_2515),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2485),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2425),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2693),
.A2(n_2011),
.B1(n_2003),
.B2(n_2385),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2519),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2540),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2693),
.A2(n_2350),
.B1(n_2368),
.B2(n_2347),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2693),
.A2(n_2376),
.B1(n_2389),
.B2(n_2368),
.Y(n_2867)
);

AOI22xp33_ASAP7_75t_L g2868 ( 
.A1(n_2658),
.A2(n_2389),
.B1(n_2376),
.B2(n_2202),
.Y(n_2868)
);

BUFx2_ASAP7_75t_L g2869 ( 
.A(n_2655),
.Y(n_2869)
);

CKINVDCx11_ASAP7_75t_R g2870 ( 
.A(n_2439),
.Y(n_2870)
);

BUFx2_ASAP7_75t_L g2871 ( 
.A(n_2655),
.Y(n_2871)
);

NAND2x1p5_ASAP7_75t_L g2872 ( 
.A(n_2430),
.B(n_2185),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2680),
.Y(n_2873)
);

BUFx8_ASAP7_75t_L g2874 ( 
.A(n_2635),
.Y(n_2874)
);

NAND2x1p5_ASAP7_75t_L g2875 ( 
.A(n_2430),
.B(n_2185),
.Y(n_2875)
);

CKINVDCx11_ASAP7_75t_R g2876 ( 
.A(n_2420),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2681),
.Y(n_2877)
);

BUFx2_ASAP7_75t_L g2878 ( 
.A(n_2679),
.Y(n_2878)
);

INVx6_ASAP7_75t_L g2879 ( 
.A(n_2487),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_2425),
.Y(n_2880)
);

INVx5_ASAP7_75t_SL g2881 ( 
.A(n_2536),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2690),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2713),
.Y(n_2883)
);

BUFx12f_ASAP7_75t_L g2884 ( 
.A(n_2441),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2544),
.Y(n_2885)
);

INVx4_ASAP7_75t_L g2886 ( 
.A(n_2608),
.Y(n_2886)
);

INVx3_ASAP7_75t_L g2887 ( 
.A(n_2644),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2630),
.B(n_2217),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2550),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2443),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2443),
.Y(n_2891)
);

BUFx8_ASAP7_75t_L g2892 ( 
.A(n_2683),
.Y(n_2892)
);

OAI22x1_ASAP7_75t_L g2893 ( 
.A1(n_2451),
.A2(n_2000),
.B1(n_2354),
.B2(n_2387),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2724),
.B(n_2217),
.Y(n_2894)
);

INVx4_ASAP7_75t_L g2895 ( 
.A(n_2480),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2554),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2421),
.B(n_2270),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2398),
.Y(n_2898)
);

INVx4_ASAP7_75t_L g2899 ( 
.A(n_2480),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2724),
.B(n_2270),
.Y(n_2900)
);

OAI22x1_ASAP7_75t_L g2901 ( 
.A1(n_2618),
.A2(n_2000),
.B1(n_2354),
.B2(n_2387),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2398),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2700),
.Y(n_2903)
);

INVx6_ASAP7_75t_L g2904 ( 
.A(n_2711),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2408),
.Y(n_2905)
);

BUFx2_ASAP7_75t_SL g2906 ( 
.A(n_2480),
.Y(n_2906)
);

AOI22xp33_ASAP7_75t_SL g2907 ( 
.A1(n_2665),
.A2(n_1707),
.B1(n_2313),
.B2(n_2129),
.Y(n_2907)
);

OAI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2479),
.A2(n_2383),
.B1(n_2061),
.B2(n_2232),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2578),
.B(n_2304),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2408),
.Y(n_2910)
);

AOI22xp33_ASAP7_75t_L g2911 ( 
.A1(n_2658),
.A2(n_2201),
.B1(n_1870),
.B2(n_2310),
.Y(n_2911)
);

BUFx4f_ASAP7_75t_SL g2912 ( 
.A(n_2689),
.Y(n_2912)
);

BUFx12f_ASAP7_75t_SL g2913 ( 
.A(n_2618),
.Y(n_2913)
);

BUFx12f_ASAP7_75t_L g2914 ( 
.A(n_2537),
.Y(n_2914)
);

OAI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2479),
.A2(n_2263),
.B1(n_2266),
.B2(n_2231),
.Y(n_2915)
);

OAI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2732),
.A2(n_1972),
.B1(n_2050),
.B2(n_2042),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2564),
.Y(n_2917)
);

CKINVDCx11_ASAP7_75t_R g2918 ( 
.A(n_2533),
.Y(n_2918)
);

OAI22xp33_ASAP7_75t_L g2919 ( 
.A1(n_2732),
.A2(n_2167),
.B1(n_2159),
.B2(n_2279),
.Y(n_2919)
);

AOI22xp33_ASAP7_75t_L g2920 ( 
.A1(n_2723),
.A2(n_1870),
.B1(n_1779),
.B2(n_2206),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2579),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2582),
.Y(n_2922)
);

OAI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_2536),
.A2(n_2294),
.B1(n_2370),
.B2(n_2195),
.Y(n_2923)
);

BUFx2_ASAP7_75t_L g2924 ( 
.A(n_2414),
.Y(n_2924)
);

BUFx12f_ASAP7_75t_L g2925 ( 
.A(n_2652),
.Y(n_2925)
);

OAI21xp33_ASAP7_75t_SL g2926 ( 
.A1(n_2651),
.A2(n_1677),
.B(n_1695),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2584),
.Y(n_2927)
);

CKINVDCx6p67_ASAP7_75t_R g2928 ( 
.A(n_2607),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_SL g2929 ( 
.A1(n_2479),
.A2(n_1707),
.B1(n_1851),
.B2(n_1737),
.Y(n_2929)
);

NAND2x1p5_ASAP7_75t_L g2930 ( 
.A(n_2490),
.B(n_2188),
.Y(n_2930)
);

BUFx10_ASAP7_75t_L g2931 ( 
.A(n_2567),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2491),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2588),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2591),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2671),
.A2(n_2353),
.B1(n_2357),
.B2(n_2304),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_2427),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2603),
.Y(n_2937)
);

INVx8_ASAP7_75t_L g2938 ( 
.A(n_2536),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2663),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2556),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2509),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_2524),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2509),
.Y(n_2943)
);

CKINVDCx11_ASAP7_75t_R g2944 ( 
.A(n_2488),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2531),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2512),
.A2(n_1870),
.B1(n_2215),
.B2(n_2214),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2547),
.Y(n_2947)
);

INVx4_ASAP7_75t_L g2948 ( 
.A(n_2530),
.Y(n_2948)
);

AOI22xp33_ASAP7_75t_SL g2949 ( 
.A1(n_2649),
.A2(n_1849),
.B1(n_1677),
.B2(n_2102),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_L g2950 ( 
.A(n_2427),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2547),
.Y(n_2951)
);

BUFx6f_ASAP7_75t_SL g2952 ( 
.A(n_2703),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_SL g2953 ( 
.A1(n_2657),
.A2(n_2154),
.B1(n_2155),
.B2(n_2106),
.Y(n_2953)
);

BUFx4f_ASAP7_75t_SL g2954 ( 
.A(n_2400),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_SL g2955 ( 
.A1(n_2670),
.A2(n_2158),
.B1(n_2157),
.B2(n_2224),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2512),
.A2(n_1732),
.B1(n_1738),
.B2(n_1725),
.Y(n_2956)
);

BUFx4f_ASAP7_75t_SL g2957 ( 
.A(n_2571),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2728),
.A2(n_1753),
.B1(n_2083),
.B2(n_1923),
.Y(n_2958)
);

CKINVDCx20_ASAP7_75t_R g2959 ( 
.A(n_2667),
.Y(n_2959)
);

INVx6_ASAP7_75t_L g2960 ( 
.A(n_2604),
.Y(n_2960)
);

OAI22x1_ASAP7_75t_L g2961 ( 
.A1(n_2548),
.A2(n_2357),
.B1(n_2353),
.B2(n_2117),
.Y(n_2961)
);

OAI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2426),
.A2(n_2388),
.B1(n_2023),
.B2(n_1926),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2538),
.Y(n_2963)
);

INVx1_ASAP7_75t_SL g2964 ( 
.A(n_2703),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_SL g2965 ( 
.A1(n_2685),
.A2(n_2121),
.B1(n_2130),
.B2(n_2118),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2545),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2552),
.Y(n_2967)
);

OAI22xp33_ASAP7_75t_L g2968 ( 
.A1(n_2426),
.A2(n_2377),
.B1(n_2378),
.B2(n_2325),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2428),
.A2(n_2498),
.B1(n_2505),
.B2(n_2465),
.Y(n_2969)
);

NAND2x1p5_ASAP7_75t_L g2970 ( 
.A(n_2490),
.B(n_2188),
.Y(n_2970)
);

INVx6_ASAP7_75t_L g2971 ( 
.A(n_2604),
.Y(n_2971)
);

AOI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_2677),
.A2(n_1925),
.B1(n_1880),
.B2(n_1901),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2551),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2650),
.A2(n_1917),
.B1(n_1905),
.B2(n_1788),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_SL g2975 ( 
.A1(n_2692),
.A2(n_2121),
.B1(n_2130),
.B2(n_2118),
.Y(n_2975)
);

CKINVDCx20_ASAP7_75t_R g2976 ( 
.A(n_2667),
.Y(n_2976)
);

INVx6_ASAP7_75t_L g2977 ( 
.A(n_2621),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2819),
.A2(n_2653),
.B1(n_2716),
.B2(n_2710),
.Y(n_2978)
);

OAI222xp33_ASAP7_75t_L g2979 ( 
.A1(n_2750),
.A2(n_2505),
.B1(n_2465),
.B2(n_2498),
.C1(n_2428),
.C2(n_2651),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2813),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2748),
.Y(n_2981)
);

INVx5_ASAP7_75t_SL g2982 ( 
.A(n_2764),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2771),
.B(n_2524),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2790),
.B(n_2589),
.Y(n_2984)
);

AOI222xp33_ASAP7_75t_L g2985 ( 
.A1(n_2952),
.A2(n_2772),
.B1(n_2854),
.B2(n_2793),
.C1(n_2799),
.C2(n_2964),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2888),
.B(n_2706),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2812),
.B(n_2654),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2736),
.A2(n_2725),
.B1(n_2733),
.B2(n_2715),
.Y(n_2988)
);

AOI222xp33_ASAP7_75t_L g2989 ( 
.A1(n_2952),
.A2(n_2656),
.B1(n_2671),
.B2(n_2454),
.C1(n_2432),
.C2(n_2450),
.Y(n_2989)
);

AOI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2846),
.A2(n_2640),
.B1(n_2645),
.B2(n_2446),
.Y(n_2990)
);

OAI21xp33_ASAP7_75t_L g2991 ( 
.A1(n_2972),
.A2(n_2561),
.B(n_2699),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2759),
.Y(n_2992)
);

CKINVDCx11_ASAP7_75t_R g2993 ( 
.A(n_2931),
.Y(n_2993)
);

BUFx6f_ASAP7_75t_L g2994 ( 
.A(n_2813),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2783),
.A2(n_2617),
.B1(n_2637),
.B2(n_2615),
.Y(n_2995)
);

AOI22xp33_ASAP7_75t_L g2996 ( 
.A1(n_2919),
.A2(n_2497),
.B1(n_2563),
.B2(n_2558),
.Y(n_2996)
);

AOI22xp33_ASAP7_75t_L g2997 ( 
.A1(n_2955),
.A2(n_2497),
.B1(n_2576),
.B2(n_2566),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2890),
.B(n_2587),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2761),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2824),
.A2(n_2643),
.B1(n_2669),
.B2(n_2590),
.Y(n_3000)
);

INVx3_ASAP7_75t_L g3001 ( 
.A(n_2780),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2953),
.A2(n_2691),
.B1(n_2705),
.B2(n_2676),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2769),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_SL g3004 ( 
.A1(n_2938),
.A2(n_2565),
.B1(n_2612),
.B2(n_2546),
.Y(n_3004)
);

OAI22xp5_ASAP7_75t_L g3005 ( 
.A1(n_2749),
.A2(n_2543),
.B1(n_2574),
.B2(n_2530),
.Y(n_3005)
);

OAI21xp33_ASAP7_75t_L g3006 ( 
.A1(n_2760),
.A2(n_2561),
.B(n_2699),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2891),
.B(n_2707),
.Y(n_3007)
);

BUFx3_ASAP7_75t_L g3008 ( 
.A(n_2734),
.Y(n_3008)
);

AOI22xp33_ASAP7_75t_L g3009 ( 
.A1(n_2776),
.A2(n_2720),
.B1(n_2726),
.B2(n_2709),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2855),
.B(n_2595),
.Y(n_3010)
);

INVx2_ASAP7_75t_SL g3011 ( 
.A(n_2892),
.Y(n_3011)
);

OAI21xp33_ASAP7_75t_L g3012 ( 
.A1(n_2974),
.A2(n_2712),
.B(n_2634),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2813),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2778),
.B(n_2530),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2892),
.Y(n_3015)
);

OAI22xp33_ASAP7_75t_L g3016 ( 
.A1(n_2935),
.A2(n_2468),
.B1(n_2574),
.B2(n_2543),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2909),
.B(n_2727),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2913),
.A2(n_2511),
.B1(n_2499),
.B2(n_2647),
.Y(n_3018)
);

INVx4_ASAP7_75t_L g3019 ( 
.A(n_2831),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2924),
.Y(n_3020)
);

BUFx4f_ASAP7_75t_SL g3021 ( 
.A(n_2874),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2915),
.A2(n_2730),
.B1(n_2396),
.B2(n_2409),
.Y(n_3022)
);

OAI222xp33_ASAP7_75t_L g3023 ( 
.A1(n_2797),
.A2(n_2610),
.B1(n_2543),
.B2(n_2614),
.C1(n_2574),
.C2(n_2461),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_SL g3024 ( 
.A1(n_2938),
.A2(n_2837),
.B1(n_2610),
.B2(n_2614),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2916),
.A2(n_2423),
.B1(n_2401),
.B2(n_2664),
.Y(n_3025)
);

OAI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2820),
.A2(n_2614),
.B1(n_2610),
.B2(n_2475),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2873),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2782),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2903),
.B(n_2702),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2877),
.Y(n_3030)
);

OAI21xp33_ASAP7_75t_L g3031 ( 
.A1(n_2757),
.A2(n_1694),
.B(n_1692),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2908),
.A2(n_2688),
.B1(n_2518),
.B2(n_2523),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_2773),
.A2(n_2520),
.B1(n_2525),
.B2(n_2461),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2816),
.A2(n_2397),
.B1(n_2402),
.B2(n_2616),
.Y(n_3034)
);

OAI21xp5_ASAP7_75t_SL g3035 ( 
.A1(n_2738),
.A2(n_2453),
.B(n_2405),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2796),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2848),
.A2(n_2616),
.B1(n_2629),
.B2(n_2626),
.Y(n_3037)
);

AOI22xp33_ASAP7_75t_L g3038 ( 
.A1(n_2923),
.A2(n_2815),
.B1(n_2747),
.B2(n_2743),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_SL g3039 ( 
.A1(n_2881),
.A2(n_2729),
.B1(n_2532),
.B2(n_2569),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2807),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2874),
.Y(n_3041)
);

BUFx3_ASAP7_75t_L g3042 ( 
.A(n_2912),
.Y(n_3042)
);

AOI21xp33_ASAP7_75t_L g3043 ( 
.A1(n_2901),
.A2(n_2390),
.B(n_2101),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2751),
.A2(n_2626),
.B1(n_2629),
.B2(n_2457),
.Y(n_3044)
);

AOI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_2843),
.A2(n_2457),
.B1(n_2419),
.B2(n_2422),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2818),
.Y(n_3046)
);

AOI222xp33_ASAP7_75t_L g3047 ( 
.A1(n_2799),
.A2(n_2735),
.B1(n_2897),
.B2(n_2742),
.C1(n_2931),
.C2(n_2741),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2904),
.Y(n_3048)
);

BUFx3_ASAP7_75t_R g3049 ( 
.A(n_2745),
.Y(n_3049)
);

BUFx4f_ASAP7_75t_SL g3050 ( 
.A(n_2795),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2857),
.A2(n_2472),
.B1(n_2627),
.B2(n_2569),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2851),
.A2(n_2532),
.B1(n_2627),
.B2(n_2405),
.Y(n_3052)
);

OAI21xp33_ASAP7_75t_L g3053 ( 
.A1(n_2800),
.A2(n_1699),
.B(n_1802),
.Y(n_3053)
);

AOI22xp33_ASAP7_75t_L g3054 ( 
.A1(n_2841),
.A2(n_2403),
.B1(n_2508),
.B2(n_2586),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2863),
.A2(n_2403),
.B1(n_2586),
.B2(n_1931),
.Y(n_3055)
);

OAI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2785),
.A2(n_2492),
.B1(n_2659),
.B2(n_2636),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2818),
.B(n_2489),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2818),
.B(n_2414),
.Y(n_3058)
);

AOI222xp33_ASAP7_75t_L g3059 ( 
.A1(n_2767),
.A2(n_2646),
.B1(n_2684),
.B2(n_1769),
.C1(n_1883),
.C2(n_1727),
.Y(n_3059)
);

CKINVDCx5p33_ASAP7_75t_R g3060 ( 
.A(n_2762),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2882),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_2803),
.A2(n_1931),
.B1(n_1929),
.B2(n_2646),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2821),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2780),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2836),
.A2(n_2791),
.B1(n_2968),
.B2(n_2828),
.Y(n_3065)
);

OAI22xp5_ASAP7_75t_L g3066 ( 
.A1(n_2817),
.A2(n_2907),
.B1(n_2975),
.B2(n_2965),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2780),
.Y(n_3067)
);

AOI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2929),
.A2(n_2722),
.B(n_1891),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2804),
.B(n_2445),
.Y(n_3069)
);

AOI22xp33_ASAP7_75t_L g3070 ( 
.A1(n_2946),
.A2(n_1929),
.B1(n_2684),
.B2(n_1734),
.Y(n_3070)
);

AOI22xp33_ASAP7_75t_L g3071 ( 
.A1(n_2809),
.A2(n_1734),
.B1(n_2171),
.B2(n_2164),
.Y(n_3071)
);

OAI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2805),
.A2(n_2492),
.B1(n_2600),
.B2(n_2636),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2898),
.B(n_2132),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2947),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2958),
.A2(n_1860),
.B1(n_2162),
.B2(n_2132),
.Y(n_3075)
);

OAI21xp33_ASAP7_75t_L g3076 ( 
.A1(n_2835),
.A2(n_2956),
.B(n_2847),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2904),
.Y(n_3077)
);

INVx4_ASAP7_75t_L g3078 ( 
.A(n_2954),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_2911),
.A2(n_2162),
.B1(n_2163),
.B2(n_2459),
.Y(n_3079)
);

CKINVDCx5p33_ASAP7_75t_R g3080 ( 
.A(n_2876),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_SL g3081 ( 
.A1(n_2881),
.A2(n_2600),
.B1(n_2659),
.B2(n_2445),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2823),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2894),
.B(n_2452),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_2868),
.A2(n_2163),
.B1(n_2464),
.B2(n_2459),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2825),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2866),
.A2(n_2464),
.B1(n_2474),
.B2(n_2098),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2902),
.B(n_2551),
.Y(n_3087)
);

AOI22xp33_ASAP7_75t_L g3088 ( 
.A1(n_2867),
.A2(n_2474),
.B1(n_1846),
.B2(n_1883),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_SL g3089 ( 
.A1(n_2789),
.A2(n_2452),
.B(n_2495),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2905),
.B(n_2910),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2826),
.Y(n_3091)
);

OAI21xp5_ASAP7_75t_SL g3092 ( 
.A1(n_2740),
.A2(n_2527),
.B(n_2495),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2961),
.A2(n_1723),
.B1(n_1891),
.B2(n_2585),
.Y(n_3093)
);

OAI21xp33_ASAP7_75t_L g3094 ( 
.A1(n_2942),
.A2(n_2438),
.B(n_2437),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2962),
.A2(n_2633),
.B1(n_2632),
.B2(n_2193),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_L g3096 ( 
.A1(n_2920),
.A2(n_2527),
.B1(n_2598),
.B2(n_2696),
.Y(n_3096)
);

INVxp67_ASAP7_75t_L g3097 ( 
.A(n_2830),
.Y(n_3097)
);

INVx5_ASAP7_75t_SL g3098 ( 
.A(n_2792),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2839),
.Y(n_3099)
);

OAI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_2798),
.A2(n_2598),
.B1(n_2704),
.B2(n_2696),
.Y(n_3100)
);

BUFx4f_ASAP7_75t_SL g3101 ( 
.A(n_2811),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2928),
.A2(n_2193),
.B1(n_2290),
.B2(n_2220),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2845),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2883),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2798),
.A2(n_2704),
.B1(n_2714),
.B2(n_2696),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2900),
.B(n_2549),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_L g3107 ( 
.A1(n_2779),
.A2(n_2220),
.B1(n_2290),
.B2(n_1926),
.Y(n_3107)
);

INVxp67_ASAP7_75t_SL g3108 ( 
.A(n_2737),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2779),
.A2(n_2250),
.B1(n_2271),
.B2(n_2240),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2802),
.B(n_2553),
.Y(n_3110)
);

HB1xp67_ASAP7_75t_L g3111 ( 
.A(n_2951),
.Y(n_3111)
);

OAI222xp33_ASAP7_75t_L g3112 ( 
.A1(n_2808),
.A2(n_2714),
.B1(n_2704),
.B2(n_2256),
.C1(n_2568),
.C2(n_2542),
.Y(n_3112)
);

AOI22xp33_ASAP7_75t_L g3113 ( 
.A1(n_2784),
.A2(n_2641),
.B1(n_2504),
.B2(n_1646),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2861),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_L g3115 ( 
.A1(n_2784),
.A2(n_2504),
.B1(n_1648),
.B2(n_1960),
.Y(n_3115)
);

OAI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2786),
.A2(n_2714),
.B1(n_2568),
.B2(n_2623),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2943),
.A2(n_2777),
.B1(n_2770),
.B2(n_2822),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2864),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2865),
.Y(n_3119)
);

OAI21xp33_ASAP7_75t_L g3120 ( 
.A1(n_2893),
.A2(n_1869),
.B(n_1907),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2885),
.B(n_2542),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2849),
.A2(n_2623),
.B1(n_2621),
.B2(n_2609),
.Y(n_3122)
);

AOI211xp5_ASAP7_75t_L g3123 ( 
.A1(n_2754),
.A2(n_1951),
.B(n_1965),
.C(n_1639),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2969),
.A2(n_1964),
.B1(n_1968),
.B2(n_1780),
.Y(n_3124)
);

OAI21xp5_ASAP7_75t_SL g3125 ( 
.A1(n_2778),
.A2(n_2609),
.B(n_2605),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2896),
.Y(n_3126)
);

AOI21xp33_ASAP7_75t_L g3127 ( 
.A1(n_2926),
.A2(n_1954),
.B(n_2541),
.Y(n_3127)
);

AOI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2801),
.A2(n_2860),
.B1(n_2878),
.B2(n_2859),
.Y(n_3128)
);

AND2x4_ASAP7_75t_L g3129 ( 
.A(n_2887),
.B(n_2596),
.Y(n_3129)
);

BUFx6f_ASAP7_75t_L g3130 ( 
.A(n_2842),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_2941),
.A2(n_2025),
.B1(n_2035),
.B2(n_2020),
.Y(n_3131)
);

AOI222xp33_ASAP7_75t_L g3132 ( 
.A1(n_2775),
.A2(n_1832),
.B1(n_1719),
.B2(n_1909),
.C1(n_2575),
.C2(n_1954),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2889),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2921),
.Y(n_3134)
);

AOI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_2960),
.A2(n_2197),
.B1(n_2259),
.B2(n_1955),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2922),
.B(n_2245),
.Y(n_3136)
);

OAI21xp5_ASAP7_75t_SL g3137 ( 
.A1(n_2887),
.A2(n_2642),
.B(n_2605),
.Y(n_3137)
);

BUFx2_ASAP7_75t_L g3138 ( 
.A(n_2960),
.Y(n_3138)
);

CKINVDCx14_ASAP7_75t_R g3139 ( 
.A(n_2959),
.Y(n_3139)
);

OAI22xp33_ASAP7_75t_L g3140 ( 
.A1(n_2858),
.A2(n_2642),
.B1(n_2364),
.B2(n_2360),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2927),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2973),
.A2(n_1903),
.B1(n_2381),
.B2(n_2364),
.Y(n_3142)
);

OAI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_2858),
.A2(n_2252),
.B1(n_2249),
.B2(n_2041),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2933),
.B(n_2249),
.Y(n_3144)
);

AOI22xp33_ASAP7_75t_SL g3145 ( 
.A1(n_2739),
.A2(n_2675),
.B1(n_2731),
.B2(n_2695),
.Y(n_3145)
);

OAI22xp33_ASAP7_75t_SL g3146 ( 
.A1(n_2971),
.A2(n_2625),
.B1(n_2731),
.B2(n_2695),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_SL g3147 ( 
.A1(n_2739),
.A2(n_2675),
.B1(n_2534),
.B2(n_2625),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2917),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2829),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2886),
.A2(n_1903),
.B1(n_2381),
.B2(n_2360),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2934),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2985),
.A2(n_2963),
.B1(n_2966),
.B2(n_2945),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_3010),
.B(n_2753),
.Y(n_3153)
);

OAI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_3065),
.A2(n_2886),
.B1(n_2971),
.B2(n_2766),
.Y(n_3154)
);

AOI222xp33_ASAP7_75t_L g3155 ( 
.A1(n_3076),
.A2(n_2829),
.B1(n_2775),
.B2(n_2944),
.C1(n_2967),
.C2(n_2752),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_3074),
.Y(n_3156)
);

AND2x2_ASAP7_75t_SL g3157 ( 
.A(n_3019),
.B(n_3014),
.Y(n_3157)
);

AOI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_2985),
.A2(n_2869),
.B1(n_2871),
.B2(n_2949),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_3019),
.A2(n_2827),
.B1(n_2788),
.B2(n_2766),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_3006),
.A2(n_2906),
.B1(n_2788),
.B2(n_2937),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2981),
.Y(n_3161)
);

OAI222xp33_ASAP7_75t_L g3162 ( 
.A1(n_3038),
.A2(n_2899),
.B1(n_2895),
.B2(n_2948),
.C1(n_2794),
.C2(n_2850),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2991),
.A2(n_2906),
.B1(n_2895),
.B2(n_2899),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_3053),
.A2(n_2948),
.B1(n_1903),
.B2(n_2977),
.Y(n_3164)
);

OAI221xp5_ASAP7_75t_SL g3165 ( 
.A1(n_2997),
.A2(n_2758),
.B1(n_2840),
.B2(n_2940),
.C(n_2932),
.Y(n_3165)
);

AOI22xp33_ASAP7_75t_L g3166 ( 
.A1(n_3066),
.A2(n_1903),
.B1(n_2977),
.B2(n_2939),
.Y(n_3166)
);

OR2x2_ASAP7_75t_L g3167 ( 
.A(n_3111),
.B(n_2763),
.Y(n_3167)
);

OAI22xp5_ASAP7_75t_L g3168 ( 
.A1(n_2996),
.A2(n_2838),
.B1(n_2879),
.B2(n_2875),
.Y(n_3168)
);

AOI22xp33_ASAP7_75t_L g3169 ( 
.A1(n_3031),
.A2(n_2774),
.B1(n_2781),
.B2(n_2765),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2992),
.Y(n_3170)
);

OA222x2_ASAP7_75t_L g3171 ( 
.A1(n_3049),
.A2(n_2814),
.B1(n_2810),
.B2(n_2856),
.C1(n_2844),
.C2(n_2853),
.Y(n_3171)
);

BUFx2_ASAP7_75t_L g3172 ( 
.A(n_2980),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2999),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3040),
.B(n_2787),
.Y(n_3174)
);

OAI22xp5_ASAP7_75t_L g3175 ( 
.A1(n_3025),
.A2(n_3092),
.B1(n_3002),
.B2(n_3045),
.Y(n_3175)
);

OAI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3092),
.A2(n_2838),
.B1(n_2879),
.B2(n_2872),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_3132),
.A2(n_1932),
.B1(n_1941),
.B2(n_1940),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_SL g3178 ( 
.A1(n_2995),
.A2(n_3052),
.B1(n_3021),
.B2(n_3020),
.Y(n_3178)
);

AOI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_3059),
.A2(n_2744),
.B1(n_2832),
.B2(n_1955),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_3043),
.A2(n_1939),
.B(n_2930),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3012),
.A2(n_2744),
.B1(n_2832),
.B2(n_2806),
.Y(n_3181)
);

AOI22xp33_ASAP7_75t_SL g3182 ( 
.A1(n_3020),
.A2(n_2752),
.B1(n_2834),
.B2(n_2976),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_L g3183 ( 
.A1(n_2983),
.A2(n_1944),
.B1(n_2534),
.B2(n_1927),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_3032),
.A2(n_2534),
.B1(n_1927),
.B2(n_2602),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_L g3185 ( 
.A1(n_3022),
.A2(n_2534),
.B1(n_2044),
.B2(n_2045),
.Y(n_3185)
);

AOI22xp5_ASAP7_75t_L g3186 ( 
.A1(n_2990),
.A2(n_2022),
.B1(n_2089),
.B2(n_1977),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2984),
.A2(n_2066),
.B1(n_2269),
.B2(n_2036),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3000),
.A2(n_2173),
.B1(n_2072),
.B2(n_2970),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_3033),
.A2(n_2311),
.B1(n_2315),
.B2(n_2281),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3110),
.B(n_2622),
.Y(n_3190)
);

INVxp67_ASAP7_75t_SL g3191 ( 
.A(n_3108),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3063),
.B(n_2252),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_L g3193 ( 
.A1(n_3047),
.A2(n_2351),
.B1(n_2380),
.B2(n_2334),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_3062),
.A2(n_2918),
.B1(n_2870),
.B2(n_2675),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_3075),
.A2(n_1837),
.B1(n_1835),
.B2(n_2675),
.Y(n_3195)
);

AOI22xp33_ASAP7_75t_L g3196 ( 
.A1(n_2989),
.A2(n_1837),
.B1(n_1835),
.B2(n_2675),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_3034),
.A2(n_1943),
.B1(n_1748),
.B2(n_1789),
.Y(n_3197)
);

OAI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_3044),
.A2(n_2755),
.B1(n_2746),
.B2(n_2719),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2986),
.B(n_2622),
.Y(n_3199)
);

NAND3xp33_ASAP7_75t_L g3200 ( 
.A(n_3120),
.B(n_2833),
.C(n_2719),
.Y(n_3200)
);

NAND3xp33_ASAP7_75t_L g3201 ( 
.A(n_2978),
.B(n_2719),
.C(n_1872),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3079),
.A2(n_3088),
.B1(n_3084),
.B2(n_3070),
.Y(n_3202)
);

AOI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3086),
.A2(n_2957),
.B1(n_2555),
.B2(n_1748),
.Y(n_3203)
);

AND2x2_ASAP7_75t_L g3204 ( 
.A(n_3069),
.B(n_2624),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_3037),
.A2(n_2678),
.B1(n_2687),
.B2(n_2662),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3089),
.A2(n_2678),
.B1(n_2687),
.B2(n_2662),
.Y(n_3206)
);

NAND3xp33_ASAP7_75t_L g3207 ( 
.A(n_3093),
.B(n_3018),
.C(n_3051),
.Y(n_3207)
);

NOR2xp67_ASAP7_75t_L g3208 ( 
.A(n_3078),
.B(n_2925),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_3089),
.A2(n_2678),
.B1(n_2687),
.B2(n_2662),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_SL g3210 ( 
.A1(n_2982),
.A2(n_2950),
.B1(n_2862),
.B2(n_2880),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_3071),
.A2(n_1943),
.B1(n_1789),
.B2(n_1695),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_3009),
.A2(n_1943),
.B1(n_1871),
.B2(n_2624),
.Y(n_3212)
);

AOI22xp33_ASAP7_75t_L g3213 ( 
.A1(n_3055),
.A2(n_3083),
.B1(n_3054),
.B2(n_3115),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3003),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_3127),
.A2(n_2631),
.B1(n_2221),
.B2(n_2150),
.Y(n_3215)
);

HB1xp67_ASAP7_75t_L g3216 ( 
.A(n_3027),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_3117),
.A2(n_2631),
.B1(n_2221),
.B2(n_2150),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3072),
.A2(n_2074),
.B1(n_2386),
.B2(n_2153),
.Y(n_3218)
);

OAI21xp5_ASAP7_75t_SL g3219 ( 
.A1(n_3125),
.A2(n_2852),
.B(n_2768),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3082),
.B(n_2842),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3085),
.B(n_2842),
.Y(n_3221)
);

AOI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3035),
.A2(n_2074),
.B1(n_1840),
.B2(n_2914),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_3016),
.A2(n_2386),
.B1(n_2153),
.B2(n_2936),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_L g3224 ( 
.A1(n_3124),
.A2(n_2386),
.B1(n_2936),
.B2(n_2950),
.Y(n_3224)
);

OAI22xp5_ASAP7_75t_L g3225 ( 
.A1(n_3035),
.A2(n_3125),
.B1(n_3137),
.B2(n_3024),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_3143),
.A2(n_2936),
.B1(n_2862),
.B2(n_2880),
.Y(n_3226)
);

AOI222xp33_ASAP7_75t_L g3227 ( 
.A1(n_2982),
.A2(n_2884),
.B1(n_2768),
.B2(n_2756),
.C1(n_2134),
.C2(n_2166),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3106),
.A2(n_2950),
.B1(n_2880),
.B2(n_2862),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_SL g3229 ( 
.A1(n_2982),
.A2(n_2756),
.B1(n_2476),
.B2(n_2694),
.Y(n_3229)
);

AOI22xp33_ASAP7_75t_SL g3230 ( 
.A1(n_3056),
.A2(n_2470),
.B1(n_2694),
.B2(n_2673),
.Y(n_3230)
);

OAI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_3137),
.A2(n_3149),
.B1(n_3128),
.B2(n_3011),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_3138),
.A2(n_2265),
.B1(n_2194),
.B2(n_2208),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_3017),
.A2(n_2260),
.B1(n_2228),
.B2(n_2211),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3058),
.B(n_311),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_L g3235 ( 
.A1(n_3094),
.A2(n_2032),
.B1(n_2034),
.B2(n_2021),
.Y(n_3235)
);

OAI21xp5_ASAP7_75t_SL g3236 ( 
.A1(n_2979),
.A2(n_2021),
.B(n_2017),
.Y(n_3236)
);

NAND3xp33_ASAP7_75t_L g3237 ( 
.A(n_3113),
.B(n_2038),
.C(n_2034),
.Y(n_3237)
);

AOI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_2988),
.A2(n_1840),
.B1(n_1799),
.B2(n_1881),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3030),
.Y(n_3239)
);

AOI22xp33_ASAP7_75t_L g3240 ( 
.A1(n_3096),
.A2(n_2032),
.B1(n_2088),
.B2(n_2103),
.Y(n_3240)
);

AOI22xp33_ASAP7_75t_SL g3241 ( 
.A1(n_3098),
.A2(n_2436),
.B1(n_2694),
.B2(n_2673),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3091),
.B(n_311),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3039),
.A2(n_2088),
.B1(n_2103),
.B2(n_2107),
.Y(n_3243)
);

AOI22xp33_ASAP7_75t_SL g3244 ( 
.A1(n_3098),
.A2(n_2447),
.B1(n_2673),
.B2(n_2628),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_3116),
.A2(n_1840),
.B1(n_1799),
.B2(n_1882),
.Y(n_3245)
);

NOR2xp33_ASAP7_75t_L g3246 ( 
.A(n_3097),
.B(n_312),
.Y(n_3246)
);

AOI22xp33_ASAP7_75t_L g3247 ( 
.A1(n_3087),
.A2(n_2107),
.B1(n_2136),
.B2(n_2147),
.Y(n_3247)
);

NAND3xp33_ASAP7_75t_L g3248 ( 
.A(n_3123),
.B(n_2436),
.C(n_2427),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_3095),
.A2(n_2136),
.B1(n_2147),
.B2(n_2087),
.Y(n_3249)
);

AOI22xp5_ASAP7_75t_L g3250 ( 
.A1(n_3122),
.A2(n_1882),
.B1(n_2087),
.B2(n_1850),
.Y(n_3250)
);

AOI22xp5_ASAP7_75t_L g3251 ( 
.A1(n_3090),
.A2(n_1850),
.B1(n_2628),
.B2(n_2606),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3099),
.B(n_313),
.Y(n_3252)
);

AOI22xp33_ASAP7_75t_L g3253 ( 
.A1(n_3028),
.A2(n_2337),
.B1(n_2349),
.B2(n_2372),
.Y(n_3253)
);

OAI22xp5_ASAP7_75t_L g3254 ( 
.A1(n_3081),
.A2(n_2494),
.B1(n_2628),
.B2(n_2606),
.Y(n_3254)
);

NAND3xp33_ASAP7_75t_L g3255 ( 
.A(n_3123),
.B(n_2447),
.C(n_2436),
.Y(n_3255)
);

OAI21xp33_ASAP7_75t_L g3256 ( 
.A1(n_3036),
.A2(n_313),
.B(n_314),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3008),
.A2(n_2337),
.B1(n_2349),
.B2(n_2372),
.Y(n_3257)
);

AOI22xp33_ASAP7_75t_L g3258 ( 
.A1(n_2993),
.A2(n_2494),
.B1(n_2606),
.B2(n_2559),
.Y(n_3258)
);

OAI222xp33_ASAP7_75t_L g3259 ( 
.A1(n_3004),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.C1(n_318),
.C2(n_319),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_3103),
.A2(n_2494),
.B1(n_2559),
.B2(n_2526),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3153),
.B(n_3216),
.Y(n_3261)
);

NOR3xp33_ASAP7_75t_L g3262 ( 
.A(n_3231),
.B(n_3078),
.C(n_3146),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3156),
.B(n_3114),
.Y(n_3263)
);

OAI21xp5_ASAP7_75t_SL g3264 ( 
.A1(n_3219),
.A2(n_3023),
.B(n_3139),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3156),
.Y(n_3265)
);

NAND2x1p5_ASAP7_75t_L g3266 ( 
.A(n_3157),
.B(n_3015),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3161),
.B(n_3118),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3170),
.B(n_3173),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3214),
.B(n_3119),
.Y(n_3269)
);

AOI22xp33_ASAP7_75t_L g3270 ( 
.A1(n_3175),
.A2(n_3133),
.B1(n_3134),
.B2(n_3151),
.Y(n_3270)
);

NAND3xp33_ASAP7_75t_SL g3271 ( 
.A(n_3227),
.B(n_3080),
.C(n_3060),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_SL g3272 ( 
.A1(n_3225),
.A2(n_3098),
.B1(n_3041),
.B2(n_3014),
.Y(n_3272)
);

OAI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3158),
.A2(n_3147),
.B1(n_3145),
.B2(n_3102),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3204),
.B(n_3057),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_3190),
.B(n_3141),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3158),
.A2(n_3140),
.B1(n_3107),
.B2(n_3129),
.Y(n_3276)
);

AOI211xp5_ASAP7_75t_L g3277 ( 
.A1(n_3231),
.A2(n_3198),
.B(n_3165),
.C(n_3162),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3216),
.B(n_3061),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_3259),
.A2(n_3068),
.B(n_3112),
.Y(n_3279)
);

NAND3xp33_ASAP7_75t_L g3280 ( 
.A(n_3152),
.B(n_2994),
.C(n_2980),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3239),
.B(n_3104),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_SL g3282 ( 
.A(n_3157),
.B(n_3042),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3191),
.B(n_2980),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3199),
.B(n_2994),
.Y(n_3284)
);

OAI221xp5_ASAP7_75t_L g3285 ( 
.A1(n_3152),
.A2(n_2998),
.B1(n_3007),
.B2(n_3109),
.C(n_3077),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3167),
.B(n_2994),
.Y(n_3286)
);

NAND3xp33_ASAP7_75t_L g3287 ( 
.A(n_3155),
.B(n_3046),
.C(n_3013),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_3207),
.B(n_3013),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_3234),
.B(n_3174),
.Y(n_3289)
);

OAI21xp33_ASAP7_75t_L g3290 ( 
.A1(n_3178),
.A2(n_3048),
.B(n_2987),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3169),
.B(n_3126),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3166),
.B(n_3148),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3172),
.B(n_3013),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3202),
.A2(n_3073),
.B1(n_3129),
.B2(n_3029),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3213),
.B(n_3220),
.Y(n_3295)
);

NAND3xp33_ASAP7_75t_L g3296 ( 
.A(n_3179),
.B(n_3046),
.C(n_3142),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3221),
.B(n_3121),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_SL g3298 ( 
.A1(n_3176),
.A2(n_3005),
.B1(n_3101),
.B2(n_3050),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3230),
.B(n_3046),
.Y(n_3299)
);

NAND3xp33_ASAP7_75t_L g3300 ( 
.A(n_3246),
.B(n_3135),
.C(n_3064),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3192),
.B(n_3136),
.Y(n_3301)
);

OAI21xp5_ASAP7_75t_SL g3302 ( 
.A1(n_3182),
.A2(n_3100),
.B(n_3105),
.Y(n_3302)
);

OAI221xp5_ASAP7_75t_L g3303 ( 
.A1(n_3177),
.A2(n_3150),
.B1(n_3067),
.B2(n_3064),
.C(n_3001),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3242),
.B(n_3252),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_SL g3305 ( 
.A(n_3222),
.B(n_3001),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3171),
.B(n_3067),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3160),
.B(n_3144),
.Y(n_3307)
);

NAND3xp33_ASAP7_75t_L g3308 ( 
.A(n_3164),
.B(n_3131),
.C(n_3130),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3181),
.Y(n_3309)
);

OAI221xp5_ASAP7_75t_SL g3310 ( 
.A1(n_3193),
.A2(n_3026),
.B1(n_316),
.B2(n_317),
.C(n_318),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3160),
.B(n_3130),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3159),
.A2(n_3130),
.B1(n_2496),
.B2(n_2559),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3187),
.B(n_315),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3228),
.B(n_319),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3185),
.B(n_3183),
.Y(n_3315)
);

INVx1_ASAP7_75t_SL g3316 ( 
.A(n_3261),
.Y(n_3316)
);

NAND3xp33_ASAP7_75t_L g3317 ( 
.A(n_3288),
.B(n_3200),
.C(n_3180),
.Y(n_3317)
);

AOI221xp5_ASAP7_75t_L g3318 ( 
.A1(n_3270),
.A2(n_3256),
.B1(n_3154),
.B2(n_3168),
.C(n_3194),
.Y(n_3318)
);

NAND4xp75_ASAP7_75t_L g3319 ( 
.A(n_3306),
.B(n_3208),
.C(n_3203),
.D(n_3188),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3263),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3261),
.B(n_3275),
.Y(n_3321)
);

AND2x2_ASAP7_75t_L g3322 ( 
.A(n_3281),
.B(n_3274),
.Y(n_3322)
);

NAND3xp33_ASAP7_75t_L g3323 ( 
.A(n_3288),
.B(n_3159),
.C(n_3201),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3265),
.B(n_3224),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3281),
.B(n_3286),
.Y(n_3325)
);

AOI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3262),
.A2(n_3194),
.B1(n_3184),
.B2(n_3232),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3262),
.A2(n_3189),
.B1(n_3237),
.B2(n_3254),
.Y(n_3327)
);

NAND3xp33_ASAP7_75t_L g3328 ( 
.A(n_3277),
.B(n_3163),
.C(n_3248),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3284),
.B(n_3289),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3270),
.B(n_3309),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3268),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_3278),
.B(n_3255),
.Y(n_3332)
);

OR2x2_ASAP7_75t_L g3333 ( 
.A(n_3267),
.B(n_3260),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_L g3334 ( 
.A(n_3272),
.B(n_3236),
.C(n_3209),
.Y(n_3334)
);

NOR4xp75_ASAP7_75t_L g3335 ( 
.A(n_3271),
.B(n_3206),
.C(n_3205),
.D(n_3229),
.Y(n_3335)
);

NAND3xp33_ASAP7_75t_L g3336 ( 
.A(n_3279),
.B(n_3260),
.C(n_3226),
.Y(n_3336)
);

AOI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3273),
.A2(n_3238),
.B1(n_3250),
.B2(n_3210),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3269),
.B(n_3251),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_3311),
.B(n_3283),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3311),
.B(n_3218),
.Y(n_3340)
);

HB1xp67_ASAP7_75t_L g3341 ( 
.A(n_3291),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3295),
.B(n_3212),
.Y(n_3342)
);

NAND4xp75_ASAP7_75t_L g3343 ( 
.A(n_3299),
.B(n_3245),
.C(n_3186),
.D(n_3244),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3307),
.B(n_3240),
.Y(n_3344)
);

NOR2x1_ASAP7_75t_L g3345 ( 
.A(n_3264),
.B(n_3241),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3297),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3301),
.B(n_3249),
.Y(n_3347)
);

OR2x2_ASAP7_75t_SL g3348 ( 
.A(n_3280),
.B(n_3258),
.Y(n_3348)
);

AO21x2_ASAP7_75t_L g3349 ( 
.A1(n_3305),
.A2(n_3197),
.B(n_3217),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3266),
.A2(n_3258),
.B1(n_3243),
.B2(n_3223),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3304),
.B(n_3233),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3293),
.B(n_3253),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3266),
.B(n_3215),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3292),
.B(n_3247),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3294),
.B(n_3196),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_L g3356 ( 
.A(n_3290),
.B(n_3235),
.Y(n_3356)
);

NOR3xp33_ASAP7_75t_L g3357 ( 
.A(n_3298),
.B(n_320),
.C(n_321),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3339),
.B(n_3299),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3346),
.Y(n_3359)
);

XOR2x2_ASAP7_75t_L g3360 ( 
.A(n_3345),
.B(n_3287),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3341),
.B(n_3294),
.Y(n_3361)
);

OR2x2_ASAP7_75t_L g3362 ( 
.A(n_3316),
.B(n_3305),
.Y(n_3362)
);

INVx1_ASAP7_75t_SL g3363 ( 
.A(n_3325),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3322),
.Y(n_3364)
);

INVx3_ASAP7_75t_L g3365 ( 
.A(n_3322),
.Y(n_3365)
);

NOR3xp33_ASAP7_75t_L g3366 ( 
.A(n_3357),
.B(n_3310),
.C(n_3314),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3321),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3346),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3339),
.B(n_3325),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3356),
.A2(n_3282),
.B1(n_3302),
.B2(n_3276),
.Y(n_3370)
);

NAND4xp75_ASAP7_75t_L g3371 ( 
.A(n_3356),
.B(n_3315),
.C(n_3313),
.D(n_3312),
.Y(n_3371)
);

INVx2_ASAP7_75t_SL g3372 ( 
.A(n_3321),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3329),
.B(n_3308),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_3320),
.B(n_3300),
.Y(n_3374)
);

NAND4xp75_ASAP7_75t_L g3375 ( 
.A(n_3318),
.B(n_3296),
.C(n_3285),
.D(n_3303),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3332),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3331),
.Y(n_3377)
);

XNOR2x2_ASAP7_75t_L g3378 ( 
.A(n_3319),
.B(n_3257),
.Y(n_3378)
);

INVx1_ASAP7_75t_SL g3379 ( 
.A(n_3333),
.Y(n_3379)
);

NAND3xp33_ASAP7_75t_SL g3380 ( 
.A(n_3335),
.B(n_3211),
.C(n_3195),
.Y(n_3380)
);

NAND4xp75_ASAP7_75t_SL g3381 ( 
.A(n_3353),
.B(n_320),
.C(n_321),
.D(n_322),
.Y(n_3381)
);

XOR2x2_ASAP7_75t_L g3382 ( 
.A(n_3334),
.B(n_322),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3338),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3341),
.Y(n_3384)
);

INVx2_ASAP7_75t_SL g3385 ( 
.A(n_3352),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3330),
.Y(n_3386)
);

XNOR2xp5_ASAP7_75t_L g3387 ( 
.A(n_3328),
.B(n_324),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3340),
.B(n_2447),
.Y(n_3388)
);

NOR4xp25_ASAP7_75t_L g3389 ( 
.A(n_3323),
.B(n_324),
.C(n_325),
.D(n_326),
.Y(n_3389)
);

NAND4xp75_ASAP7_75t_L g3390 ( 
.A(n_3337),
.B(n_326),
.C(n_327),
.D(n_328),
.Y(n_3390)
);

NOR4xp75_ASAP7_75t_L g3391 ( 
.A(n_3343),
.B(n_3355),
.C(n_3350),
.D(n_3342),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3324),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3351),
.Y(n_3393)
);

NAND4xp75_ASAP7_75t_L g3394 ( 
.A(n_3340),
.B(n_328),
.C(n_329),
.D(n_330),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3347),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3344),
.B(n_330),
.Y(n_3396)
);

NAND4xp75_ASAP7_75t_SL g3397 ( 
.A(n_3348),
.B(n_3336),
.C(n_3327),
.D(n_3354),
.Y(n_3397)
);

BUFx3_ASAP7_75t_L g3398 ( 
.A(n_3365),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3365),
.Y(n_3399)
);

XOR2x2_ASAP7_75t_L g3400 ( 
.A(n_3382),
.B(n_3397),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3383),
.Y(n_3401)
);

XOR2x2_ASAP7_75t_L g3402 ( 
.A(n_3382),
.B(n_3326),
.Y(n_3402)
);

AO22x2_ASAP7_75t_L g3403 ( 
.A1(n_3397),
.A2(n_3317),
.B1(n_3354),
.B2(n_3352),
.Y(n_3403)
);

AND2x4_ASAP7_75t_L g3404 ( 
.A(n_3383),
.B(n_3349),
.Y(n_3404)
);

HB1xp67_ASAP7_75t_L g3405 ( 
.A(n_3376),
.Y(n_3405)
);

XOR2x2_ASAP7_75t_L g3406 ( 
.A(n_3391),
.B(n_3326),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3386),
.B(n_3349),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3359),
.Y(n_3408)
);

XNOR2xp5_ASAP7_75t_L g3409 ( 
.A(n_3360),
.B(n_3327),
.Y(n_3409)
);

INVx1_ASAP7_75t_SL g3410 ( 
.A(n_3379),
.Y(n_3410)
);

XNOR2x1_ASAP7_75t_L g3411 ( 
.A(n_3360),
.B(n_331),
.Y(n_3411)
);

XNOR2xp5_ASAP7_75t_L g3412 ( 
.A(n_3370),
.B(n_332),
.Y(n_3412)
);

NAND2x1_ASAP7_75t_L g3413 ( 
.A(n_3358),
.B(n_2470),
.Y(n_3413)
);

XOR2x2_ASAP7_75t_L g3414 ( 
.A(n_3378),
.B(n_333),
.Y(n_3414)
);

XOR2x2_ASAP7_75t_L g3415 ( 
.A(n_3387),
.B(n_334),
.Y(n_3415)
);

XOR2x2_ASAP7_75t_L g3416 ( 
.A(n_3375),
.B(n_335),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3368),
.Y(n_3417)
);

INVxp67_ASAP7_75t_L g3418 ( 
.A(n_3393),
.Y(n_3418)
);

XOR2x2_ASAP7_75t_L g3419 ( 
.A(n_3381),
.B(n_335),
.Y(n_3419)
);

OA22x2_ASAP7_75t_L g3420 ( 
.A1(n_3385),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_3420)
);

XNOR2x2_ASAP7_75t_L g3421 ( 
.A(n_3371),
.B(n_339),
.Y(n_3421)
);

XNOR2x1_ASAP7_75t_L g3422 ( 
.A(n_3390),
.B(n_339),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3398),
.Y(n_3423)
);

INVx4_ASAP7_75t_SL g3424 ( 
.A(n_3416),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3403),
.A2(n_3385),
.B1(n_3361),
.B2(n_3363),
.Y(n_3425)
);

OAI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3403),
.A2(n_3409),
.B1(n_3410),
.B2(n_3411),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3405),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3401),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3413),
.Y(n_3429)
);

INVx1_ASAP7_75t_SL g3430 ( 
.A(n_3420),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3399),
.B(n_3376),
.Y(n_3431)
);

INVx2_ASAP7_75t_SL g3432 ( 
.A(n_3400),
.Y(n_3432)
);

AND2x4_ASAP7_75t_L g3433 ( 
.A(n_3418),
.B(n_3377),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3408),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3408),
.Y(n_3435)
);

XNOR2xp5_ASAP7_75t_L g3436 ( 
.A(n_3414),
.B(n_3381),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3417),
.Y(n_3437)
);

AOI22xp5_ASAP7_75t_L g3438 ( 
.A1(n_3402),
.A2(n_3380),
.B1(n_3366),
.B2(n_3395),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3417),
.Y(n_3439)
);

OA22x2_ASAP7_75t_L g3440 ( 
.A1(n_3412),
.A2(n_3361),
.B1(n_3392),
.B2(n_3373),
.Y(n_3440)
);

INVx1_ASAP7_75t_SL g3441 ( 
.A(n_3421),
.Y(n_3441)
);

OA22x2_ASAP7_75t_L g3442 ( 
.A1(n_3404),
.A2(n_3407),
.B1(n_3406),
.B2(n_3413),
.Y(n_3442)
);

CKINVDCx14_ASAP7_75t_R g3443 ( 
.A(n_3415),
.Y(n_3443)
);

INVx3_ASAP7_75t_SL g3444 ( 
.A(n_3419),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3404),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3422),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3410),
.Y(n_3447)
);

OA22x2_ASAP7_75t_L g3448 ( 
.A1(n_3409),
.A2(n_3384),
.B1(n_3372),
.B2(n_3364),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3398),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3447),
.Y(n_3450)
);

XOR2x2_ASAP7_75t_L g3451 ( 
.A(n_3444),
.B(n_3380),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3427),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3434),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3435),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3433),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3433),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3423),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3449),
.Y(n_3458)
);

INVxp67_ASAP7_75t_L g3459 ( 
.A(n_3446),
.Y(n_3459)
);

INVx1_ASAP7_75t_SL g3460 ( 
.A(n_3441),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3437),
.Y(n_3461)
);

BUFx2_ASAP7_75t_L g3462 ( 
.A(n_3448),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3439),
.Y(n_3463)
);

OA22x2_ASAP7_75t_L g3464 ( 
.A1(n_3426),
.A2(n_3364),
.B1(n_3367),
.B2(n_3369),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3445),
.Y(n_3465)
);

HB1xp67_ASAP7_75t_L g3466 ( 
.A(n_3441),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3431),
.Y(n_3467)
);

OAI322xp33_ASAP7_75t_L g3468 ( 
.A1(n_3426),
.A2(n_3374),
.A3(n_3396),
.B1(n_3362),
.B2(n_3367),
.C1(n_3389),
.C2(n_3366),
.Y(n_3468)
);

AOI22x1_ASAP7_75t_L g3469 ( 
.A1(n_3466),
.A2(n_3432),
.B1(n_3436),
.B2(n_3430),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3466),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3457),
.Y(n_3471)
);

INVxp67_ASAP7_75t_L g3472 ( 
.A(n_3460),
.Y(n_3472)
);

INVx1_ASAP7_75t_SL g3473 ( 
.A(n_3460),
.Y(n_3473)
);

AOI22xp33_ASAP7_75t_L g3474 ( 
.A1(n_3464),
.A2(n_3440),
.B1(n_3448),
.B2(n_3425),
.Y(n_3474)
);

AO22x2_ASAP7_75t_L g3475 ( 
.A1(n_3459),
.A2(n_3424),
.B1(n_3425),
.B2(n_3430),
.Y(n_3475)
);

AOI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3464),
.A2(n_3440),
.B1(n_3438),
.B2(n_3424),
.Y(n_3476)
);

AOI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3462),
.A2(n_3438),
.B1(n_3442),
.B2(n_3443),
.Y(n_3477)
);

AOI31xp33_ASAP7_75t_L g3478 ( 
.A1(n_3459),
.A2(n_3442),
.A3(n_3428),
.B(n_3394),
.Y(n_3478)
);

OAI222xp33_ASAP7_75t_L g3479 ( 
.A1(n_3465),
.A2(n_3429),
.B1(n_3388),
.B2(n_342),
.C1(n_344),
.C2(n_345),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3458),
.Y(n_3480)
);

AOI22xp5_ASAP7_75t_L g3481 ( 
.A1(n_3451),
.A2(n_3455),
.B1(n_3456),
.B2(n_3450),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3452),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3453),
.Y(n_3483)
);

AOI22xp5_ASAP7_75t_L g3484 ( 
.A1(n_3467),
.A2(n_3429),
.B1(n_2496),
.B2(n_2526),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3470),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3473),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3472),
.Y(n_3487)
);

OA22x2_ASAP7_75t_SL g3488 ( 
.A1(n_3469),
.A2(n_3468),
.B1(n_3454),
.B2(n_3461),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3471),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3480),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3482),
.Y(n_3491)
);

O2A1O1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_3478),
.A2(n_3463),
.B(n_341),
.C(n_345),
.Y(n_3492)
);

AND4x1_ASAP7_75t_L g3493 ( 
.A(n_3477),
.B(n_340),
.C(n_341),
.D(n_346),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3475),
.Y(n_3494)
);

INVxp67_ASAP7_75t_SL g3495 ( 
.A(n_3481),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3475),
.Y(n_3496)
);

AOI211xp5_ASAP7_75t_SL g3497 ( 
.A1(n_3476),
.A2(n_3479),
.B(n_3483),
.C(n_3484),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3486),
.Y(n_3498)
);

AOI22xp5_ASAP7_75t_L g3499 ( 
.A1(n_3495),
.A2(n_3474),
.B1(n_2496),
.B2(n_2526),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3495),
.B(n_346),
.Y(n_3500)
);

OAI221xp5_ASAP7_75t_L g3501 ( 
.A1(n_3488),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.C(n_350),
.Y(n_3501)
);

AOI221xp5_ASAP7_75t_L g3502 ( 
.A1(n_3492),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.C(n_351),
.Y(n_3502)
);

NOR4xp25_ASAP7_75t_L g3503 ( 
.A(n_3494),
.B(n_352),
.C(n_353),
.D(n_355),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3493),
.B(n_352),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3487),
.A2(n_2476),
.B1(n_2522),
.B2(n_2507),
.Y(n_3505)
);

OA22x2_ASAP7_75t_L g3506 ( 
.A1(n_3496),
.A2(n_353),
.B1(n_356),
.B2(n_357),
.Y(n_3506)
);

AOI22xp5_ASAP7_75t_L g3507 ( 
.A1(n_3485),
.A2(n_2476),
.B1(n_2522),
.B2(n_2507),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3489),
.Y(n_3508)
);

INVxp67_ASAP7_75t_SL g3509 ( 
.A(n_3504),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3498),
.Y(n_3510)
);

AOI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_3501),
.A2(n_3490),
.B1(n_3491),
.B2(n_3497),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3506),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3500),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_SL g3514 ( 
.A(n_3508),
.B(n_3492),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3499),
.B(n_358),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3502),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3503),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3507),
.B(n_359),
.Y(n_3518)
);

INVx1_ASAP7_75t_SL g3519 ( 
.A(n_3505),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3512),
.Y(n_3520)
);

AOI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_3516),
.A2(n_2477),
.B1(n_2522),
.B2(n_2507),
.Y(n_3521)
);

NAND4xp25_ASAP7_75t_L g3522 ( 
.A(n_3511),
.B(n_3514),
.C(n_3517),
.D(n_3519),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_3509),
.Y(n_3523)
);

INVx4_ASAP7_75t_L g3524 ( 
.A(n_3510),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3515),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3520),
.Y(n_3526)
);

NOR2x1_ASAP7_75t_L g3527 ( 
.A(n_3522),
.B(n_3513),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_SL g3528 ( 
.A1(n_3523),
.A2(n_3518),
.B1(n_360),
.B2(n_2501),
.Y(n_3528)
);

OAI211xp5_ASAP7_75t_L g3529 ( 
.A1(n_3524),
.A2(n_360),
.B(n_2501),
.C(n_2477),
.Y(n_3529)
);

OAI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3525),
.A2(n_2501),
.B1(n_2477),
.B2(n_2470),
.Y(n_3530)
);

AOI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3521),
.A2(n_2708),
.B1(n_2373),
.B2(n_2372),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3528),
.Y(n_3532)
);

OAI22x1_ASAP7_75t_L g3533 ( 
.A1(n_3527),
.A2(n_482),
.B1(n_483),
.B2(n_486),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3526),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3534),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3532),
.Y(n_3536)
);

AOI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3536),
.A2(n_3529),
.B1(n_3533),
.B2(n_3530),
.Y(n_3537)
);

INVxp67_ASAP7_75t_L g3538 ( 
.A(n_3537),
.Y(n_3538)
);

AOI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_3538),
.A2(n_3535),
.B1(n_3531),
.B2(n_2708),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3539),
.Y(n_3540)
);

AOI221xp5_ASAP7_75t_L g3541 ( 
.A1(n_3540),
.A2(n_2708),
.B1(n_2373),
.B2(n_2349),
.C(n_495),
.Y(n_3541)
);

AOI211xp5_ASAP7_75t_L g3542 ( 
.A1(n_3541),
.A2(n_487),
.B(n_491),
.C(n_494),
.Y(n_3542)
);


endmodule