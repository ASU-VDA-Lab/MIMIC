module fake_jpeg_13257_n_482 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_482);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_482;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_17),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_10),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_58),
.B(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_61),
.Y(n_128)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_66),
.Y(n_182)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_21),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_71),
.B(n_78),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_18),
.Y(n_76)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_93),
.Y(n_162)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_34),
.A2(n_1),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_27),
.B(n_13),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_51),
.Y(n_100)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_43),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_103),
.Y(n_195)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_10),
.Y(n_103)
);

INVx2_ASAP7_75t_R g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_49),
.B(n_1),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_26),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_30),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_111),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_26),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_114),
.B(n_115),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_4),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_35),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_120),
.Y(n_187)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_23),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_57),
.B1(n_56),
.B2(n_42),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_122),
.A2(n_132),
.B(n_135),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_108),
.B1(n_99),
.B2(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_123),
.A2(n_130),
.B1(n_136),
.B2(n_142),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_28),
.B1(n_56),
.B2(n_22),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_57),
.B1(n_22),
.B2(n_42),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_55),
.B1(n_54),
.B2(n_46),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_55),
.B1(n_28),
.B2(n_47),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_66),
.A2(n_55),
.B1(n_28),
.B2(n_47),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_41),
.B1(n_25),
.B2(n_29),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_153),
.B1(n_160),
.B2(n_177),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_41),
.B1(n_25),
.B2(n_29),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_148),
.A2(n_164),
.B1(n_193),
.B2(n_135),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_39),
.B1(n_33),
.B2(n_38),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_65),
.A2(n_35),
.B1(n_46),
.B2(n_39),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_157),
.A2(n_170),
.B(n_179),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_33),
.B1(n_35),
.B2(n_46),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_50),
.B1(n_46),
.B2(n_7),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_116),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_63),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_64),
.A2(n_100),
.B1(n_70),
.B2(n_80),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_189),
.B1(n_191),
.B2(n_121),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_77),
.B(n_104),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_188),
.B(n_181),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_83),
.A2(n_107),
.B1(n_74),
.B2(n_82),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_175),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_119),
.A2(n_89),
.B1(n_76),
.B2(n_77),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_94),
.A2(n_59),
.B1(n_52),
.B2(n_78),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_196),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_199),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_200),
.A2(n_205),
.B(n_209),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

AND2x4_ASAP7_75t_SL g203 ( 
.A(n_139),
.B(n_174),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_203),
.B(n_224),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_129),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_128),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_207),
.B(n_216),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_126),
.A2(n_163),
.B1(n_138),
.B2(n_192),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_210),
.A2(n_211),
.B1(n_244),
.B2(n_247),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_169),
.B1(n_194),
.B2(n_155),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_125),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g309 ( 
.A(n_214),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_150),
.B(n_145),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_195),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_152),
.B(n_137),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_203),
.C(n_251),
.Y(n_271)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_158),
.Y(n_220)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_161),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_222),
.B(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_157),
.B(n_172),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_223),
.A2(n_198),
.B(n_231),
.Y(n_305)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_136),
.A2(n_142),
.B1(n_123),
.B2(n_156),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_231),
.B1(n_257),
.B2(n_204),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_227),
.Y(n_261)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_228),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_236),
.Y(n_267)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_230),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_131),
.A2(n_159),
.B1(n_168),
.B2(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_235),
.B(n_238),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_158),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_245),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_140),
.B(n_121),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_131),
.B(n_159),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_240),
.B(n_258),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_164),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_241),
.B(n_246),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_242),
.Y(n_300)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_121),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_155),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_122),
.A2(n_132),
.B1(n_179),
.B2(n_168),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_170),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_248),
.B(n_253),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_182),
.B(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_254),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_151),
.B(n_178),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_151),
.A2(n_142),
.B1(n_136),
.B2(n_123),
.Y(n_252)
);

AO21x2_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_239),
.B(n_249),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_151),
.B(n_178),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_221),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_128),
.B(n_58),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_259),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_136),
.A2(n_142),
.B1(n_99),
.B2(n_108),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_133),
.B(n_128),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_128),
.B(n_58),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_234),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_244),
.B(n_223),
.C(n_232),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_271),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_200),
.A2(n_254),
.B1(n_233),
.B2(n_252),
.Y(n_263)
);

AO21x2_ASAP7_75t_L g311 ( 
.A1(n_263),
.A2(n_265),
.B(n_196),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_204),
.B1(n_219),
.B2(n_205),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_250),
.B1(n_227),
.B2(n_259),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_205),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_270),
.B(n_294),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_277),
.A2(n_282),
.B1(n_297),
.B2(n_271),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_209),
.B(n_203),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_285),
.B(n_307),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_237),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_299),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_202),
.B(n_212),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_214),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_305),
.A2(n_268),
.B(n_306),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_198),
.B(n_196),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_224),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_230),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_318),
.B1(n_323),
.B2(n_330),
.Y(n_355)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_287),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_324),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_308),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_264),
.A2(n_245),
.B1(n_217),
.B2(n_199),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_319),
.A2(n_344),
.B1(n_283),
.B2(n_309),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_218),
.B(n_243),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_320),
.A2(n_321),
.B(n_337),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_228),
.B(n_243),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_331),
.B(n_292),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_206),
.B1(n_208),
.B2(n_213),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_224),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_326),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_286),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_329),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_242),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_242),
.B1(n_262),
.B2(n_264),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_305),
.B(n_288),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_262),
.B1(n_282),
.B2(n_285),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_334),
.A2(n_290),
.B1(n_293),
.B2(n_295),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_281),
.B(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_339),
.A2(n_343),
.B1(n_292),
.B2(n_279),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_280),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_281),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_341),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_277),
.A2(n_261),
.B1(n_279),
.B2(n_278),
.Y(n_343)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_345),
.A2(n_309),
.B(n_296),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_347),
.A2(n_348),
.B(n_370),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_339),
.A2(n_292),
.B1(n_272),
.B2(n_284),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_351),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_284),
.B1(n_290),
.B2(n_295),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_357),
.A2(n_311),
.B1(n_327),
.B2(n_328),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_346),
.A2(n_293),
.B(n_275),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_358),
.A2(n_361),
.B(n_323),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_275),
.B(n_276),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_300),
.C(n_276),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_321),
.C(n_333),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_300),
.B(n_283),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_369),
.B(n_320),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_310),
.A2(n_291),
.B1(n_315),
.B2(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_336),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_371),
.Y(n_375)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_368),
.B(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_373),
.B(n_385),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_374),
.A2(n_361),
.B(n_352),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_378),
.C(n_379),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_377),
.A2(n_311),
.B1(n_351),
.B2(n_365),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_313),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_313),
.C(n_331),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_329),
.C(n_310),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_383),
.C(n_384),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_348),
.C(n_370),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_317),
.C(n_325),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_354),
.B(n_335),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_386),
.A2(n_390),
.B(n_367),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_314),
.Y(n_387)
);

AOI21xp33_ASAP7_75t_L g417 ( 
.A1(n_387),
.A2(n_388),
.B(n_393),
.Y(n_417)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_363),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_317),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_391),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_361),
.A2(n_330),
.B(n_322),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_324),
.C(n_314),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_332),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_312),
.Y(n_394)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_394),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_332),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_401),
.A2(n_411),
.B(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_381),
.A2(n_361),
.B1(n_355),
.B2(n_365),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_405),
.A2(n_395),
.B1(n_311),
.B2(n_347),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_376),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_409),
.Y(n_419)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_392),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_413),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_353),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_353),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_410),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_384),
.B(n_350),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_414),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_347),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_416),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_357),
.Y(n_416)
);

BUFx12_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_430),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_383),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_434),
.C(n_406),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_416),
.B(n_396),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_374),
.B(n_367),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_427),
.B(n_431),
.Y(n_448)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_429),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_418),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_363),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_396),
.B1(n_395),
.B2(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_432),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_358),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_435),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_381),
.C(n_358),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_362),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_415),
.Y(n_437)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_437),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_422),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_427),
.B(n_425),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_404),
.C(n_406),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_443),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_428),
.A2(n_400),
.B1(n_311),
.B2(n_399),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_442),
.A2(n_444),
.B1(n_445),
.B2(n_429),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_404),
.C(n_414),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_400),
.B1(n_311),
.B2(n_412),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_426),
.A2(n_413),
.B1(n_381),
.B2(n_356),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_440),
.B(n_437),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_432),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_456),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_453),
.C(n_441),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_422),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_398),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_454),
.B(n_455),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_398),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_457),
.B(n_420),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_458),
.B(n_420),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_449),
.B(n_426),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_465),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_463),
.B(n_464),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_450),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_439),
.C(n_419),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g473 ( 
.A1(n_467),
.A2(n_471),
.A3(n_421),
.B1(n_444),
.B2(n_447),
.C1(n_438),
.C2(n_445),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_469),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_459),
.B(n_442),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_473),
.A2(n_471),
.B(n_433),
.Y(n_477)
);

AOI322xp5_ASAP7_75t_L g475 ( 
.A1(n_472),
.A2(n_421),
.A3(n_447),
.B1(n_466),
.B2(n_438),
.C1(n_424),
.C2(n_403),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_476),
.Y(n_478)
);

AOI322xp5_ASAP7_75t_L g476 ( 
.A1(n_468),
.A2(n_421),
.A3(n_424),
.B1(n_408),
.B2(n_456),
.C1(n_355),
.C2(n_417),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_474),
.C(n_470),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_479),
.A2(n_480),
.B(n_453),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_478),
.B(n_451),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_409),
.Y(n_482)
);


endmodule