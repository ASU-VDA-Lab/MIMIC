module fake_netlist_6_1154_n_893 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_893);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_893;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_685;
wire n_832;
wire n_280;
wire n_287;
wire n_597;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_852;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_201;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_857;
wire n_674;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_SL g191 ( 
.A(n_135),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_52),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_45),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_43),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_1),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_35),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g205 ( 
.A(n_97),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_58),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_44),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_60),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_121),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_154),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_65),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_122),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_29),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_66),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_11),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_1),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_23),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_90),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_100),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_87),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_180),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_152),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_101),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_81),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_91),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_128),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_15),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_186),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_168),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_46),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_179),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_200),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_0),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_204),
.A2(n_21),
.B(n_20),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_204),
.B(n_22),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_2),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_191),
.B(n_3),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_193),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_206),
.B(n_4),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_219),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_195),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_222),
.B(n_25),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_223),
.A2(n_4),
.B(n_5),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_6),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_201),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_202),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_265),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_245),
.A2(n_7),
.B(n_9),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_211),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_212),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_9),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_292),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_194),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_R g322 ( 
.A(n_290),
.B(n_304),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_317),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_270),
.B(n_197),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_298),
.B(n_242),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_313),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_313),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_270),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_313),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_281),
.A2(n_279),
.B(n_306),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_315),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_315),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_315),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_276),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_R g345 ( 
.A(n_298),
.B(n_255),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_273),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_311),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_R g350 ( 
.A(n_316),
.B(n_213),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_318),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_214),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_276),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_309),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_301),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_215),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_294),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_294),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_288),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_288),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_270),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_270),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_271),
.Y(n_372)
);

AO221x1_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_316),
.B1(n_287),
.B2(n_308),
.C(n_307),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_271),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_287),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_287),
.Y(n_377)
);

NAND2xp33_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_274),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_271),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_271),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_283),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

AO21x2_ASAP7_75t_L g384 ( 
.A1(n_329),
.A2(n_275),
.B(n_302),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_321),
.B(n_282),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_289),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_321),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_341),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_293),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_305),
.Y(n_390)
);

OR2x6_ASAP7_75t_L g391 ( 
.A(n_319),
.B(n_267),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_345),
.B(n_336),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_328),
.B(n_268),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_277),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_L g398 ( 
.A1(n_343),
.A2(n_314),
.B1(n_272),
.B2(n_286),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_339),
.B(n_286),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_303),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_306),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_287),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_333),
.B(n_281),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_347),
.B(n_291),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_296),
.C(n_291),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_351),
.A2(n_300),
.B(n_316),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_291),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_354),
.A2(n_300),
.B1(n_217),
.B2(n_248),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_320),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_344),
.B(n_300),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_291),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_341),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_360),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_323),
.B(n_221),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_296),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_325),
.B(n_224),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_327),
.B(n_225),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_364),
.B(n_296),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_296),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_321),
.B(n_299),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_349),
.B(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_363),
.B(n_308),
.C(n_307),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_353),
.B(n_307),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_367),
.B(n_226),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_353),
.B(n_308),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_367),
.B(n_227),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_353),
.B(n_308),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_R g444 ( 
.A(n_415),
.B(n_228),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_277),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_229),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_382),
.Y(n_450)
);

OR2x2_ASAP7_75t_SL g451 ( 
.A(n_417),
.B(n_10),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_399),
.B(n_231),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_386),
.B(n_277),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_233),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_429),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_433),
.A2(n_277),
.B1(n_266),
.B2(n_262),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_398),
.A2(n_256),
.B1(n_239),
.B2(n_240),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

O2A1O1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_414),
.A2(n_277),
.B(n_260),
.C(n_259),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_234),
.Y(n_470)
);

O2A1O1Ixp5_ASAP7_75t_L g471 ( 
.A1(n_412),
.A2(n_253),
.B(n_252),
.C(n_251),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_385),
.B(n_241),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_403),
.B(n_243),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_434),
.A2(n_250),
.B(n_249),
.C(n_246),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_378),
.A2(n_98),
.B1(n_189),
.B2(n_188),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_389),
.B(n_11),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_390),
.B(n_12),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_394),
.B(n_12),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_373),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_427),
.B(n_13),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_371),
.B(n_14),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_405),
.B(n_26),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_391),
.B(n_16),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_410),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_431),
.B(n_372),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_440),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_391),
.B(n_16),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_396),
.B(n_27),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_416),
.B(n_30),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_431),
.B(n_17),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_412),
.B(n_31),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_409),
.B(n_374),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_395),
.B(n_17),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_32),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_431),
.B(n_34),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_395),
.A2(n_18),
.B1(n_19),
.B2(n_37),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_395),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_413),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_379),
.B(n_18),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_381),
.B(n_38),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_39),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_425),
.B(n_19),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_426),
.B(n_40),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_428),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_450),
.A2(n_388),
.B(n_421),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_494),
.A2(n_436),
.B1(n_441),
.B2(n_439),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_423),
.B1(n_442),
.B2(n_408),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_455),
.B(n_408),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_497),
.A2(n_424),
.B(n_384),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_497),
.A2(n_384),
.B1(n_50),
.B2(n_51),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_445),
.B(n_49),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_446),
.A2(n_53),
.B(n_54),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_489),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_446),
.A2(n_448),
.B(n_505),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_463),
.B(n_59),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_61),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_482),
.A2(n_62),
.B(n_63),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_471),
.A2(n_64),
.B(n_67),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_483),
.A2(n_490),
.B(n_487),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_461),
.B(n_68),
.Y(n_538)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_498),
.A2(n_69),
.B(n_70),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_470),
.B(n_393),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_488),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_477),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_444),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_513),
.A2(n_495),
.B1(n_473),
.B2(n_458),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_459),
.B(n_74),
.Y(n_546)
);

NOR3xp33_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_393),
.C(n_76),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_460),
.A2(n_75),
.B(n_77),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_466),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_449),
.B(n_78),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_462),
.B(n_79),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_468),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_456),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_502),
.B(n_85),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_506),
.B(n_88),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_485),
.A2(n_89),
.B(n_92),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_507),
.A2(n_94),
.B(n_95),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_500),
.B(n_96),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_491),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_454),
.B(n_99),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_105),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_478),
.A2(n_106),
.B(n_107),
.C(n_108),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_510),
.A2(n_110),
.B(n_112),
.Y(n_567)
);

O2A1O1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_474),
.A2(n_113),
.B(n_114),
.C(n_117),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_467),
.B(n_119),
.C(n_120),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_451),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_472),
.B(n_123),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_502),
.A2(n_480),
.B1(n_465),
.B2(n_503),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_512),
.A2(n_127),
.B(n_129),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_495),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_499),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_522),
.A2(n_514),
.B(n_501),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_529),
.A2(n_499),
.B(n_457),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_532),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_530),
.B(n_491),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_530),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_562),
.B(n_502),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_535),
.A2(n_453),
.B(n_457),
.Y(n_588)
);

BUFx2_ASAP7_75t_SL g589 ( 
.A(n_525),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_549),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_540),
.Y(n_592)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_520),
.A2(n_481),
.B(n_484),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_537),
.B(n_479),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_509),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_557),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_536),
.B(n_502),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_570),
.Y(n_598)
);

BUFx8_ASAP7_75t_SL g599 ( 
.A(n_544),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_519),
.Y(n_600)
);

AO21x2_ASAP7_75t_L g601 ( 
.A1(n_523),
.A2(n_493),
.B(n_469),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_509),
.Y(n_602)
);

NOR2xp67_ASAP7_75t_SL g603 ( 
.A(n_569),
.B(n_453),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_528),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_576),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_576),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_531),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_531),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_565),
.A2(n_475),
.B(n_515),
.Y(n_610)
);

NAND2x1p5_ASAP7_75t_L g611 ( 
.A(n_554),
.B(n_504),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_517),
.A2(n_504),
.B(n_138),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_524),
.A2(n_509),
.B(n_139),
.Y(n_613)
);

AO21x1_ASAP7_75t_L g614 ( 
.A1(n_572),
.A2(n_137),
.B(n_140),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_541),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_563),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_521),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_546),
.A2(n_142),
.B(n_145),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_545),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_551),
.A2(n_146),
.B(n_147),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_526),
.A2(n_568),
.B(n_548),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_550),
.B(n_190),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_534),
.A2(n_150),
.B(n_153),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_533),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_590),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_602),
.A2(n_575),
.B1(n_538),
.B2(n_518),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_613),
.A2(n_564),
.B1(n_571),
.B2(n_539),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_547),
.Y(n_631)
);

CKINVDCx14_ASAP7_75t_R g632 ( 
.A(n_579),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_580),
.Y(n_633)
);

NAND2x1_ASAP7_75t_L g634 ( 
.A(n_580),
.B(n_561),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_600),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_599),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_604),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_607),
.B(n_555),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_591),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_618),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_602),
.A2(n_527),
.B1(n_553),
.B2(n_559),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_618),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_603),
.A2(n_567),
.B(n_573),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_619),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_607),
.B(n_566),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_620),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_602),
.A2(n_543),
.B1(n_156),
.B2(n_158),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_581),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_607),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_625),
.B(n_155),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_581),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_605),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_599),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_608),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_605),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_592),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_606),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_602),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_594),
.A2(n_166),
.B(n_167),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_611),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_608),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_586),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_628),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_657),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

BUFx6f_ASAP7_75t_SL g674 ( 
.A(n_633),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_653),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_R g676 ( 
.A(n_632),
.B(n_579),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_SL g677 ( 
.A(n_657),
.B(n_615),
.C(n_621),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_653),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_637),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_646),
.B(n_635),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_635),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_637),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_640),
.B(n_595),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_638),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_665),
.B(n_627),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_631),
.B(n_586),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_632),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_660),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_667),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_668),
.B(n_595),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_648),
.B(n_596),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_652),
.B(n_586),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_SL g694 ( 
.A1(n_629),
.A2(n_627),
.B(n_614),
.C(n_593),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_666),
.B(n_586),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_633),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_630),
.A2(n_596),
.B1(n_589),
.B2(n_583),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_669),
.B(n_584),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_641),
.B(n_584),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_642),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_652),
.B(n_583),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_633),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_R g703 ( 
.A(n_647),
.B(n_585),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_650),
.B(n_583),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_649),
.A2(n_614),
.B1(n_625),
.B2(n_583),
.Y(n_705)
);

AND3x1_ASAP7_75t_L g706 ( 
.A(n_663),
.B(n_615),
.C(n_616),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_659),
.Y(n_707)
);

INVx4_ASAP7_75t_SL g708 ( 
.A(n_633),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_644),
.B(n_617),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_654),
.B(n_617),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_654),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_656),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_647),
.B(n_615),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_639),
.B(n_580),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_634),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_656),
.B(n_585),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_639),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_662),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_662),
.B(n_580),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_717),
.B(n_683),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_722),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_675),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_671),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_612),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_717),
.B(n_612),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_686),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_686),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_707),
.B(n_670),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_686),
.Y(n_732)
);

AND2x4_ASAP7_75t_SL g733 ( 
.A(n_680),
.B(n_585),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_704),
.B(n_587),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_675),
.Y(n_735)
);

AOI211xp5_ASAP7_75t_L g736 ( 
.A1(n_697),
.A2(n_658),
.B(n_626),
.C(n_624),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_673),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_700),
.B(n_670),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_687),
.B(n_623),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_678),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_685),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_718),
.B(n_664),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_711),
.B(n_664),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_711),
.B(n_623),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_719),
.Y(n_745)
);

AOI33xp33_ASAP7_75t_L g746 ( 
.A1(n_691),
.A2(n_643),
.A3(n_601),
.B1(n_645),
.B2(n_626),
.B3(n_176),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_719),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_712),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_720),
.B(n_601),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_681),
.B(n_588),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_721),
.B(n_587),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_715),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_709),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_684),
.B(n_588),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_686),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_689),
.B(n_577),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_710),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_701),
.B(n_587),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_716),
.B(n_587),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_716),
.B(n_610),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_749),
.B(n_713),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_749),
.B(n_713),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_757),
.B(n_690),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_726),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_756),
.B(n_753),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_756),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_724),
.B(n_692),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_750),
.B(n_693),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_723),
.B(n_737),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_738),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_741),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_677),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_731),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_715),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_750),
.B(n_688),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_738),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_748),
.B(n_695),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_754),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_761),
.B(n_708),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_754),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_734),
.B(n_695),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_725),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_761),
.B(n_696),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_735),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_734),
.B(n_699),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_742),
.B(n_702),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_742),
.B(n_705),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_727),
.B(n_714),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_785),
.B(n_758),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_779),
.B(n_739),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_771),
.B(n_727),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_771),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_781),
.B(n_767),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_772),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_777),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_766),
.B(n_743),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_770),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_783),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_785),
.B(n_758),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_784),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_788),
.B(n_728),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_SL g806 ( 
.A(n_773),
.B(n_736),
.C(n_746),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_788),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_776),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_786),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_806),
.A2(n_706),
.B1(n_789),
.B2(n_703),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_806),
.A2(n_789),
.B(n_688),
.C(n_762),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_792),
.B(n_729),
.Y(n_812)
);

AOI32xp33_ASAP7_75t_L g813 ( 
.A1(n_808),
.A2(n_762),
.A3(n_763),
.B1(n_790),
.B2(n_775),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_795),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_801),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_798),
.B(n_764),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_796),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_795),
.Y(n_818)
);

OAI22xp33_ASAP7_75t_L g819 ( 
.A1(n_798),
.A2(n_703),
.B1(n_729),
.B2(n_755),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_797),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_810),
.A2(n_763),
.B1(n_780),
.B2(n_734),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_816),
.Y(n_822)
);

XOR2x2_ASAP7_75t_L g823 ( 
.A(n_817),
.B(n_679),
.Y(n_823)
);

NOR4xp25_ASAP7_75t_L g824 ( 
.A(n_811),
.B(n_778),
.C(n_796),
.D(n_799),
.Y(n_824)
);

XNOR2xp5_ASAP7_75t_L g825 ( 
.A(n_819),
.B(n_679),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_814),
.A2(n_820),
.B(n_818),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_812),
.A2(n_729),
.B1(n_755),
.B2(n_800),
.Y(n_827)
);

OAI21xp33_ASAP7_75t_L g828 ( 
.A1(n_824),
.A2(n_813),
.B(n_815),
.Y(n_828)
);

OAI322xp33_ASAP7_75t_L g829 ( 
.A1(n_825),
.A2(n_800),
.A3(n_774),
.B1(n_804),
.B2(n_797),
.C1(n_768),
.C2(n_769),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_821),
.A2(n_812),
.B1(n_755),
.B2(n_729),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_822),
.A2(n_729),
.B1(n_755),
.B2(n_807),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_823),
.B(n_791),
.Y(n_832)
);

AO22x2_ASAP7_75t_L g833 ( 
.A1(n_826),
.A2(n_794),
.B1(n_809),
.B2(n_802),
.Y(n_833)
);

NAND2x1_ASAP7_75t_L g834 ( 
.A(n_827),
.B(n_793),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_828),
.B(n_803),
.Y(n_835)
);

NAND4xp25_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_782),
.C(n_787),
.D(n_790),
.Y(n_836)
);

AOI221x1_ASAP7_75t_L g837 ( 
.A1(n_833),
.A2(n_794),
.B1(n_805),
.B2(n_752),
.C(n_760),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_834),
.Y(n_838)
);

AOI22x1_ASAP7_75t_SL g839 ( 
.A1(n_829),
.A2(n_682),
.B1(n_672),
.B2(n_676),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_835),
.B(n_831),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_SL g841 ( 
.A1(n_838),
.A2(n_830),
.B(n_780),
.Y(n_841)
);

AND3x1_ASAP7_75t_L g842 ( 
.A(n_840),
.B(n_839),
.C(n_836),
.Y(n_842)
);

AOI211xp5_ASAP7_75t_L g843 ( 
.A1(n_841),
.A2(n_676),
.B(n_682),
.C(n_672),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_SL g844 ( 
.A(n_840),
.B(n_714),
.C(n_837),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_844),
.B(n_805),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_842),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_843),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_842),
.B(n_793),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_844),
.B(n_780),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_842),
.Y(n_850)
);

NAND4xp75_ASAP7_75t_L g851 ( 
.A(n_846),
.B(n_698),
.C(n_728),
.D(n_775),
.Y(n_851)
);

NAND4xp75_ASAP7_75t_L g852 ( 
.A(n_850),
.B(n_759),
.C(n_743),
.D(n_744),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_SL g853 ( 
.A1(n_847),
.A2(n_733),
.B(n_739),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_849),
.B(n_733),
.Y(n_854)
);

AND3x4_ASAP7_75t_L g855 ( 
.A(n_845),
.B(n_848),
.C(n_751),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_846),
.B(n_694),
.C(n_760),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_856),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_853),
.B(n_735),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_854),
.B(n_755),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_851),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_852),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_862),
.A2(n_730),
.B1(n_732),
.B2(n_752),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_858),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_861),
.Y(n_866)
);

XNOR2x2_ASAP7_75t_L g867 ( 
.A(n_857),
.B(n_610),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_859),
.Y(n_868)
);

XNOR2x1_ASAP7_75t_L g869 ( 
.A(n_860),
.B(n_169),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_860),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_862),
.A2(n_674),
.B1(n_751),
.B2(n_686),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_861),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_866),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_872),
.Y(n_874)
);

AOI31xp33_ASAP7_75t_L g875 ( 
.A1(n_869),
.A2(n_597),
.A3(n_708),
.B(n_674),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_863),
.B(n_686),
.Y(n_876)
);

OAI31xp33_ASAP7_75t_SL g877 ( 
.A1(n_870),
.A2(n_708),
.A3(n_759),
.B(n_674),
.Y(n_877)
);

OAI22xp33_ASAP7_75t_L g878 ( 
.A1(n_868),
.A2(n_732),
.B1(n_730),
.B2(n_745),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_868),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_865),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_867),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_879),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_873),
.A2(n_871),
.B1(n_864),
.B2(n_730),
.Y(n_883)
);

OAI22x1_ASAP7_75t_L g884 ( 
.A1(n_874),
.A2(n_732),
.B1(n_597),
.B2(n_751),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_880),
.Y(n_885)
);

AO22x2_ASAP7_75t_L g886 ( 
.A1(n_881),
.A2(n_747),
.B1(n_745),
.B2(n_740),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_875),
.B(n_171),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_882),
.A2(n_877),
.B(n_876),
.Y(n_888)
);

OAI22x1_ASAP7_75t_L g889 ( 
.A1(n_885),
.A2(n_878),
.B1(n_747),
.B2(n_740),
.Y(n_889)
);

XNOR2xp5_ASAP7_75t_L g890 ( 
.A(n_888),
.B(n_887),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_890),
.A2(n_883),
.B1(n_886),
.B2(n_884),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_891),
.B(n_889),
.Y(n_892)
);

AOI211xp5_ASAP7_75t_L g893 ( 
.A1(n_892),
.A2(n_172),
.B(n_173),
.C(n_178),
.Y(n_893)
);


endmodule