module fake_jpeg_10484_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_25),
.B1(n_13),
.B2(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_12),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_57),
.B(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_29),
.C(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_72),
.B1(n_79),
.B2(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_15),
.B1(n_13),
.B2(n_29),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_54),
.B1(n_55),
.B2(n_15),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_87),
.B1(n_95),
.B2(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_63),
.B1(n_66),
.B2(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_48),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_75),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_24),
.B(n_2),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_83),
.C(n_77),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_105),
.B1(n_91),
.B2(n_96),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_75),
.C(n_46),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_109),
.C(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

OAI322xp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_94),
.A3(n_89),
.B1(n_92),
.B2(n_87),
.C1(n_85),
.C2(n_99),
.Y(n_114)
);

OA21x2_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_86),
.B(n_23),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_5),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.C(n_109),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_50),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_102),
.B1(n_100),
.B2(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.C(n_80),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_6),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_126),
.B1(n_133),
.B2(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_3),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_9),
.B(n_10),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_9),
.C(n_3),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.C(n_134),
.Y(n_141)
);


endmodule