module fake_jpeg_15425_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_45),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_54),
.Y(n_96)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_21),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_8),
.Y(n_114)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_29),
.B1(n_32),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_87),
.B1(n_98),
.B2(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_86),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_29),
.B1(n_32),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_73),
.A2(n_83),
.B1(n_85),
.B2(n_48),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_79),
.A2(n_94),
.B1(n_33),
.B2(n_30),
.Y(n_135)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_47),
.B1(n_55),
.B2(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_16),
.C(n_28),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_11),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_22),
.B1(n_33),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_41),
.B(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_89),
.B(n_100),
.Y(n_149)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_16),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_9),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_48),
.A2(n_9),
.B1(n_13),
.B2(n_11),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_8),
.Y(n_157)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_11),
.Y(n_118)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_160),
.B1(n_105),
.B2(n_72),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_63),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_59),
.B(n_56),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_127),
.A2(n_150),
.B(n_107),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_131),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_134),
.A2(n_142),
.B(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_137),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_71),
.B(n_16),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_143),
.Y(n_176)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_51),
.B(n_42),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_51),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_68),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_146),
.B(n_147),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_69),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_80),
.A2(n_91),
.B1(n_101),
.B2(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_167),
.B1(n_108),
.B2(n_104),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_77),
.B(n_10),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_69),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_154),
.B(n_157),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_114),
.B(n_96),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_10),
.B1(n_8),
.B2(n_45),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_161),
.B1(n_109),
.B2(n_108),
.Y(n_174)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_44),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

AO22x2_ASAP7_75t_L g161 ( 
.A1(n_87),
.A2(n_45),
.B1(n_44),
.B2(n_2),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_0),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_0),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_1),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_72),
.C(n_82),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_187),
.C(n_208),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_174),
.A2(n_184),
.B1(n_182),
.B2(n_211),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_189),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_193),
.B(n_195),
.Y(n_233)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_107),
.B1(n_115),
.B2(n_111),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_191),
.B1(n_195),
.B2(n_216),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_184),
.A2(n_204),
.B1(n_133),
.B2(n_153),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_72),
.C(n_82),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_104),
.B1(n_97),
.B2(n_75),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_97),
.B1(n_75),
.B2(n_105),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_1),
.B(n_3),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_198),
.B(n_203),
.Y(n_224)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_88),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_161),
.A2(n_88),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_143),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_4),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_209),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_131),
.B(n_6),
.C(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_4),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_200),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_128),
.A2(n_5),
.B1(n_124),
.B2(n_120),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_162),
.B1(n_5),
.B2(n_157),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_127),
.A2(n_5),
.B1(n_125),
.B2(n_167),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_123),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_217),
.B(n_232),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_125),
.B1(n_150),
.B2(n_152),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_218),
.A2(n_221),
.B1(n_226),
.B2(n_229),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_123),
.B1(n_122),
.B2(n_124),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_220),
.A2(n_228),
.B(n_238),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_169),
.B1(n_129),
.B2(n_130),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_168),
.B(n_164),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_225),
.A2(n_233),
.B(n_242),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_129),
.B1(n_130),
.B2(n_136),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_132),
.B1(n_151),
.B2(n_144),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_136),
.B1(n_140),
.B2(n_148),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_192),
.B(n_132),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_241),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_183),
.B(n_144),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_234),
.B(n_248),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_239),
.B1(n_226),
.B2(n_220),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_149),
.C(n_148),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_249),
.C(n_208),
.Y(n_268)
);

AOI32xp33_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_133),
.A3(n_147),
.B1(n_154),
.B2(n_149),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_186),
.A2(n_139),
.B1(n_158),
.B2(n_140),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_5),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_162),
.B(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_194),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_176),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_253),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_172),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_176),
.B(n_173),
.C(n_187),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_202),
.A2(n_191),
.B(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_188),
.B(n_200),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_197),
.A2(n_213),
.B(n_196),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_199),
.B(n_213),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_177),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_178),
.B(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_174),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_259),
.A2(n_254),
.B(n_258),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_178),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_282),
.Y(n_307)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_268),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_206),
.B1(n_171),
.B2(n_190),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_263),
.A2(n_266),
.B1(n_289),
.B2(n_221),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_265),
.B(n_269),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_219),
.A2(n_171),
.B1(n_190),
.B2(n_186),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_288),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_177),
.A3(n_180),
.B1(n_194),
.B2(n_201),
.C1(n_230),
.C2(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_201),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_279),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_244),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_252),
.B1(n_250),
.B2(n_225),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_222),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_237),
.C(n_247),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_287),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_235),
.A2(n_233),
.B1(n_218),
.B2(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_245),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_248),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_242),
.C(n_227),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_228),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_304),
.B1(n_308),
.B2(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_293),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_312),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_284),
.B(n_259),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_301),
.A2(n_302),
.B(n_305),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_224),
.B(n_255),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_300),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_225),
.B1(n_244),
.B2(n_256),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_253),
.B1(n_257),
.B2(n_227),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_311),
.C(n_321),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_241),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_280),
.A2(n_259),
.B1(n_265),
.B2(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_222),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_317),
.B(n_277),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_274),
.A2(n_229),
.B1(n_239),
.B2(n_232),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_295),
.B1(n_304),
.B2(n_308),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_263),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_319),
.A2(n_320),
.B(n_303),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_286),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_268),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_281),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_342),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_276),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_328),
.C(n_341),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_289),
.B1(n_271),
.B2(n_278),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_327),
.B1(n_329),
.B2(n_330),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_260),
.B1(n_281),
.B2(n_280),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_282),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_291),
.B1(n_288),
.B2(n_272),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_296),
.A2(n_291),
.B1(n_272),
.B2(n_264),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_301),
.A2(n_264),
.B1(n_287),
.B2(n_283),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_331),
.A2(n_314),
.B1(n_294),
.B2(n_298),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_302),
.B(n_270),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_297),
.C(n_337),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_334),
.B(n_313),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_336),
.A2(n_338),
.B1(n_299),
.B2(n_310),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_270),
.B1(n_277),
.B2(n_293),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_337),
.B(n_324),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_340),
.A2(n_305),
.B1(n_300),
.B2(n_294),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_307),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_311),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_297),
.C(n_333),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_309),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_348),
.C(n_356),
.Y(n_362)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_338),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_354),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_347),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_306),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_350),
.A2(n_360),
.B1(n_354),
.B2(n_344),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_355),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_329),
.B(n_310),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_353),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_357),
.A2(n_360),
.B1(n_326),
.B2(n_340),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_342),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_358),
.A2(n_359),
.B(n_330),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_343),
.C(n_333),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_367),
.C(n_368),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_361),
.Y(n_365)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_323),
.C(n_327),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_339),
.C(n_332),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_349),
.B(n_355),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_371),
.A2(n_349),
.B1(n_357),
.B2(n_326),
.Y(n_380)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_345),
.C(n_352),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_380),
.C(n_367),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_371),
.B(n_373),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_381),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_383),
.A2(n_384),
.B(n_366),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_387),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_382),
.A2(n_379),
.B(n_375),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_372),
.B(n_369),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_389),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_390),
.B(n_388),
.Y(n_391)
);

AOI321xp33_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_376),
.A3(n_380),
.B1(n_378),
.B2(n_374),
.C(n_362),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_392),
.A2(n_376),
.B(n_368),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_364),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_348),
.Y(n_395)
);


endmodule