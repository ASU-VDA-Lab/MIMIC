module fake_jpeg_2777_n_193 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_20),
.B1(n_23),
.B2(n_27),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_79),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_20),
.B1(n_27),
.B2(n_23),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_63),
.B1(n_75),
.B2(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_28),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_19),
.C(n_15),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_82),
.C(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_29),
.B1(n_30),
.B2(n_19),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_44),
.B1(n_42),
.B2(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_22),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_2),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_48),
.B1(n_49),
.B2(n_25),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_70),
.B1(n_58),
.B2(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_1),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_65),
.B1(n_77),
.B2(n_51),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_77),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_93),
.B1(n_97),
.B2(n_101),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_25),
.C(n_4),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_25),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

OAI22x1_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_67),
.B1(n_65),
.B2(n_59),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_113),
.B1(n_53),
.B2(n_54),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_93),
.B1(n_88),
.B2(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_51),
.B(n_74),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_100),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_9),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_84),
.B1(n_102),
.B2(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_66),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_134),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_145),
.B(n_131),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_117),
.B(n_122),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_92),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_141),
.C(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_94),
.B1(n_72),
.B2(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_137),
.B1(n_127),
.B2(n_124),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_72),
.B1(n_103),
.B2(n_77),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_10),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_53),
.C(n_54),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_144),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_13),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_115),
.C(n_114),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_141),
.C(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_138),
.B(n_119),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_144),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_122),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_143),
.C(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_130),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_150),
.C(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_169),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_159),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_164),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_152),
.B1(n_128),
.B2(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_7),
.B1(n_123),
.B2(n_171),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_166),
.CI(n_7),
.CON(n_179),
.SN(n_179)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_180),
.B1(n_172),
.B2(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_173),
.C(n_176),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.C(n_176),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_178),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_184),
.C(n_183),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_190),
.B1(n_179),
.B2(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_179),
.C(n_7),
.Y(n_193)
);


endmodule