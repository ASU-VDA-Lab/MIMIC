module fake_jpeg_15045_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_1),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_61),
.Y(n_84)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_48),
.Y(n_103)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_43),
.B1(n_41),
.B2(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_42),
.B1(n_78),
.B2(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_2),
.Y(n_98)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_94),
.B1(n_100),
.B2(n_102),
.Y(n_110)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_53),
.Y(n_94)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_106),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_60),
.B1(n_61),
.B2(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_52),
.B1(n_44),
.B2(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_48),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_46),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_45),
.B1(n_55),
.B2(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_114),
.B1(n_119),
.B2(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_22),
.B1(n_39),
.B2(n_38),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_123),
.B1(n_125),
.B2(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_115),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_129),
.B1(n_111),
.B2(n_105),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_103),
.B(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_110),
.B1(n_126),
.B2(n_114),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_134),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_2),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_5),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_132),
.C(n_9),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_138),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_26),
.C(n_11),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_27),
.B(n_12),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_29),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_19),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_30),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_18),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_31),
.B(n_13),
.C(n_14),
.Y(n_153)
);


endmodule