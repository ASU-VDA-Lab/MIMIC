module fake_jpeg_17781_n_354 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_38),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_68),
.B1(n_67),
.B2(n_54),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_45),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_19),
.B1(n_27),
.B2(n_40),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_19),
.B1(n_27),
.B2(n_33),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_34),
.B1(n_25),
.B2(n_31),
.Y(n_87)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_36),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_18),
.C(n_22),
.Y(n_112)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_0),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_29),
.B(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_30),
.B(n_35),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

BUFx2_ASAP7_75t_SL g109 ( 
.A(n_91),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_130),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_101),
.Y(n_137)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_133),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_121),
.B(n_47),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_0),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_98),
.B1(n_104),
.B2(n_82),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_90),
.Y(n_154)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_77),
.C(n_42),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_45),
.C(n_42),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_104),
.B1(n_88),
.B2(n_91),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_76),
.B1(n_61),
.B2(n_36),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_134),
.B1(n_88),
.B2(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_41),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_76),
.B1(n_46),
.B2(n_41),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_57),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_45),
.B1(n_42),
.B2(n_49),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_100),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_134),
.C(n_117),
.Y(n_176)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_143),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_93),
.B(n_94),
.C(n_101),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_151),
.B(n_35),
.Y(n_186)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_49),
.B1(n_44),
.B2(n_47),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_99),
.B1(n_92),
.B2(n_79),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_90),
.B(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_157),
.B(n_161),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_113),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_102),
.B1(n_89),
.B2(n_75),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_162),
.B1(n_132),
.B2(n_120),
.Y(n_166)
);

OR2x6_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_89),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_75),
.B1(n_100),
.B2(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_130),
.B(n_106),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_171),
.B(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_140),
.B1(n_160),
.B2(n_150),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_146),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_118),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_184),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_127),
.C(n_112),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_189),
.C(n_156),
.Y(n_210)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_129),
.B1(n_115),
.B2(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_117),
.C(n_77),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_120),
.B(n_113),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_152),
.B1(n_163),
.B2(n_158),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_135),
.C(n_103),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_135),
.C(n_103),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_148),
.B(n_151),
.Y(n_202)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_202),
.B(n_186),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_164),
.B(n_141),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_206),
.C(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_204),
.B1(n_211),
.B2(n_114),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_178),
.B1(n_182),
.B2(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

OR2x2_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_176),
.B1(n_174),
.B2(n_166),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_145),
.B1(n_162),
.B2(n_152),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_24),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_136),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_35),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_178),
.B1(n_174),
.B2(n_182),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_220),
.B(n_234),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_238),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_177),
.B1(n_183),
.B2(n_187),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_165),
.B1(n_175),
.B2(n_116),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_233),
.B1(n_237),
.B2(n_244),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.C(n_240),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_155),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_125),
.B1(n_24),
.B2(n_23),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_11),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_105),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_105),
.C(n_22),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_0),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_257),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_210),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_250),
.B(n_30),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_255),
.C(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_191),
.C(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_197),
.C(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_235),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_263),
.C(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_197),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_196),
.C(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_199),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_201),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_22),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_244),
.B1(n_233),
.B2(n_224),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_23),
.B1(n_21),
.B2(n_4),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_219),
.CI(n_244),
.CON(n_270),
.SN(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_227),
.B1(n_219),
.B2(n_196),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_282),
.B1(n_280),
.B2(n_261),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_219),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_275),
.C(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_212),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_251),
.B(n_13),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_263),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_24),
.C(n_23),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_287),
.C(n_264),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_24),
.C(n_23),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_292),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_262),
.B(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_280),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_250),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_262),
.B1(n_264),
.B2(n_3),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_286),
.B1(n_271),
.B2(n_287),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_22),
.C(n_18),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_1),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_22),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_22),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.C(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_2),
.C(n_3),
.Y(n_304)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_314),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_268),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_316),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_310),
.B1(n_5),
.B2(n_6),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_285),
.C(n_4),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_315),
.C(n_288),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_16),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_14),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_291),
.A2(n_295),
.B1(n_301),
.B2(n_302),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_2),
.C(n_4),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_16),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_296),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_292),
.B(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_14),
.B(n_13),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_331),
.B(n_7),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_311),
.B(n_308),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_5),
.C(n_6),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_330),
.C(n_315),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_8),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_5),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_7),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_321),
.A2(n_328),
.B(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_333),
.A2(n_326),
.B(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_336),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_338),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_310),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_340),
.B(n_327),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g340 ( 
.A1(n_325),
.A2(n_319),
.B(n_9),
.C(n_10),
.Y(n_340)
);

AO21x2_ASAP7_75t_L g349 ( 
.A1(n_341),
.A2(n_345),
.B(n_332),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_344),
.B(n_346),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_8),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_8),
.B(n_9),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_342),
.C(n_349),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_347),
.C(n_9),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_10),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_353),
.Y(n_354)
);


endmodule