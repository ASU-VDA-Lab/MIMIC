module fake_jpeg_28_n_227 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_56),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_78),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

BUFx6f_ASAP7_75t_SL g88 ( 
.A(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_60),
.B1(n_64),
.B2(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_77),
.B1(n_59),
.B2(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_66),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_87),
.B1(n_80),
.B2(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_84),
.B1(n_80),
.B2(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_93),
.Y(n_109)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_115),
.B1(n_97),
.B2(n_70),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_88),
.B1(n_61),
.B2(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_121),
.B1(n_63),
.B2(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_96),
.C(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_54),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_55),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_69),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_119),
.B(n_76),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_77),
.B1(n_73),
.B2(n_75),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_125),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_128),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_62),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_136),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_25),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_24),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_8),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_103),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_115),
.B1(n_116),
.B2(n_105),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_30),
.B1(n_50),
.B2(n_48),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_1),
.B(n_4),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_163),
.B(n_11),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_6),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_8),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_10),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_11),
.B(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_10),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_137),
.B1(n_13),
.B2(n_14),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_187),
.B1(n_149),
.B2(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_151),
.B1(n_147),
.B2(n_156),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_29),
.B(n_47),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_176),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_35),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_184),
.C(n_161),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_27),
.B(n_46),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_26),
.C(n_44),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_161),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_52),
.B(n_23),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_148),
.B1(n_162),
.B2(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_185),
.A3(n_183),
.B1(n_181),
.B2(n_179),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_171),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_187),
.B1(n_174),
.B2(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_200),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_199),
.C(n_198),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.C(n_172),
.Y(n_200)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_175),
.B1(n_180),
.B2(n_173),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_184),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_21),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_191),
.B1(n_36),
.B2(n_17),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_15),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_213),
.B1(n_219),
.B2(n_211),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_201),
.B(n_210),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_218),
.A3(n_202),
.B1(n_212),
.B2(n_20),
.C1(n_38),
.C2(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_15),
.B(n_16),
.C(n_19),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_40),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_42),
.Y(n_227)
);


endmodule