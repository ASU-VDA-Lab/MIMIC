module real_aes_8679_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_635;
wire n_905;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_638;
wire n_519;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_938;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_960;
wire n_973;
wire n_504;
wire n_671;
wire n_725;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_0), .A2(n_171), .B1(n_959), .B2(n_960), .Y(n_958) );
INVx1_ASAP7_75t_L g825 ( .A(n_1), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_2), .A2(n_216), .B1(n_401), .B2(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_3), .A2(n_162), .B1(n_297), .B2(n_431), .C1(n_455), .C2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_4), .A2(n_228), .B1(n_501), .B2(n_557), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_5), .A2(n_97), .B1(n_354), .B2(n_370), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_6), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_7), .A2(n_147), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_8), .A2(n_86), .B1(n_485), .B2(n_488), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_9), .A2(n_70), .B1(n_431), .B2(n_689), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_10), .B(n_533), .Y(n_532) );
AO22x2_ASAP7_75t_L g369 ( .A1(n_11), .A2(n_199), .B1(n_360), .B2(n_365), .Y(n_369) );
INVx1_ASAP7_75t_L g985 ( .A(n_11), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_12), .A2(n_156), .B1(n_498), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_13), .A2(n_318), .B1(n_452), .B2(n_611), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_14), .A2(n_143), .B1(n_372), .B2(n_544), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_15), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_16), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_17), .A2(n_177), .B1(n_410), .B2(n_506), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_18), .A2(n_224), .B1(n_372), .B2(n_514), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_19), .A2(n_285), .B1(n_390), .B2(n_393), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_20), .A2(n_286), .B1(n_480), .B2(n_737), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g517 ( .A1(n_21), .A2(n_57), .B1(n_249), .B2(n_452), .C1(n_518), .C2(n_520), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_22), .A2(n_274), .B1(n_605), .B2(n_891), .Y(n_890) );
AOI22xp5_ASAP7_75t_SL g853 ( .A1(n_23), .A2(n_221), .B1(n_544), .B2(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_24), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_25), .A2(n_272), .B1(n_370), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_26), .A2(n_227), .B1(n_557), .B2(n_603), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_27), .A2(n_322), .B1(n_516), .B2(n_540), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_28), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_29), .A2(n_219), .B1(n_488), .B2(n_498), .Y(n_668) );
AO22x2_ASAP7_75t_L g367 ( .A1(n_30), .A2(n_112), .B1(n_360), .B2(n_361), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_31), .A2(n_159), .B1(n_384), .B2(n_402), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_32), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_33), .A2(n_945), .B1(n_966), .B2(n_967), .Y(n_944) );
INVx1_ASAP7_75t_L g967 ( .A(n_33), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_34), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_35), .A2(n_53), .B1(n_479), .B2(n_603), .Y(n_671) );
INVx1_ASAP7_75t_L g803 ( .A(n_36), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_37), .A2(n_259), .B1(n_431), .B2(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_38), .A2(n_54), .B1(n_356), .B2(n_597), .Y(n_772) );
INVx1_ASAP7_75t_L g577 ( .A(n_39), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_40), .A2(n_151), .B1(n_498), .B2(n_911), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_41), .A2(n_269), .B1(n_354), .B2(n_401), .Y(n_964) );
INVx1_ASAP7_75t_L g998 ( .A(n_42), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_43), .A2(n_191), .B1(n_420), .B2(n_432), .Y(n_801) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_44), .A2(n_266), .B1(n_284), .B2(n_424), .C1(n_426), .C2(n_430), .Y(n_423) );
AOI22xp5_ASAP7_75t_SL g852 ( .A1(n_45), .A2(n_281), .B1(n_501), .B2(n_692), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_46), .Y(n_615) );
AOI22xp5_ASAP7_75t_SL g771 ( .A1(n_47), .A2(n_198), .B1(n_372), .B2(n_692), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_48), .A2(n_64), .B1(n_585), .B2(n_877), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_49), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_50), .A2(n_292), .B1(n_508), .B2(n_509), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g918 ( .A(n_51), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_52), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_55), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_56), .A2(n_220), .B1(n_572), .B2(n_648), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_58), .A2(n_85), .B1(n_431), .B2(n_509), .Y(n_999) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_59), .A2(n_121), .B1(n_512), .B2(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g823 ( .A(n_60), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g812 ( .A(n_61), .B(n_777), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_62), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_63), .A2(n_185), .B1(n_648), .B2(n_650), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_65), .A2(n_84), .B1(n_644), .B2(n_646), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_66), .A2(n_196), .B1(n_410), .B2(n_414), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_67), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_68), .A2(n_206), .B1(n_474), .B2(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g635 ( .A(n_69), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_71), .A2(n_204), .B1(n_502), .B2(n_775), .Y(n_848) );
AOI22xp5_ASAP7_75t_SL g774 ( .A1(n_72), .A2(n_91), .B1(n_488), .B2(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g587 ( .A(n_73), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_74), .A2(n_142), .B1(n_570), .B2(n_572), .Y(n_569) );
AO22x2_ASAP7_75t_L g364 ( .A1(n_75), .A2(n_231), .B1(n_360), .B2(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g982 ( .A(n_75), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_240), .B1(n_384), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_77), .A2(n_78), .B1(n_644), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_79), .A2(n_313), .B1(n_520), .B2(n_581), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_80), .A2(n_311), .B1(n_499), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_81), .A2(n_262), .B1(n_413), .B2(n_505), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g949 ( .A1(n_82), .A2(n_194), .B1(n_430), .B2(n_950), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_83), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_87), .A2(n_257), .B1(n_478), .B2(n_480), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_88), .A2(n_276), .B1(n_537), .B2(n_597), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g988 ( .A1(n_89), .A2(n_989), .B1(n_990), .B2(n_1007), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_89), .Y(n_1007) );
OA22x2_ASAP7_75t_L g349 ( .A1(n_90), .A2(n_350), .B1(n_351), .B2(n_434), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_90), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_92), .A2(n_186), .B1(n_401), .B2(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g1003 ( .A1(n_93), .A2(n_108), .B1(n_488), .B2(n_512), .Y(n_1003) );
INVx1_ASAP7_75t_L g575 ( .A(n_94), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_95), .A2(n_102), .B1(n_426), .B2(n_611), .Y(n_664) );
INVx1_ASAP7_75t_L g768 ( .A(n_96), .Y(n_768) );
INVx1_ASAP7_75t_L g558 ( .A(n_98), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_99), .A2(n_120), .B1(n_487), .B2(n_962), .Y(n_961) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_100), .A2(n_336), .B(n_344), .C(n_987), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_101), .A2(n_145), .B1(n_416), .B2(n_838), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_103), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_104), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_105), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_106), .B(n_994), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_107), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_109), .A2(n_248), .B1(n_502), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g564 ( .A(n_110), .Y(n_564) );
INVx1_ASAP7_75t_L g687 ( .A(n_111), .Y(n_687) );
INVx1_ASAP7_75t_L g986 ( .A(n_112), .Y(n_986) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_113), .A2(n_132), .B1(n_379), .B2(n_480), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_114), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_115), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_116), .A2(n_183), .B1(n_417), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_117), .A2(n_123), .B1(n_401), .B2(n_694), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_118), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_119), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_119), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_122), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_124), .Y(n_748) );
AOI211xp5_ASAP7_75t_L g920 ( .A1(n_125), .A2(n_424), .B(n_921), .C(n_927), .Y(n_920) );
INVx1_ASAP7_75t_L g697 ( .A(n_126), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_127), .Y(n_808) );
INVx1_ASAP7_75t_L g1015 ( .A(n_128), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_129), .A2(n_299), .B1(n_399), .B2(n_404), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_130), .A2(n_158), .B1(n_512), .B2(n_598), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_131), .A2(n_230), .B1(n_585), .B2(n_612), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_133), .A2(n_320), .B1(n_452), .B2(n_611), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_134), .A2(n_553), .B1(n_591), .B2(n_592), .Y(n_552) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_134), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_135), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_136), .A2(n_236), .B1(n_393), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_137), .A2(n_168), .B1(n_384), .B2(n_479), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_138), .A2(n_319), .B1(n_416), .B2(n_838), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_139), .A2(n_243), .B1(n_416), .B2(n_420), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_140), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_141), .A2(n_210), .B1(n_478), .B2(n_572), .Y(n_965) );
AND2x6_ASAP7_75t_L g338 ( .A(n_144), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_144), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_146), .A2(n_271), .B1(n_401), .B2(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_148), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_149), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_150), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_152), .A2(n_315), .B1(n_479), .B2(n_886), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_153), .A2(n_215), .B1(n_420), .B2(n_431), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_154), .A2(n_325), .B1(n_488), .B2(n_498), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_155), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_157), .A2(n_239), .B1(n_379), .B2(n_383), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_160), .A2(n_331), .B1(n_458), .B2(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g639 ( .A(n_161), .Y(n_639) );
INVx1_ASAP7_75t_L g582 ( .A(n_163), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_164), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_165), .A2(n_169), .B1(n_605), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_166), .A2(n_238), .B1(n_390), .B2(n_889), .Y(n_888) );
AO22x2_ASAP7_75t_L g359 ( .A1(n_167), .A2(n_222), .B1(n_360), .B2(n_361), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_167), .B(n_984), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_170), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_172), .A2(n_237), .B1(n_501), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_173), .A2(n_225), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_174), .A2(n_273), .B1(n_585), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_175), .A2(n_309), .B1(n_372), .B2(n_598), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_176), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_178), .A2(n_334), .B1(n_452), .B2(n_585), .Y(n_636) );
INVx1_ASAP7_75t_L g630 ( .A(n_179), .Y(n_630) );
INVx1_ASAP7_75t_L g638 ( .A(n_180), .Y(n_638) );
AOI22xp5_ASAP7_75t_SL g856 ( .A1(n_181), .A2(n_245), .B1(n_562), .B2(n_777), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_182), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_184), .A2(n_213), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_187), .A2(n_304), .B1(n_384), .B2(n_399), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_188), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_189), .B(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_190), .A2(n_729), .B1(n_764), .B2(n_765), .Y(n_728) );
INVx1_ASAP7_75t_L g764 ( .A(n_190), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_192), .A2(n_223), .B1(n_416), .B2(n_838), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_193), .A2(n_327), .B1(n_354), .B2(n_692), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_195), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_197), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_200), .A2(n_439), .B1(n_489), .B2(n_490), .Y(n_438) );
INVx1_ASAP7_75t_L g489 ( .A(n_200), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_201), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_202), .A2(n_214), .B1(n_603), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_203), .A2(n_316), .B1(n_399), .B2(n_404), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_205), .B(n_506), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_207), .A2(n_264), .B1(n_838), .B2(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_208), .A2(n_324), .B1(n_499), .B2(n_605), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_209), .Y(n_866) );
XNOR2xp5_ASAP7_75t_L g871 ( .A(n_211), .B(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_212), .A2(n_241), .B1(n_562), .B2(n_845), .Y(n_844) );
AND2x2_ASAP7_75t_L g342 ( .A(n_217), .B(n_343), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_218), .A2(n_291), .B1(n_432), .B2(n_452), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_226), .A2(n_235), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_229), .A2(n_279), .B1(n_512), .B2(n_514), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_232), .A2(n_278), .B1(n_539), .B2(n_572), .Y(n_935) );
INVx1_ASAP7_75t_L g800 ( .A(n_233), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_234), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_242), .A2(n_283), .B1(n_409), .B2(n_413), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_244), .B(n_506), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_246), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_247), .A2(n_323), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_250), .A2(n_333), .B1(n_557), .B2(n_644), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_251), .Y(n_782) );
INVx1_ASAP7_75t_L g360 ( .A(n_252), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_252), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_253), .A2(n_258), .B1(n_409), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g632 ( .A(n_254), .Y(n_632) );
INVx1_ASAP7_75t_L g705 ( .A(n_255), .Y(n_705) );
INVx1_ASAP7_75t_L g579 ( .A(n_256), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_260), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_261), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_263), .A2(n_302), .B1(n_404), .B2(n_512), .Y(n_696) );
INVx1_ASAP7_75t_L g704 ( .A(n_265), .Y(n_704) );
INVx1_ASAP7_75t_L g568 ( .A(n_267), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_268), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_270), .A2(n_310), .B1(n_417), .B2(n_509), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_275), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_277), .A2(n_303), .B1(n_611), .B2(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g882 ( .A(n_280), .B(n_410), .Y(n_882) );
AO22x2_ASAP7_75t_L g893 ( .A1(n_282), .A2(n_894), .B1(n_912), .B2(n_913), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_282), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_287), .Y(n_829) );
INVx1_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_289), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g339 ( .A(n_290), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_293), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_294), .B(n_609), .Y(n_995) );
INVx1_ASAP7_75t_L g590 ( .A(n_295), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_296), .B(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g826 ( .A(n_298), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_300), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_301), .B(n_505), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_305), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_306), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_307), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_308), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_312), .Y(n_712) );
INVx1_ASAP7_75t_L g942 ( .A(n_314), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_317), .B(n_609), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_321), .Y(n_939) );
INVx1_ASAP7_75t_L g560 ( .A(n_326), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_328), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_329), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_330), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_332), .Y(n_660) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_339), .Y(n_978) );
OAI21xp5_ASAP7_75t_L g1013 ( .A1(n_340), .A2(n_977), .B(n_1014), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_723), .B1(n_972), .B2(n_973), .C(n_974), .Y(n_344) );
INVx1_ASAP7_75t_L g972 ( .A(n_345), .Y(n_972) );
AOI22xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B1(n_618), .B2(n_619), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
XNOR2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_549), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_435), .B1(n_547), .B2(n_548), .Y(n_348) );
INVx1_ASAP7_75t_L g547 ( .A(n_349), .Y(n_547) );
INVx1_ASAP7_75t_SL g434 ( .A(n_351), .Y(n_434) );
NAND4xp75_ASAP7_75t_L g351 ( .A(n_352), .B(n_388), .C(n_407), .D(n_423), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_378), .Y(n_352) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g483 ( .A(n_355), .Y(n_483) );
INVx2_ASAP7_75t_L g502 ( .A(n_355), .Y(n_502) );
OAI221xp5_ASAP7_75t_SL g563 ( .A1(n_355), .A2(n_564), .B1(n_565), .B2(n_568), .C(n_569), .Y(n_563) );
INVx3_ASAP7_75t_L g603 ( .A(n_355), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g813 ( .A1(n_355), .A2(n_513), .B1(n_814), .B2(n_815), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_355), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
INVx6_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g544 ( .A(n_356), .Y(n_544) );
BUFx3_ASAP7_75t_L g886 ( .A(n_356), .Y(n_886) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_366), .Y(n_356) );
AND2x2_ASAP7_75t_L g392 ( .A(n_357), .B(n_376), .Y(n_392) );
AND2x6_ASAP7_75t_L g395 ( .A(n_357), .B(n_396), .Y(n_395) );
AND2x6_ASAP7_75t_L g425 ( .A(n_357), .B(n_422), .Y(n_425) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_363), .Y(n_357) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_364), .Y(n_403) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_359), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_359), .B(n_364), .Y(n_387) );
AND2x2_ASAP7_75t_L g419 ( .A(n_359), .B(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_362), .Y(n_365) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g375 ( .A(n_364), .Y(n_375) );
INVx1_ASAP7_75t_L g429 ( .A(n_364), .Y(n_429) );
AND2x2_ASAP7_75t_L g382 ( .A(n_366), .B(n_374), .Y(n_382) );
AND2x6_ASAP7_75t_L g414 ( .A(n_366), .B(n_403), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_366), .B(n_403), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_366), .B(n_374), .Y(n_821) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g377 ( .A(n_367), .Y(n_377) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
OR2x2_ASAP7_75t_L g397 ( .A(n_367), .B(n_368), .Y(n_397) );
AND2x2_ASAP7_75t_L g422 ( .A(n_367), .B(n_369), .Y(n_422) );
AND2x2_ASAP7_75t_L g376 ( .A(n_368), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g745 ( .A(n_372), .Y(n_745) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g487 ( .A(n_373), .Y(n_487) );
BUFx3_ASAP7_75t_L g498 ( .A(n_373), .Y(n_498) );
BUFx3_ASAP7_75t_L g645 ( .A(n_373), .Y(n_645) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_374), .B(n_376), .Y(n_567) );
INVx1_ASAP7_75t_L g421 ( .A(n_375), .Y(n_421) );
AND2x4_ASAP7_75t_L g402 ( .A(n_376), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g405 ( .A(n_376), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g428 ( .A(n_377), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g464 ( .A(n_377), .Y(n_464) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g649 ( .A(n_380), .Y(n_649) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx5_ASAP7_75t_L g479 ( .A(n_381), .Y(n_479) );
INVx2_ASAP7_75t_L g516 ( .A(n_381), .Y(n_516) );
INVx1_ASAP7_75t_L g539 ( .A(n_381), .Y(n_539) );
BUFx3_ASAP7_75t_L g571 ( .A(n_381), .Y(n_571) );
INVx3_ASAP7_75t_L g692 ( .A(n_381), .Y(n_692) );
INVx8_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx4f_ASAP7_75t_SL g480 ( .A(n_384), .Y(n_480) );
BUFx2_ASAP7_75t_L g540 ( .A(n_384), .Y(n_540) );
BUFx2_ASAP7_75t_L g650 ( .A(n_384), .Y(n_650) );
INVx6_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g572 ( .A(n_385), .Y(n_572) );
INVx1_ASAP7_75t_SL g694 ( .A(n_385), .Y(n_694) );
OR2x6_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
INVx1_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_398), .Y(n_388) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx3_ASAP7_75t_L g474 ( .A(n_391), .Y(n_474) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_391), .Y(n_557) );
INVx3_ASAP7_75t_L g739 ( .A(n_391), .Y(n_739) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g513 ( .A(n_392), .Y(n_513) );
BUFx2_ASAP7_75t_SL g854 ( .A(n_392), .Y(n_854) );
BUFx2_ASAP7_75t_SL g962 ( .A(n_392), .Y(n_962) );
INVx1_ASAP7_75t_L g559 ( .A(n_393), .Y(n_559) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g501 ( .A(n_394), .Y(n_501) );
OAI221xp5_ASAP7_75t_SL g731 ( .A1(n_394), .A2(n_732), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_731) );
INVx4_ASAP7_75t_L g775 ( .A(n_394), .Y(n_775) );
INVx11_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx11_ASAP7_75t_L g599 ( .A(n_395), .Y(n_599) );
AND2x4_ASAP7_75t_L g412 ( .A(n_396), .B(n_403), .Y(n_412) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g445 ( .A(n_397), .B(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g476 ( .A(n_402), .Y(n_476) );
BUFx3_ASAP7_75t_L g514 ( .A(n_402), .Y(n_514) );
BUFx3_ASAP7_75t_L g537 ( .A(n_402), .Y(n_537) );
BUFx3_ASAP7_75t_L g605 ( .A(n_402), .Y(n_605) );
INVx1_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g488 ( .A(n_405), .Y(n_488) );
BUFx3_ASAP7_75t_L g499 ( .A(n_405), .Y(n_499) );
BUFx3_ASAP7_75t_L g562 ( .A(n_405), .Y(n_562) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_405), .Y(n_646) );
BUFx3_ASAP7_75t_L g734 ( .A(n_405), .Y(n_734) );
INVx1_ASAP7_75t_L g819 ( .A(n_405), .Y(n_819) );
BUFx2_ASAP7_75t_SL g960 ( .A(n_405), .Y(n_960) );
AND2x2_ASAP7_75t_L g777 ( .A(n_406), .B(n_464), .Y(n_777) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_408), .B(n_415), .Y(n_407) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx5_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g505 ( .A(n_411), .Y(n_505) );
INVx2_ASAP7_75t_L g533 ( .A(n_411), .Y(n_533) );
INVx2_ASAP7_75t_L g609 ( .A(n_411), .Y(n_609) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx4f_ASAP7_75t_L g506 ( .A(n_414), .Y(n_506) );
INVx1_ASAP7_75t_SL g842 ( .A(n_414), .Y(n_842) );
BUFx2_ASAP7_75t_L g994 ( .A(n_414), .Y(n_994) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g508 ( .A(n_417), .Y(n_508) );
BUFx3_ASAP7_75t_L g611 ( .A(n_417), .Y(n_611) );
INVx1_ASAP7_75t_L g955 ( .A(n_417), .Y(n_955) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x4_ASAP7_75t_L g427 ( .A(n_419), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g432 ( .A(n_419), .B(n_433), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_419), .B(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g509 ( .A(n_420), .Y(n_509) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_420), .Y(n_612) );
BUFx2_ASAP7_75t_SL g662 ( .A(n_420), .Y(n_662) );
BUFx2_ASAP7_75t_SL g689 ( .A(n_420), .Y(n_689) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVx1_ASAP7_75t_L g469 ( .A(n_422), .Y(n_469) );
INVx3_ASAP7_75t_L g901 ( .A(n_424), .Y(n_901) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_425), .Y(n_455) );
INVx4_ASAP7_75t_L g519 ( .A(n_425), .Y(n_519) );
INVx2_ASAP7_75t_L g527 ( .A(n_425), .Y(n_527) );
INVx2_ASAP7_75t_SL g807 ( .A(n_425), .Y(n_807) );
INVx2_ASAP7_75t_L g861 ( .A(n_425), .Y(n_861) );
INVx1_ASAP7_75t_L g711 ( .A(n_426), .Y(n_711) );
BUFx4f_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
BUFx2_ASAP7_75t_L g581 ( .A(n_427), .Y(n_581) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_427), .Y(n_614) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_427), .Y(n_685) );
INVx1_ASAP7_75t_L g433 ( .A(n_429), .Y(n_433) );
BUFx4f_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
BUFx12f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_432), .Y(n_458) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_432), .Y(n_585) );
INVx3_ASAP7_75t_L g548 ( .A(n_435), .Y(n_548) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_491), .B2(n_492), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_471), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_450), .C(n_460), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_447), .B2(n_448), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_443), .A2(n_750), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g576 ( .A(n_444), .Y(n_576) );
INVx2_ASAP7_75t_L g631 ( .A(n_444), .Y(n_631) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_445), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_445), .A2(n_800), .B(n_801), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_448), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
OA211x2_ASAP7_75t_L g606 ( .A1(n_448), .A2(n_607), .B(n_608), .C(n_610), .Y(n_606) );
BUFx3_ASAP7_75t_L g633 ( .A(n_448), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_448), .A2(n_576), .B1(n_704), .B2(n_705), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_448), .A2(n_463), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx2_ASAP7_75t_L g924 ( .A(n_448), .Y(n_924) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g751 ( .A(n_449), .Y(n_751) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_456), .C1(n_457), .C2(n_459), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_451), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
INVx3_ASAP7_75t_L g877 ( .A(n_451), .Y(n_877) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g789 ( .A(n_452), .Y(n_789) );
BUFx2_ASAP7_75t_L g835 ( .A(n_452), .Y(n_835) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_454), .A2(n_579), .B1(n_580), .B2(n_582), .C(n_583), .Y(n_578) );
OAI21xp33_ASAP7_75t_SL g634 ( .A1(n_454), .A2(n_635), .B(n_636), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_454), .A2(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g755 ( .A(n_455), .Y(n_755) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g758 ( .A(n_458), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_465), .B2(n_466), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_462), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx4_ASAP7_75t_L g589 ( .A(n_463), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_463), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_637) );
BUFx3_ASAP7_75t_L g762 ( .A(n_463), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_466), .A2(n_587), .B1(n_588), .B2(n_590), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_466), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g640 ( .A(n_468), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_468), .A2(n_588), .B1(n_904), .B2(n_905), .Y(n_903) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_477), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI21xp5_ASAP7_75t_SL g810 ( .A1(n_476), .A2(n_811), .B(n_812), .Y(n_810) );
INVx2_ASAP7_75t_L g845 ( .A(n_476), .Y(n_845) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AO22x2_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_523), .B2(n_546), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
XOR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_522), .Y(n_494) );
NAND4xp75_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .C(n_510), .D(n_517), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g938 ( .A(n_501), .Y(n_938) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx1_ASAP7_75t_L g881 ( .A(n_506), .Y(n_881) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g597 ( .A(n_513), .Y(n_597) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_514), .Y(n_742) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_516), .Y(n_737) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g787 ( .A1(n_519), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g931 ( .A(n_520), .Y(n_931) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx4_ASAP7_75t_SL g546 ( .A(n_523), .Y(n_546) );
XOR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_545), .Y(n_523) );
NAND3x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .C(n_541), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
OAI21xp5_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_527), .A2(n_660), .B(n_661), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_527), .A2(n_687), .B(n_688), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g947 ( .A1(n_527), .A2(n_948), .B(n_949), .Y(n_947) );
OAI21xp5_ASAP7_75t_SL g997 ( .A1(n_527), .A2(n_998), .B(n_999), .Y(n_997) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .C(n_534), .Y(n_530) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_593), .B1(n_616), .B2(n_617), .Y(n_549) );
INVx1_ASAP7_75t_SL g616 ( .A(n_550), .Y(n_616) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g592 ( .A(n_553), .Y(n_592) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_554), .B(n_573), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_563), .Y(n_554) );
OAI221xp5_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_558), .B1(n_559), .B2(n_560), .C(n_561), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_556), .A2(n_565), .B1(n_941), .B2(n_942), .Y(n_940) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_567), .B(n_823), .Y(n_822) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .C(n_586), .Y(n_573) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx3_ASAP7_75t_SL g781 ( .A(n_589), .Y(n_781) );
INVx2_ASAP7_75t_SL g617 ( .A(n_593), .Y(n_617) );
XOR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_615), .Y(n_593) );
NAND4xp75_ASAP7_75t_L g594 ( .A(n_595), .B(n_601), .C(n_606), .D(n_613), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g654 ( .A(n_598), .Y(n_654) );
INVx5_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_599), .B(n_825), .Y(n_824) );
INVx4_ASAP7_75t_L g889 ( .A(n_599), .Y(n_889) );
INVx2_ASAP7_75t_SL g911 ( .A(n_599), .Y(n_911) );
INVx2_ASAP7_75t_L g959 ( .A(n_599), .Y(n_959) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_SL g839 ( .A(n_612), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_614), .Y(n_753) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_675), .B2(n_722), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AO22x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_656), .B2(n_674), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_641), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .C(n_637), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_631), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_651), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
BUFx4f_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx3_ASAP7_75t_SL g674 ( .A(n_656), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_656), .A2(n_674), .B1(n_699), .B2(n_700), .Y(n_698) );
XOR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_673), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_658), .B(n_666), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_663), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx2_ASAP7_75t_L g722 ( .A(n_675), .Y(n_722) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OA22x2_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_698), .B2(n_721), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
XOR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_697), .Y(n_678) );
NAND4xp75_ASAP7_75t_SL g679 ( .A(n_680), .B(n_690), .C(n_695), .D(n_696), .Y(n_679) );
NOR2xp67_ASAP7_75t_SL g680 ( .A(n_681), .B(n_686), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .C(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g929 ( .A(n_685), .Y(n_929) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_685), .Y(n_950) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g721 ( .A(n_698), .Y(n_721) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
XNOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_720), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_713), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .C(n_709), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g973 ( .A(n_723), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_792), .B2(n_971), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_727), .B1(n_766), .B2(n_791), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g765 ( .A(n_729), .Y(n_765) );
AND2x2_ASAP7_75t_SL g729 ( .A(n_730), .B(n_746), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_738), .Y(n_730) );
INVx2_ASAP7_75t_L g891 ( .A(n_733), .Y(n_891) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI221xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_740), .B1(n_741), .B2(n_743), .C(n_744), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_752), .C(n_760), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_750), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_779) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI222xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .C1(n_757), .C2(n_759), .Y(n_752) );
OAI21xp5_ASAP7_75t_SL g832 ( .A1(n_755), .A2(n_833), .B(n_834), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_755), .A2(n_875), .B(n_876), .Y(n_874) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g791 ( .A(n_766), .Y(n_791) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NAND3x1_ASAP7_75t_SL g769 ( .A(n_770), .B(n_773), .C(n_778), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_783), .C(n_787), .Y(n_778) );
OAI21xp5_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_785), .B(n_786), .Y(n_783) );
INVx1_ASAP7_75t_L g971 ( .A(n_792), .Y(n_971) );
XOR2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_867), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_827), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
XNOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_826), .Y(n_796) );
AND3x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_809), .C(n_816), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .C(n_805), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .Y(n_809) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_822), .C(n_824), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_817) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_850), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_843), .C(n_847), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_836), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_840), .Y(n_836) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .Y(n_843) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
XOR2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_866), .Y(n_850) );
NAND4xp75_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .C(n_855), .D(n_858), .Y(n_851) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_863), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B(n_862), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_914), .B1(n_969), .B2(n_970), .Y(n_867) );
INVx1_ASAP7_75t_L g969 ( .A(n_868), .Y(n_969) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AO22x1_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B1(n_892), .B2(n_893), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND4xp75_ASAP7_75t_SL g872 ( .A(n_873), .B(n_884), .C(n_888), .D(n_890), .Y(n_872) );
NOR2xp67_ASAP7_75t_L g873 ( .A(n_874), .B(n_878), .Y(n_873) );
NAND3xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_882), .C(n_883), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
XNOR2x2_ASAP7_75t_L g943 ( .A(n_893), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_SL g912 ( .A(n_894), .Y(n_912) );
AND2x2_ASAP7_75t_SL g894 ( .A(n_895), .B(n_906), .Y(n_894) );
NOR3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .C(n_903), .Y(n_895) );
OAI21xp33_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .B(n_902), .Y(n_899) );
AND4x1_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .C(n_909), .D(n_910), .Y(n_906) );
INVx2_ASAP7_75t_SL g970 ( .A(n_914), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B1(n_943), .B2(n_968), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
XNOR2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_932), .Y(n_919) );
OAI211xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B(n_925), .C(n_926), .Y(n_921) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_927) );
NOR3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .C(n_940), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx2_ASAP7_75t_L g968 ( .A(n_943), .Y(n_968) );
INVx2_ASAP7_75t_SL g966 ( .A(n_945), .Y(n_966) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_956), .Y(n_945) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_951), .Y(n_946) );
NAND2xp5_ASAP7_75t_SL g951 ( .A(n_952), .B(n_953), .Y(n_951) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_963), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_961), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
NOR2x1_ASAP7_75t_L g975 ( .A(n_976), .B(n_980), .Y(n_975) );
OR2x2_ASAP7_75t_SL g1021 ( .A(n_976), .B(n_981), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_979), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_978), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_978), .B(n_1011), .Y(n_1014) );
CKINVDCx16_ASAP7_75t_R g1011 ( .A(n_979), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
OAI322xp33_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_1008), .A3(n_1009), .B1(n_1012), .B2(n_1015), .C1(n_1016), .C2(n_1019), .Y(n_987) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
XOR2x2_ASAP7_75t_SL g1018 ( .A(n_990), .B(n_1015), .Y(n_1018) );
NAND2x1p5_ASAP7_75t_L g990 ( .A(n_991), .B(n_1000), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_997), .Y(n_991) );
NAND3xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_995), .C(n_996), .Y(n_992) );
NOR2x1_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
CKINVDCx16_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_SL g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_1020), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_1021), .Y(n_1020) );
endmodule