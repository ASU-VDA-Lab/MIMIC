module fake_jpeg_21610_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_15),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_13),
.A2(n_17),
.B1(n_9),
.B2(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_18),
.B1(n_10),
.B2(n_0),
.Y(n_19)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

XNOR2x1_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_9),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.C(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_20),
.B1(n_13),
.B2(n_12),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_8),
.B1(n_6),
.B2(n_11),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_17),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_16),
.C(n_15),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

AOI221xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.C(n_25),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_27),
.C(n_20),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_35),
.C(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

AO221x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_5),
.B2(n_11),
.C(n_21),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_29),
.C(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_5),
.Y(n_39)
);


endmodule