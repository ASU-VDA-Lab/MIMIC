module fake_jpeg_31372_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_27),
.B(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_18),
.B1(n_43),
.B2(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_57),
.B1(n_56),
.B2(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_0),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_0),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_59),
.B1(n_49),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_58),
.B1(n_48),
.B2(n_51),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_55),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_5),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_22),
.B1(n_39),
.B2(n_38),
.Y(n_92)
);

FAx1_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_50),
.CI(n_56),
.CON(n_81),
.SN(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_87),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_88),
.B1(n_92),
.B2(n_44),
.Y(n_106)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_10),
.Y(n_101)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_11),
.Y(n_103)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_80),
.B1(n_7),
.B2(n_6),
.Y(n_98)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_106),
.B1(n_28),
.B2(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_103),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_12),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_15),
.B(n_16),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_35),
.B(n_26),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_20),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_119),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_34),
.B1(n_108),
.B2(n_112),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_100),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_107),
.B(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_122),
.A3(n_123),
.B1(n_121),
.B2(n_125),
.C(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_125),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_131),
.B(n_133),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_121),
.C(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);


endmodule