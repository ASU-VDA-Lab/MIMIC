module fake_jpeg_28358_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_32),
.B1(n_24),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_59),
.B1(n_20),
.B2(n_23),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_17),
.B1(n_29),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_40),
.B1(n_17),
.B2(n_20),
.Y(n_77)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_41),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_79),
.B1(n_85),
.B2(n_88),
.Y(n_91)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_87),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_38),
.B1(n_37),
.B2(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_38),
.B1(n_37),
.B2(n_43),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_69),
.B1(n_86),
.B2(n_54),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_54),
.B(n_2),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_31),
.B(n_78),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_34),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_1),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_49),
.B1(n_55),
.B2(n_45),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_103),
.B1(n_106),
.B2(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_47),
.B1(n_30),
.B2(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_58),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_47),
.B1(n_23),
.B2(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_68),
.B1(n_76),
.B2(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_47),
.B1(n_33),
.B2(n_25),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_73),
.B1(n_66),
.B2(n_81),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_74),
.C(n_68),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_124),
.C(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_84),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_25),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_99),
.B(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_107),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_136),
.B1(n_105),
.B2(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_18),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_25),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_28),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_1),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_105),
.B(n_109),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_149),
.B(n_155),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_109),
.B(n_90),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_90),
.B1(n_93),
.B2(n_97),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_130),
.B(n_115),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_124),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_176),
.C(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_126),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_164),
.B1(n_148),
.B2(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_147),
.B1(n_157),
.B2(n_142),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_120),
.C(n_123),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_140),
.C(n_131),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_168),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_136),
.B(n_139),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_159),
.B(n_146),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_158),
.C(n_163),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_146),
.C(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_118),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_138),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_194),
.C(n_186),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_172),
.B(n_183),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_192),
.B1(n_167),
.B2(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_147),
.B1(n_144),
.B2(n_141),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_161),
.B1(n_121),
.B2(n_149),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_149),
.C(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_203),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_156),
.B1(n_93),
.B2(n_99),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_178),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_208),
.A2(n_216),
.B1(n_200),
.B2(n_201),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_213),
.Y(n_222)
);

AOI31xp67_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_182),
.A3(n_172),
.B(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_189),
.C(n_202),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_187),
.C(n_194),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_176),
.C(n_15),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_15),
.B1(n_3),
.B2(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_202),
.C(n_191),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_200),
.B1(n_28),
.B2(n_5),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_226),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_9),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_209),
.A3(n_215),
.B1(n_216),
.B2(n_208),
.C1(n_205),
.C2(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_211),
.B(n_7),
.C(n_8),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_230),
.B(n_233),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_218),
.B(n_221),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_9),
.B(n_10),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_226),
.C(n_222),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_228),
.B1(n_14),
.B2(n_11),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_222),
.B(n_13),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_239),
.B1(n_14),
.B2(n_31),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_14),
.C(n_242),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_246),
.B(n_244),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_247),
.B(n_245),
.CI(n_241),
.CON(n_248),
.SN(n_248)
);


endmodule