module fake_jpeg_16668_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_52),
.Y(n_57)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_1),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_3),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_34),
.B1(n_40),
.B2(n_37),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_53),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_18),
.B1(n_33),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_36),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_1),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_2),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

AOI22x1_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_13),
.B1(n_28),
.B2(n_27),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_5),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_72),
.B1(n_64),
.B2(n_6),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_78),
.B1(n_76),
.B2(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_7),
.C(n_9),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_82),
.C(n_11),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_91),
.B(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_92),
.C(n_76),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_88),
.B1(n_12),
.B2(n_19),
.Y(n_95)
);

AOI31xp33_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_10),
.A3(n_20),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_24),
.Y(n_99)
);


endmodule