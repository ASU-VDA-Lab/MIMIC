module fake_jpeg_6446_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_33),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_24),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_36),
.C(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_38),
.B1(n_42),
.B2(n_32),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_25),
.B1(n_32),
.B2(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_28),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_18),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_56),
.Y(n_82)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_71),
.B1(n_27),
.B2(n_61),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_74),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_41),
.B1(n_26),
.B2(n_29),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_86),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_93),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_54),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_92),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_51),
.B(n_46),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_97),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_35),
.B(n_23),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_103),
.Y(n_124)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_27),
.B1(n_66),
.B2(n_63),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_47),
.B(n_55),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_109),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_79),
.Y(n_122)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_18),
.C(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_118),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_117),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_62),
.B1(n_80),
.B2(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_130),
.B1(n_133),
.B2(n_81),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_116),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_88),
.B(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_62),
.B1(n_67),
.B2(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_87),
.B1(n_95),
.B2(n_32),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_65),
.B1(n_73),
.B2(n_25),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_88),
.B(n_107),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_144),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_128),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_148),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_123),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_96),
.B1(n_90),
.B2(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_154),
.B1(n_155),
.B2(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_99),
.C(n_109),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_158),
.C(n_149),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_157),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_97),
.B1(n_95),
.B2(n_81),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_98),
.B(n_87),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_116),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_60),
.C(n_106),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_113),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_165),
.B(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_124),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_170),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_156),
.B(n_147),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_173),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_146),
.B1(n_135),
.B2(n_30),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_30),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_178),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_18),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_93),
.B(n_25),
.C(n_24),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_161),
.B(n_158),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_106),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_30),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_154),
.B1(n_153),
.B2(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_189),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_151),
.B1(n_141),
.B2(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_196),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_30),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_167),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_20),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_163),
.C(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_214),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_215),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_180),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_166),
.C(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_164),
.C(n_176),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_169),
.C(n_174),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_185),
.B(n_172),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_187),
.B1(n_198),
.B2(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_222),
.B1(n_227),
.B2(n_206),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_224),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_225),
.C(n_12),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_193),
.B1(n_197),
.B2(n_200),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_198),
.B(n_192),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_219),
.B(n_226),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_195),
.Y(n_224)
);

OAI322xp33_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_202),
.A3(n_179),
.B1(n_181),
.B2(n_22),
.C1(n_15),
.C2(n_5),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_235),
.B1(n_230),
.B2(n_234),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_206),
.B1(n_209),
.B2(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_212),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_0),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_227),
.C(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_0),
.B1(n_4),
.B2(n_7),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

AOI21x1_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_4),
.B(n_7),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_9),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_242),
.B(n_238),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_248),
.B(n_9),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_7),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_249),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_251),
.B(n_9),
.C(n_10),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_245),
.B(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_10),
.C(n_11),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_252),
.B(n_11),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_12),
.Y(n_256)
);


endmodule