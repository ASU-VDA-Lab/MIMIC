module fake_jpeg_10719_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_21),
.B1(n_36),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_48),
.B1(n_46),
.B2(n_42),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_58),
.Y(n_59)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_47),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_45),
.B1(n_24),
.B2(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_3),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_79),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_45),
.C(n_23),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_81),
.C(n_6),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_78),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_65),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_86),
.B1(n_27),
.B2(n_29),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_45),
.C(n_20),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_5),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_15),
.B1(n_33),
.B2(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_13),
.B(n_30),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_93),
.C(n_98),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_11),
.B(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_74),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_91),
.C(n_88),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_102),
.B(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_87),
.B(n_100),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_108),
.A3(n_105),
.B1(n_98),
.B2(n_89),
.C1(n_101),
.C2(n_37),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_7),
.Y(n_114)
);


endmodule