module fake_jpeg_18144_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_66),
.B1(n_67),
.B2(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_61),
.B1(n_37),
.B2(n_45),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_17),
.B(n_26),
.C(n_25),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_21),
.B(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_36),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_36),
.B(n_23),
.Y(n_109)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_73),
.B(n_84),
.Y(n_123)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_88),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_40),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_104),
.B(n_107),
.Y(n_124)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_56),
.B1(n_72),
.B2(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_57),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_46),
.B1(n_38),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_86),
.B1(n_108),
.B2(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_25),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_137)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_93),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_44),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_42),
.C(n_57),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_46),
.B1(n_38),
.B2(n_45),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_101),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_109),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_21),
.B1(n_17),
.B2(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_65),
.B1(n_68),
.B2(n_54),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_71),
.B1(n_77),
.B2(n_89),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_65),
.B1(n_68),
.B2(n_56),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_118),
.B1(n_137),
.B2(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_68),
.B1(n_56),
.B2(n_43),
.Y(n_118)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_76),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_139),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_94),
.C(n_107),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_12),
.B(n_16),
.Y(n_138)
);

AOI22x1_ASAP7_75t_R g171 ( 
.A1(n_138),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_42),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_145),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_109),
.B(n_96),
.C(n_75),
.D(n_85),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_156),
.B(n_170),
.Y(n_186)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_149),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_78),
.A3(n_105),
.B1(n_75),
.B2(n_80),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_164),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_100),
.B1(n_98),
.B2(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_113),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_167),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_172),
.B1(n_115),
.B2(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_36),
.B(n_30),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_88),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_79),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_19),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_30),
.B(n_19),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_49),
.B(n_90),
.C(n_19),
.D(n_30),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_133),
.Y(n_201)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_119),
.C(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_185),
.C(n_195),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_118),
.A3(n_116),
.B1(n_137),
.B2(n_112),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_196),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_131),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_148),
.B(n_164),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_142),
.B1(n_154),
.B2(n_165),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_117),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_188),
.B(n_170),
.C(n_162),
.D(n_145),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_113),
.C(n_136),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_130),
.Y(n_188)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_136),
.Y(n_196)
);

AO21x2_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_90),
.B(n_49),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_76),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_146),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_169),
.B1(n_172),
.B2(n_157),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_220),
.B(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_143),
.C(n_151),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_143),
.B(n_133),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_147),
.C(n_168),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_106),
.C(n_125),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_125),
.B1(n_11),
.B2(n_12),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_222),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_188),
.B(n_203),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_24),
.B1(n_27),
.B2(n_9),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_121),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_27),
.C(n_24),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_7),
.B(n_15),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_229),
.B1(n_184),
.B2(n_199),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_28),
.C(n_10),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_6),
.C(n_5),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_243),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_248),
.B1(n_252),
.B2(n_202),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_209),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_204),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_197),
.B1(n_190),
.B2(n_178),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_205),
.B1(n_197),
.B2(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_215),
.C(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_228),
.B1(n_190),
.B2(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_259),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_234),
.B1(n_239),
.B2(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_211),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_211),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_264),
.C(n_269),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_224),
.C(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_268),
.A2(n_241),
.B(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_192),
.B1(n_206),
.B2(n_191),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_220),
.B1(n_189),
.B2(n_217),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_245),
.B(n_231),
.C(n_230),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_240),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_236),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_237),
.C(n_184),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_275),
.B(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_278),
.C(n_264),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_255),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_251),
.B(n_182),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_258),
.B1(n_260),
.B2(n_270),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_292),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_263),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_279),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_259),
.C(n_258),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_274),
.B1(n_284),
.B2(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_204),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_272),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_283),
.B(n_187),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_290),
.A2(n_283),
.B(n_187),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_302),
.B(n_295),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_266),
.B1(n_200),
.B2(n_245),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_292),
.C(n_294),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_298),
.Y(n_309)
);

OAI221xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_200),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_310)
);

A2O1A1O1Ixp25_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_299),
.B(n_304),
.C(n_302),
.D(n_3),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_0),
.CI(n_1),
.CON(n_314),
.SN(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_2),
.B(n_3),
.Y(n_315)
);

OAI21x1_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_312),
.B(n_315),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_3),
.B1(n_4),
.B2(n_312),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);


endmodule