module fake_jpeg_9036_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_30),
.Y(n_44)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_16),
.B(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_43),
.B1(n_25),
.B2(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_21),
.Y(n_54)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_31),
.B1(n_30),
.B2(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_42),
.C(n_48),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_4),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_32),
.C(n_26),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_38),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_50),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_35),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_68),
.B(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_70),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_11),
.C(n_4),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_7),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_52),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_81),
.C(n_84),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_84),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_52),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_32),
.C(n_41),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_68),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_76),
.C(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_92),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_51),
.B1(n_36),
.B2(n_47),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_90),
.B(n_80),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_74),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_81),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_32),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_85),
.C(n_91),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_89),
.B1(n_86),
.B2(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_47),
.B1(n_41),
.B2(n_29),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_100),
.B(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_99),
.C(n_41),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_12),
.B(n_2),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_9),
.CI(n_15),
.CON(n_107),
.SN(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.B1(n_2),
.B2(n_19),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_19),
.Y(n_110)
);


endmodule