module fake_jpeg_28690_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_1),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_29),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_0),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_77),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_1),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_2),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_91),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_60),
.B1(n_68),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_56),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_68),
.B1(n_60),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_88),
.B1(n_92),
.B2(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_62),
.B1(n_63),
.B2(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_62),
.B1(n_57),
.B2(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_109),
.Y(n_112)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_106),
.Y(n_111)
);

OAI22x1_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_59),
.B1(n_52),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_23),
.B(n_49),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_13),
.B(n_14),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_10),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_127),
.B1(n_108),
.B2(n_14),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_8),
.B(n_9),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_129),
.Y(n_137)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2x1_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_11),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_131),
.B(n_112),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_12),
.B(n_13),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_38),
.B(n_41),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_33),
.B1(n_48),
.B2(n_45),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_30),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_12),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_108),
.B(n_110),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_140),
.B(n_143),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_27),
.C1(n_32),
.C2(n_35),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_138),
.B(n_139),
.C(n_144),
.D(n_145),
.Y(n_148)
);

XOR2x1_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_36),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_50),
.C(n_39),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_118),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_131),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_137),
.C(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_122),
.B(n_113),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_134),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_154),
.B(n_156),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_152),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_150),
.A3(n_151),
.B1(n_139),
.B2(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_137),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_157),
.B(n_122),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_142),
.C(n_128),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_123),
.Y(n_163)
);


endmodule