module fake_jpeg_21510_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_37),
.B1(n_36),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_47),
.B1(n_36),
.B2(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_65),
.B1(n_53),
.B2(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_76),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_78),
.B1(n_96),
.B2(n_103),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_46),
.B1(n_17),
.B2(n_25),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_79),
.A2(n_90),
.B1(n_100),
.B2(n_59),
.Y(n_139)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_45),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_21),
.B1(n_31),
.B2(n_35),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_42),
.C(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_101),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_37),
.B1(n_36),
.B2(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_31),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_40),
.C(n_44),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_45),
.C(n_44),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_40),
.B1(n_27),
.B2(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_77),
.B1(n_78),
.B2(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_22),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_34),
.CI(n_27),
.CON(n_119),
.SN(n_119)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_18),
.B(n_22),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_128),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_59),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_119),
.B(n_29),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_126),
.B1(n_129),
.B2(n_141),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_41),
.B1(n_45),
.B2(n_44),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_38),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.C(n_41),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_45),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_94),
.B1(n_85),
.B2(n_84),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_96),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_34),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_27),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_144),
.B(n_151),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_81),
.B1(n_76),
.B2(n_98),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_148),
.A2(n_162),
.B1(n_171),
.B2(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_93),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_118),
.B1(n_158),
.B2(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_159),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_95),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_28),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_116),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_109),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_94),
.B1(n_84),
.B2(n_85),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_172),
.B1(n_169),
.B2(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_71),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_71),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_19),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_74),
.B1(n_73),
.B2(n_67),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_41),
.B1(n_74),
.B2(n_86),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_20),
.B1(n_30),
.B2(n_19),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_73),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_132),
.B(n_134),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_193),
.B(n_199),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_204),
.B1(n_172),
.B2(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_198),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_203),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_118),
.B(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_147),
.C(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_33),
.C(n_16),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_154),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_116),
.B(n_141),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_129),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_9),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_124),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_168),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_130),
.C(n_113),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_125),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_216),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_211),
.A2(n_212),
.B1(n_218),
.B2(n_235),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_130),
.B1(n_127),
.B2(n_113),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_221),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_148),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_162),
.B1(n_171),
.B2(n_130),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_223),
.B1(n_225),
.B2(n_229),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_199),
.B1(n_178),
.B2(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_124),
.B1(n_127),
.B2(n_137),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_197),
.B1(n_194),
.B2(n_175),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_230),
.C(n_181),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_137),
.B1(n_156),
.B2(n_150),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_156),
.B1(n_30),
.B2(n_24),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_33),
.B(n_16),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_33),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_33),
.B1(n_16),
.B2(n_2),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_15),
.C(n_8),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_9),
.B(n_14),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_181),
.B1(n_188),
.B2(n_187),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_190),
.A2(n_0),
.B(n_1),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_176),
.B(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_176),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_239),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_175),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_255),
.B1(n_258),
.B2(n_238),
.Y(n_272)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_183),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.C(n_219),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_256),
.C(n_218),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_231),
.B1(n_230),
.B2(n_226),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_211),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_179),
.B1(n_192),
.B2(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_207),
.C(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_185),
.B1(n_188),
.B2(n_187),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_264),
.C(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_272),
.B1(n_273),
.B2(n_277),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_210),
.C(n_225),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_210),
.C(n_220),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_232),
.B1(n_233),
.B2(n_213),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_276),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_213),
.B1(n_185),
.B2(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_228),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_264),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_246),
.B1(n_251),
.B2(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_15),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_236),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_289),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_268),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_256),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_240),
.B1(n_241),
.B2(n_250),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_265),
.B1(n_261),
.B2(n_10),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_248),
.CI(n_245),
.CON(n_289),
.SN(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_292),
.B1(n_265),
.B2(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_186),
.C(n_7),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_277),
.C(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_304),
.B1(n_0),
.B2(n_2),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_261),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.C(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_15),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_281),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_0),
.C(n_1),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_280),
.C(n_289),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_278),
.B(n_293),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_288),
.B(n_283),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_311),
.B(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_313),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_281),
.B(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_2),
.C(n_4),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_320),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_294),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_321),
.B(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_322),
.Y(n_326)
);

OAI21x1_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_318),
.B(n_308),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_326),
.B(n_295),
.C(n_294),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_295),
.C(n_303),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_319),
.B(n_301),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_4),
.B(n_5),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_5),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_6),
.B(n_326),
.Y(n_332)
);


endmodule