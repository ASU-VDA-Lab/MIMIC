module fake_jpeg_4224_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_24),
.B1(n_16),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_59),
.B1(n_31),
.B2(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_24),
.B1(n_38),
.B2(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_56),
.B1(n_57),
.B2(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_24),
.B1(n_19),
.B2(n_30),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_18),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_29),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_17),
.B1(n_19),
.B2(n_25),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_83),
.B1(n_55),
.B2(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_85),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_22),
.B(n_27),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_21),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_56),
.B1(n_17),
.B2(n_47),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_26),
.B1(n_20),
.B2(n_23),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_45),
.B1(n_54),
.B2(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_22),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_50),
.C(n_52),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_55),
.C(n_44),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_91),
.B1(n_93),
.B2(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_51),
.B1(n_62),
.B2(n_41),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_63),
.B(n_13),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_58),
.CON(n_123),
.SN(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_62),
.B1(n_21),
.B2(n_23),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_84),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_66),
.C(n_65),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_55),
.B1(n_20),
.B2(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_82),
.B(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_117),
.B1(n_27),
.B2(n_1),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_128),
.C(n_130),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_27),
.B(n_60),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_121),
.B1(n_122),
.B2(n_93),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_79),
.B1(n_81),
.B2(n_41),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_80),
.B(n_44),
.C(n_58),
.D(n_60),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_0),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_92),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_87),
.B1(n_77),
.B2(n_20),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_89),
.B1(n_109),
.B2(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_87),
.B1(n_65),
.B2(n_66),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_100),
.B1(n_102),
.B2(n_90),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_71),
.C(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_78),
.B1(n_71),
.B2(n_75),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_63),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_144),
.B1(n_122),
.B2(n_132),
.Y(n_176)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_145),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_153),
.B1(n_115),
.B2(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_91),
.B1(n_99),
.B2(n_109),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_29),
.B(n_60),
.C(n_58),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_148),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_130),
.Y(n_148)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_119),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_110),
.C(n_95),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_135),
.C(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_145),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_177),
.C(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_112),
.B1(n_127),
.B2(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_176),
.B1(n_153),
.B2(n_154),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_167),
.C(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_116),
.C(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_179),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_119),
.C(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_150),
.B(n_140),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_0),
.C(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_196),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_191),
.B1(n_198),
.B2(n_175),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_147),
.B(n_155),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_200),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_193),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_146),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_136),
.B(n_149),
.Y(n_219)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_144),
.B1(n_155),
.B2(n_159),
.Y(n_198)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_172),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_182),
.B1(n_138),
.B2(n_136),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_142),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_166),
.C(n_167),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_212),
.C(n_197),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_165),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_165),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_161),
.B1(n_164),
.B2(n_174),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_178),
.C(n_168),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_190),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_216),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_184),
.B1(n_198),
.B2(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_201),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_187),
.B1(n_183),
.B2(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_204),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_203),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_212),
.C(n_208),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_158),
.B(n_13),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_206),
.B1(n_219),
.B2(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_231),
.B1(n_2),
.B2(n_4),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_195),
.B1(n_196),
.B2(n_202),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_210),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_238),
.B(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_239),
.C(n_244),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_214),
.CI(n_158),
.CON(n_237),
.SN(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_13),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_12),
.C(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_221),
.B1(n_233),
.B2(n_226),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_225),
.B(n_227),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_251),
.B(n_9),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_244),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_250),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_224),
.B(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_259),
.B(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_236),
.A3(n_226),
.B1(n_243),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_252),
.B(n_254),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_2),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_9),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_10),
.B(n_5),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_265),
.B(n_266),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_4),
.B(n_5),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_256),
.B(n_6),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_5),
.C(n_6),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_269),
.C1(n_204),
.C2(n_235),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_270),
.C(n_7),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_7),
.B(n_8),
.Y(n_274)
);


endmodule