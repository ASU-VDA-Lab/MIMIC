module fake_jpeg_13310_n_453 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_57),
.B(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_68),
.Y(n_127)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_95),
.Y(n_132)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g151 ( 
.A(n_70),
.Y(n_151)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_73),
.Y(n_130)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_75),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_76),
.B(n_78),
.Y(n_148)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_77),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_14),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_25),
.B(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_83),
.B(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_10),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_18),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_37),
.B1(n_44),
.B2(n_48),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_41),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_94),
.B(n_116),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_32),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_36),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_110),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_55),
.B(n_4),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_4),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_5),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_27),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_115),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_27),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_94),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_56),
.B1(n_22),
.B2(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_56),
.B1(n_52),
.B2(n_51),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_22),
.B1(n_43),
.B2(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_128),
.A2(n_136),
.B1(n_141),
.B2(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_133),
.A2(n_151),
.B1(n_145),
.B2(n_129),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_50),
.B1(n_46),
.B2(n_49),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_79),
.A2(n_49),
.B1(n_46),
.B2(n_7),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_7),
.B1(n_49),
.B2(n_72),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_149),
.A2(n_182),
.B1(n_167),
.B2(n_142),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_69),
.A2(n_7),
.B1(n_91),
.B2(n_77),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_7),
.B1(n_100),
.B2(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_171),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_71),
.B(n_87),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_144),
.B(n_147),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_70),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_188),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_92),
.A2(n_65),
.B1(n_89),
.B2(n_82),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_75),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_121),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_81),
.A2(n_62),
.B1(n_104),
.B2(n_73),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_63),
.A2(n_97),
.B1(n_101),
.B2(n_96),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_105),
.A2(n_113),
.B1(n_116),
.B2(n_86),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_88),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_74),
.A2(n_29),
.B1(n_31),
.B2(n_92),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_95),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_190),
.B(n_213),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_192),
.Y(n_290)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_127),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_194),
.B(n_195),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_148),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_226),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_197),
.B(n_198),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_199),
.B(n_214),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_200),
.B(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_221),
.Y(n_252)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_146),
.A2(n_135),
.B(n_161),
.C(n_160),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_248),
.B(n_201),
.C(n_196),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_168),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_205),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_208),
.A2(n_210),
.B1(n_214),
.B2(n_212),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_137),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_149),
.B1(n_175),
.B2(n_128),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_211),
.B(n_219),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_215),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_129),
.A2(n_145),
.B1(n_166),
.B2(n_141),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_216),
.Y(n_257)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_139),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_149),
.B(n_126),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_126),
.B(n_118),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_225),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_134),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_130),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_140),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_234),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_180),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_162),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_140),
.B(n_154),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_181),
.A2(n_176),
.B1(n_179),
.B2(n_186),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_251),
.B1(n_208),
.B2(n_221),
.Y(n_265)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_154),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_239),
.Y(n_271)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_R g286 ( 
.A(n_240),
.B(n_242),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_142),
.C(n_167),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_236),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_119),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_250),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_158),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_247),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

OR2x2_ASAP7_75t_SL g248 ( 
.A(n_163),
.B(n_68),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_233),
.Y(n_292)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_119),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_133),
.A2(n_68),
.B1(n_77),
.B2(n_75),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_261),
.B(n_296),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_265),
.A2(n_273),
.B1(n_279),
.B2(n_282),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_254),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_203),
.A2(n_199),
.B(n_244),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_222),
.B(n_233),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_250),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_204),
.B(n_203),
.C(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_291),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_226),
.B1(n_240),
.B2(n_190),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_240),
.A2(n_223),
.B1(n_241),
.B2(n_234),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_225),
.A2(n_229),
.B1(n_245),
.B2(n_191),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_239),
.B(n_237),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_202),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_292),
.A2(n_260),
.B(n_259),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_192),
.B(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_308),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_301),
.A2(n_298),
.B(n_285),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_222),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_309),
.C(n_317),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_252),
.A2(n_275),
.B1(n_279),
.B2(n_255),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_305),
.B1(n_267),
.B2(n_264),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_238),
.B1(n_232),
.B2(n_207),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_257),
.A2(n_218),
.B1(n_215),
.B2(n_193),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_285),
.B(n_267),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_205),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_269),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_314),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_276),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_327),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_220),
.B1(n_217),
.B2(n_224),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_316),
.B1(n_322),
.B2(n_285),
.Y(n_347)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_228),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_227),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_319),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_235),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_276),
.B(n_206),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_321),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_282),
.B1(n_265),
.B2(n_294),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_277),
.A2(n_256),
.B(n_286),
.C(n_278),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_325),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_284),
.C(n_281),
.Y(n_351)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_330),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_270),
.B(n_261),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_291),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_332),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_268),
.B(n_288),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_254),
.B(n_268),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_253),
.Y(n_339)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_253),
.A3(n_286),
.B1(n_271),
.B2(n_287),
.C1(n_285),
.C2(n_283),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_334),
.B(n_333),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_340),
.A2(n_350),
.B(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_305),
.B1(n_300),
.B2(n_328),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_264),
.B(n_297),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_352),
.C(n_360),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_298),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_293),
.B1(n_281),
.B2(n_297),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_293),
.B1(n_283),
.B2(n_284),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_299),
.A2(n_274),
.B1(n_287),
.B2(n_315),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_274),
.B(n_302),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_302),
.A2(n_301),
.B(n_318),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_318),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_310),
.C(n_311),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_331),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_363),
.C(n_377),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_332),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_347),
.A2(n_329),
.B1(n_322),
.B2(n_320),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_374),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_346),
.Y(n_365)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

BUFx12_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_379),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_349),
.B(n_303),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_378),
.C(n_327),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_313),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_307),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_376),
.Y(n_386)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_329),
.C(n_319),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_317),
.Y(n_378)
);

BUFx12_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_381),
.B(n_342),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_382),
.B(n_344),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_359),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_393),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_335),
.Y(n_387)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_357),
.B1(n_350),
.B2(n_344),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_388),
.A2(n_399),
.B1(n_361),
.B2(n_364),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_380),
.A2(n_344),
.B(n_358),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_391),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_396),
.B(n_398),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_337),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_369),
.A2(n_359),
.B1(n_348),
.B2(n_328),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_371),
.B(n_366),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_400),
.A2(n_412),
.B(n_386),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_370),
.C(n_379),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_394),
.C(n_379),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_390),
.B1(n_385),
.B2(n_397),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_383),
.A2(n_371),
.B(n_366),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_399),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_384),
.B(n_367),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_411),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_377),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_362),
.Y(n_415)
);

BUFx12_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_388),
.A2(n_382),
.B(n_345),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_419),
.C(n_408),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_417),
.Y(n_429)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_420),
.A2(n_424),
.B(n_406),
.Y(n_426)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_391),
.C(n_393),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_422),
.B(n_410),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_408),
.B(n_363),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_415),
.B(n_338),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_426),
.A2(n_430),
.B(n_432),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_420),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_419),
.B(n_401),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_367),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_404),
.B1(n_413),
.B2(n_414),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_433),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_434),
.B(n_439),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_416),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_429),
.A2(n_422),
.B1(n_413),
.B2(n_431),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_418),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_426),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_437),
.Y(n_441)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_441),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_442),
.B(n_444),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_427),
.B(n_400),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_443),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_448),
.A2(n_434),
.B1(n_389),
.B2(n_395),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_446),
.A2(n_436),
.B1(n_447),
.B2(n_405),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_450),
.B(n_386),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_449),
.C(n_387),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_375),
.Y(n_453)
);


endmodule