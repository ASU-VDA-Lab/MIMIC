module fake_jpeg_21156_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_48),
.Y(n_55)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_66),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_43),
.C(n_44),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_99),
.C(n_40),
.Y(n_109)
);

AND2x4_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_44),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_39),
.Y(n_124)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_33),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_88),
.Y(n_126)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_84),
.B1(n_98),
.B2(n_100),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_85),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_87),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_92),
.Y(n_127)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_45),
.B1(n_41),
.B2(n_38),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_43),
.C(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_49),
.B1(n_47),
.B2(n_31),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_49),
.B1(n_45),
.B2(n_47),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_46),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_132),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_46),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_46),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_19),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_116),
.B1(n_41),
.B2(n_59),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_49),
.B1(n_47),
.B2(n_42),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_36),
.B(n_19),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_124),
.B(n_104),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_21),
.B(n_30),
.Y(n_125)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_26),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_49),
.B1(n_41),
.B2(n_38),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_134),
.B(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_142),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_122),
.B1(n_105),
.B2(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_147),
.B1(n_116),
.B2(n_132),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_26),
.B(n_19),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_74),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_154),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_160),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_149),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_74),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_20),
.B(n_23),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_39),
.Y(n_157)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_77),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_120),
.B(n_132),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_162),
.A2(n_167),
.B(n_180),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_138),
.B1(n_159),
.B2(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_115),
.B1(n_103),
.B2(n_132),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_178),
.B1(n_144),
.B2(n_10),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_117),
.B(n_106),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_121),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_182),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_128),
.B1(n_118),
.B2(n_84),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_112),
.B1(n_40),
.B2(n_17),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_128),
.B1(n_118),
.B2(n_72),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_175),
.B1(n_153),
.B2(n_145),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_183),
.B(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_41),
.B1(n_28),
.B2(n_38),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_140),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_159),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_42),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_186),
.B(n_40),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_123),
.C(n_39),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_40),
.Y(n_210)
);

OAI211xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_151),
.B(n_156),
.C(n_154),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_197),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_207),
.B1(n_172),
.B2(n_174),
.Y(n_228)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_202),
.B1(n_199),
.B2(n_184),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_147),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_191),
.B(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_138),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_29),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_6),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_204),
.B(n_217),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_32),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_32),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_15),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_32),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_112),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_85),
.CI(n_80),
.CON(n_249),
.SN(n_249)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_32),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_193),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_77),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_18),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_89),
.B1(n_27),
.B2(n_24),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_164),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_227),
.A2(n_229),
.B(n_242),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_243),
.B1(n_199),
.B2(n_206),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_162),
.B1(n_167),
.B2(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_239),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_168),
.B1(n_169),
.B2(n_29),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_248),
.B(n_197),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_168),
.C(n_53),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_210),
.C(n_203),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_223),
.B1(n_222),
.B2(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_29),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_27),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_255),
.B1(n_266),
.B2(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_258),
.C(n_261),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_208),
.B1(n_213),
.B2(n_214),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_194),
.C(n_205),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_257),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_226),
.A2(n_221),
.B1(n_215),
.B2(n_194),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_201),
.C(n_203),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_248),
.B1(n_252),
.B2(n_267),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.C(n_232),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_27),
.B1(n_24),
.B2(n_17),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_235),
.B1(n_238),
.B2(n_234),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_27),
.B1(n_24),
.B2(n_17),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_279),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_248),
.B1(n_245),
.B2(n_233),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_280),
.B1(n_289),
.B2(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_240),
.B(n_243),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_244),
.C(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_291),
.C(n_258),
.Y(n_300)
);

XNOR2x2_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_249),
.Y(n_288)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_253),
.A2(n_238),
.B1(n_251),
.B2(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_251),
.C(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_296),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_286),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_299),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_289),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_271),
.B(n_17),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_290),
.B1(n_282),
.B2(n_280),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_18),
.C(n_8),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.C(n_279),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_18),
.C(n_8),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_276),
.B1(n_1),
.B2(n_2),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_274),
.B(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_310),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_284),
.B(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_9),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_301),
.B1(n_307),
.B2(n_306),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_292),
.Y(n_320)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_323),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_306),
.C(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_326),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_9),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_328),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_11),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_324),
.A2(n_315),
.B(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_322),
.B(n_316),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_314),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_308),
.C(n_319),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_337),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_330),
.A3(n_329),
.B1(n_338),
.B2(n_335),
.C1(n_333),
.C2(n_2),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_0),
.B(n_3),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_341),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_4),
.C(n_342),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_4),
.Y(n_345)
);


endmodule