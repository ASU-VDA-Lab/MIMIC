module fake_jpeg_11876_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_42),
.B(n_34),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_71),
.C(n_76),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_6),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_1),
.B(n_2),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_4),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_16),
.B(n_30),
.C(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.C(n_90),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_76),
.B1(n_9),
.B2(n_7),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_18),
.C(n_26),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_88),
.C(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_68),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_94),
.B(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_76),
.C(n_77),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_87),
.B1(n_76),
.B2(n_81),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_80),
.B(n_82),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_91),
.B(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_97),
.B1(n_12),
.B2(n_13),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_10),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_20),
.C(n_21),
.Y(n_104)
);

NOR2xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_23),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_24),
.Y(n_106)
);


endmodule