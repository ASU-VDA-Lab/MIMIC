module real_jpeg_25255_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_86),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_86),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_96)
);

INVx8_ASAP7_75t_SL g78 ( 
.A(n_5),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_81),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_6),
.A2(n_57),
.B(n_60),
.C(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_158),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_28),
.C(n_47),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_158),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_6),
.A2(n_31),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_149),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_64),
.B1(n_70),
.B2(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_64),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_70),
.B1(n_71),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_9),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_136),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_136),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_136),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_69),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_69),
.Y(n_238)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_16),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_16),
.A2(n_32),
.B1(n_123),
.B2(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_16),
.A2(n_32),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_20),
.B(n_114),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_113),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.C(n_66),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_25),
.A2(n_38),
.B1(n_39),
.B2(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_25),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_26),
.A2(n_31),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_33),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_27),
.B(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_35),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_31),
.A2(n_165),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_31),
.A2(n_238),
.B(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_32),
.B(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_37),
.B(n_158),
.Y(n_242)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_37),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_37),
.A2(n_212),
.B(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_50),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_42),
.A2(n_58),
.B(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_43),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_45),
.A2(n_51),
.B1(n_53),
.B2(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_45),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_45),
.A2(n_53),
.B1(n_205),
.B2(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_50),
.A2(n_128),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_50),
.B(n_158),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_50),
.A2(n_153),
.B(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_53),
.B(n_154),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_54),
.B(n_66),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_65),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_55),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_55),
.A2(n_183),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_63),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_56),
.A2(n_131),
.B(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_60),
.B(n_78),
.C(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_61),
.A2(n_77),
.B(n_159),
.C(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_82),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_75),
.B1(n_81),
.B2(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_71),
.Y(n_169)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_73),
.B(n_158),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_75),
.A2(n_83),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_80),
.A2(n_111),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_93),
.A2(n_204),
.B(n_206),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_93),
.A2(n_206),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_115),
.B(n_118),
.Y(n_291)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_119),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.C(n_134),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_120),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_127),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_149),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_288),
.B(n_292),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_191),
.B(n_275),
.C(n_287),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_178),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_142),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_160),
.C(n_170),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_143),
.A2(n_144),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_151),
.C(n_155),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B(n_159),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_160),
.A2(n_161),
.B1(n_170),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_166),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_170),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_177),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_179),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.CI(n_184),
.CON(n_179),
.SN(n_179)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_180),
.B(n_181),
.C(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_268),
.B(n_274),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_223),
.B(n_267),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_215),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_215),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_214),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_197),
.B(n_203),
.C(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_261),
.B(n_266),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_251),
.B(n_260),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_239),
.B(n_250),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_246),
.B(n_249),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_259),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_286),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);


endmodule