module fake_jpeg_818_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_63),
.Y(n_223)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_70),
.Y(n_192)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_75),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_76),
.B(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_19),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_85),
.Y(n_156)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_19),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_47),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_105),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_102),
.B(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_27),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_107),
.B(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_37),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_21),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_113),
.Y(n_217)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_44),
.B(n_17),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_17),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_23),
.B(n_0),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_124),
.B(n_31),
.C(n_20),
.Y(n_180)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_48),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_0),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_50),
.Y(n_131)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_48),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_136),
.B(n_171),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_59),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_142),
.B(n_149),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_101),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_161),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_214),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g294 ( 
.A(n_169),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_183),
.Y(n_244)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_59),
.B1(n_53),
.B2(n_50),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_63),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

INVx2_ASAP7_75t_R g194 ( 
.A(n_71),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_207),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_196),
.Y(n_288)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_51),
.B(n_58),
.C(n_52),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_52),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_205),
.B(n_206),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_118),
.B(n_58),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_125),
.B(n_39),
.C(n_54),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_114),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_62),
.Y(n_220)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

HAxp5_ASAP7_75t_SL g221 ( 
.A(n_113),
.B(n_59),
.CON(n_221),
.SN(n_221)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_221),
.Y(n_256)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_224),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_61),
.A2(n_39),
.B1(n_54),
.B2(n_31),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_99),
.B1(n_72),
.B2(n_68),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_142),
.A2(n_95),
.B1(n_40),
.B2(n_43),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_228),
.A2(n_229),
.B1(n_254),
.B2(n_257),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_147),
.B1(n_151),
.B2(n_188),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_183),
.A2(n_70),
.B1(n_69),
.B2(n_73),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_237),
.A2(n_252),
.B1(n_295),
.B2(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

CKINVDCx12_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_250),
.B(n_261),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_251),
.B(n_253),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_163),
.A2(n_151),
.B1(n_147),
.B2(n_157),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_157),
.A2(n_36),
.B1(n_33),
.B2(n_20),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_146),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_255),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_146),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_45),
.B1(n_34),
.B2(n_33),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_269),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_45),
.B1(n_53),
.B2(n_59),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_178),
.A2(n_81),
.B1(n_66),
.B2(n_78),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_65),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_138),
.Y(n_262)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_156),
.B(n_90),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_263),
.B(n_265),
.Y(n_371)
);

CKINVDCx12_ASAP7_75t_R g265 ( 
.A(n_199),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_156),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_266),
.B(n_276),
.Y(n_355)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_132),
.Y(n_267)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_279),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_188),
.B(n_90),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_143),
.B(n_87),
.Y(n_273)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_275),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_136),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_87),
.B1(n_97),
.B2(n_17),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_277),
.A2(n_292),
.B1(n_160),
.B2(n_139),
.Y(n_339)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_140),
.Y(n_278)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_217),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_168),
.Y(n_281)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_175),
.B(n_79),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_286),
.C(n_223),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_133),
.B(n_162),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_284),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_148),
.B(n_0),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_164),
.Y(n_285)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_182),
.B(n_127),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_150),
.B(n_0),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_297),
.Y(n_336)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_184),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_221),
.A2(n_117),
.B1(n_2),
.B2(n_3),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_217),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_152),
.B(n_155),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_304),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g300 ( 
.A1(n_134),
.A2(n_211),
.B1(n_186),
.B2(n_174),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_211),
.Y(n_301)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_193),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_185),
.B(n_1),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_6),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_194),
.A2(n_2),
.B(n_4),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_210),
.B(n_177),
.Y(n_362)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_197),
.Y(n_308)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_200),
.Y(n_309)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_256),
.A2(n_219),
.B1(n_181),
.B2(n_226),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_244),
.B(n_223),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_315),
.Y(n_381)
);

OR2x2_ASAP7_75t_SL g316 ( 
.A(n_244),
.B(n_166),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_316),
.B(n_321),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

FAx1_ASAP7_75t_L g322 ( 
.A(n_244),
.B(n_177),
.CI(n_216),
.CON(n_322),
.SN(n_322)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_322),
.A2(n_286),
.B(n_272),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_212),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_323),
.B(n_330),
.C(n_347),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_141),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_325),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_189),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_329),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_158),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_135),
.C(n_222),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_246),
.A2(n_192),
.B1(n_186),
.B2(n_216),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_346),
.B1(n_295),
.B2(n_230),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_249),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_343),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_339),
.A2(n_294),
.B1(n_298),
.B2(n_264),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_249),
.B(n_238),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_246),
.A2(n_192),
.B1(n_134),
.B2(n_212),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_177),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_167),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_363),
.Y(n_416)
);

BUFx6f_ASAP7_75t_SL g351 ( 
.A(n_235),
.Y(n_351)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_233),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_354),
.B(n_359),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_252),
.B(n_224),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_357),
.B(n_360),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_239),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_271),
.B(n_195),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_364),
.B(n_282),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_218),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_237),
.A2(n_144),
.B(n_170),
.C(n_169),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_236),
.Y(n_366)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_241),
.B(n_195),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_368),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_248),
.B(n_196),
.Y(n_368)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_372),
.Y(n_460)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

INVx3_ASAP7_75t_SL g377 ( 
.A(n_327),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_322),
.A2(n_300),
.B1(n_262),
.B2(n_255),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_413),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_243),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_239),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_384),
.B(n_400),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_385),
.A2(n_398),
.B(n_325),
.Y(n_440)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_389),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_391),
.A2(n_403),
.B1(n_320),
.B2(n_352),
.Y(n_452)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_286),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_406),
.Y(n_423)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_268),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_369),
.A2(n_287),
.B1(n_274),
.B2(n_285),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_420),
.B1(n_340),
.B2(n_351),
.Y(n_436)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

AO21x2_ASAP7_75t_L g403 ( 
.A1(n_331),
.A2(n_308),
.B(n_291),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_405),
.B(n_409),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_313),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_365),
.B1(n_294),
.B2(n_298),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_272),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_334),
.B(n_302),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_411),
.Y(n_433)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_414),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_280),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_323),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_355),
.Y(n_439)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_365),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_369),
.A2(n_301),
.B1(n_240),
.B2(n_278),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_422),
.B(n_386),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_343),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_434),
.C(n_407),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_398),
.A2(n_363),
.B(n_362),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_428),
.B(n_444),
.Y(n_466)
);

AND2x2_ASAP7_75t_SL g431 ( 
.A(n_416),
.B(n_325),
.Y(n_431)
);

NAND2x1_ASAP7_75t_SL g475 ( 
.A(n_431),
.B(n_373),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_317),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_381),
.A2(n_328),
.B1(n_314),
.B2(n_315),
.Y(n_435)
);

OAI22x1_ASAP7_75t_L g482 ( 
.A1(n_435),
.A2(n_430),
.B1(n_437),
.B2(n_428),
.Y(n_482)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_317),
.B1(n_315),
.B2(n_364),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_437),
.A2(n_446),
.B1(n_458),
.B2(n_375),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_439),
.B(n_376),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_440),
.A2(n_456),
.B(n_378),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_416),
.A2(n_326),
.B1(n_329),
.B2(n_348),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_445),
.B1(n_449),
.B2(n_452),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_385),
.A2(n_330),
.B(n_319),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_388),
.A2(n_316),
.B1(n_312),
.B2(n_321),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_401),
.A2(n_347),
.B1(n_358),
.B2(n_340),
.Y(n_446)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_388),
.A2(n_358),
.B1(n_345),
.B2(n_370),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_370),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_461),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_345),
.B(n_324),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_383),
.A2(n_361),
.B1(n_356),
.B2(n_310),
.Y(n_458)
);

AO22x1_ASAP7_75t_L g461 ( 
.A1(n_396),
.A2(n_281),
.B1(n_361),
.B2(n_309),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_413),
.B(n_378),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_462),
.A2(n_482),
.B(n_438),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_443),
.B(n_429),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_463),
.Y(n_524)
);

MAJx2_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_453),
.C(n_426),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_467),
.A2(n_496),
.B1(n_498),
.B2(n_491),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_395),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_470),
.B(n_473),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_419),
.Y(n_471)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_383),
.C(n_404),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_477),
.C(n_431),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_399),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_474),
.B(n_487),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_480),
.C(n_494),
.Y(n_523)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_374),
.C(n_389),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_478),
.Y(n_527)
);

INVx13_ASAP7_75t_L g479 ( 
.A(n_424),
.Y(n_479)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_479),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_447),
.Y(n_480)
);

INVx13_ASAP7_75t_L g484 ( 
.A(n_424),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_484),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_485),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_486),
.B(n_445),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_439),
.B(n_337),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_488),
.B(n_490),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_456),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_489),
.B(n_497),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_430),
.A2(n_405),
.B(n_387),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_435),
.A2(n_391),
.B1(n_414),
.B2(n_403),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_491),
.A2(n_493),
.B1(n_403),
.B2(n_426),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_402),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_499),
.Y(n_507)
);

INVx11_ASAP7_75t_L g493 ( 
.A(n_425),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_433),
.B(n_380),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_231),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_450),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_423),
.A2(n_403),
.B1(n_380),
.B2(n_379),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_372),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_431),
.A2(n_403),
.B1(n_380),
.B2(n_412),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_441),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_500),
.B(n_520),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_505),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_485),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_502),
.B(n_519),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_465),
.A2(n_431),
.B1(n_446),
.B2(n_436),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_506),
.Y(n_537)
);

AO22x1_ASAP7_75t_L g506 ( 
.A1(n_498),
.A2(n_461),
.B1(n_454),
.B2(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_458),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_509),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_510),
.A2(n_511),
.B1(n_532),
.B2(n_512),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_461),
.Y(n_512)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_512),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_515),
.B(n_476),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_441),
.Y(n_516)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_337),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_517),
.A2(n_534),
.B(n_462),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_471),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_464),
.B(n_453),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_522),
.A2(n_482),
.B(n_494),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_472),
.B(n_432),
.C(n_438),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_530),
.C(n_533),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_465),
.A2(n_481),
.B1(n_468),
.B2(n_490),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_536),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_477),
.B(n_459),
.C(n_457),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_469),
.B(n_459),
.Y(n_532)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_532),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_495),
.B(n_457),
.C(n_318),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_486),
.B(n_442),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_SL g535 ( 
.A(n_466),
.B(n_397),
.C(n_332),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_488),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_481),
.A2(n_442),
.B1(n_460),
.B2(n_425),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_516),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_539),
.B(n_536),
.Y(n_577)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_542),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_544),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_518),
.Y(n_545)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_508),
.A2(n_483),
.B1(n_496),
.B2(n_468),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_546),
.A2(n_506),
.B1(n_460),
.B2(n_393),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_522),
.A2(n_489),
.B(n_475),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_563),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_518),
.Y(n_549)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_549),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_466),
.C(n_475),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_553),
.C(n_560),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_525),
.B(n_467),
.C(n_482),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_530),
.B(n_521),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_556),
.B(n_557),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_529),
.B(n_492),
.Y(n_557)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_507),
.Y(n_559)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_559),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_501),
.B(n_469),
.C(n_478),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_513),
.Y(n_561)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_561),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_497),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_562),
.B(n_505),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_523),
.A2(n_524),
.B(n_531),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_564),
.A2(n_504),
.B1(n_506),
.B2(n_511),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_565),
.B(n_500),
.Y(n_579)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_507),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_568),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_514),
.B(n_535),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_567),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_514),
.A2(n_493),
.B1(n_484),
.B2(n_479),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_533),
.B(n_332),
.C(n_310),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_526),
.C(n_503),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_560),
.B(n_528),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_570),
.B(n_589),
.C(n_567),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_SL g607 ( 
.A(n_576),
.B(n_579),
.Y(n_607)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_577),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_583),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_526),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_503),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_592),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_543),
.B(n_527),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_586),
.A2(n_563),
.B(n_566),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_588),
.A2(n_538),
.B1(n_537),
.B2(n_540),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_550),
.B(n_390),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_590),
.A2(n_593),
.B1(n_549),
.B2(n_545),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_551),
.B(n_484),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_543),
.A2(n_479),
.B1(n_377),
.B2(n_264),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_550),
.B(n_235),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_592),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_555),
.B(n_305),
.C(n_234),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_552),
.C(n_555),
.Y(n_601)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

INVx13_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_600),
.B(n_608),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_582),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_553),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_602),
.B(n_613),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_603),
.A2(n_267),
.B1(n_288),
.B2(n_245),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_569),
.C(n_565),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_604),
.B(n_612),
.C(n_579),
.Y(n_627)
);

HAxp5_ASAP7_75t_SL g605 ( 
.A(n_572),
.B(n_538),
.CON(n_605),
.SN(n_605)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_605),
.A2(n_234),
.B(n_245),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_606),
.A2(n_611),
.B1(n_615),
.B2(n_573),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_609),
.A2(n_574),
.B1(n_588),
.B2(n_581),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_584),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_575),
.B(n_562),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_578),
.B(n_548),
.C(n_542),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_544),
.Y(n_613)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_571),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_617),
.Y(n_631)
);

AOI221xp5_ASAP7_75t_L g615 ( 
.A1(n_580),
.A2(n_558),
.B1(n_559),
.B2(n_547),
.C(n_537),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_596),
.B(n_561),
.C(n_558),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_576),
.B(n_547),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_618),
.B(n_231),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_634),
.Y(n_648)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_620),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_616),
.A2(n_573),
.B(n_574),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_621),
.A2(n_636),
.B(n_632),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_622),
.B(n_607),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_623),
.B(n_630),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_597),
.A2(n_591),
.B1(n_586),
.B2(n_594),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_625),
.B(n_627),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_608),
.A2(n_587),
.B1(n_585),
.B2(n_590),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_626),
.A2(n_598),
.B1(n_607),
.B2(n_288),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_602),
.B(n_613),
.C(n_604),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_629),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_601),
.B(n_593),
.C(n_232),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_616),
.B(n_275),
.C(n_293),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_633),
.B(n_635),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_612),
.B(n_290),
.Y(n_635)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_636),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_SL g640 ( 
.A1(n_637),
.A2(n_605),
.B(n_624),
.C(n_600),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_SL g654 ( 
.A(n_640),
.B(n_646),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_618),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_642),
.B(n_242),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_643),
.B(n_649),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_644),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_622),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_645),
.A2(n_619),
.B1(n_633),
.B2(n_247),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_628),
.B(n_632),
.C(n_627),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_630),
.A2(n_247),
.B(n_242),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_652),
.A2(n_394),
.B(n_9),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_638),
.A2(n_629),
.B1(n_635),
.B2(n_634),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_653),
.B(n_655),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_646),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_656),
.B(n_657),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_645),
.B(n_6),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_659),
.B(n_660),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_651),
.A2(n_394),
.B(n_9),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_662),
.B(n_647),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_639),
.B(n_8),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_663),
.B(n_664),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_647),
.B(n_8),
.Y(n_664)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_666),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_650),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_667),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_656),
.B(n_648),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_661),
.C(n_640),
.Y(n_677)
);

AOI322xp5_ASAP7_75t_L g672 ( 
.A1(n_658),
.A2(n_640),
.A3(n_641),
.B1(n_649),
.B2(n_648),
.C1(n_14),
.C2(n_8),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_672),
.A2(n_665),
.B(n_670),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_674),
.B(n_677),
.Y(n_678)
);

AO21x1_ASAP7_75t_L g676 ( 
.A1(n_668),
.A2(n_654),
.B(n_640),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_676),
.A2(n_10),
.B(n_11),
.Y(n_680)
);

AOI332xp33_ASAP7_75t_L g679 ( 
.A1(n_673),
.A2(n_661),
.A3(n_671),
.B1(n_666),
.B2(n_669),
.B3(n_10),
.C1(n_14),
.C2(n_12),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_680),
.B(n_676),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_678),
.B(n_675),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_681),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_682),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_SL g685 ( 
.A1(n_684),
.A2(n_14),
.B(n_16),
.C(n_681),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_14),
.B(n_16),
.Y(n_686)
);


endmodule