module fake_jpeg_27001_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_39),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_35),
.B1(n_39),
.B2(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_38),
.B1(n_34),
.B2(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_46),
.B1(n_32),
.B2(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_38),
.B1(n_46),
.B2(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_75),
.Y(n_92)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_29),
.B1(n_19),
.B2(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_76),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_80),
.B1(n_38),
.B2(n_17),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_32),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_27),
.C(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_26),
.B1(n_31),
.B2(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_28),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_88),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_95),
.B1(n_103),
.B2(n_104),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_60),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_99),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_69),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_61),
.C(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_56),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_114),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_76),
.B(n_58),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_108),
.B(n_37),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_111),
.B1(n_112),
.B2(n_1),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_59),
.B(n_64),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_100),
.B1(n_89),
.B2(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_67),
.B1(n_57),
.B2(n_66),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_104),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_18),
.C(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_14),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_118),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_66),
.B1(n_61),
.B2(n_73),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_84),
.B1(n_25),
.B2(n_27),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_30),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_13),
.B(n_10),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_101),
.B(n_97),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_84),
.B(n_94),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_97),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_113),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_1),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_27),
.C(n_13),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_3),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_139),
.C(n_141),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_3),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_155),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_107),
.A3(n_110),
.B1(n_114),
.B2(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_153),
.B(n_134),
.Y(n_162)
);

NAND2x1_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_127),
.Y(n_157)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_131),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_6),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_135),
.B1(n_144),
.B2(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_129),
.B1(n_121),
.B2(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_129),
.C(n_5),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_156),
.C(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_149),
.B1(n_145),
.B2(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_153),
.B(n_152),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_4),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_6),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_168),
.C(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_9),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_160),
.B1(n_169),
.B2(n_164),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_167),
.C1(n_177),
.C2(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_170),
.C(n_160),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_186),
.B(n_9),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_165),
.B1(n_173),
.B2(n_172),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_191),
.B1(n_182),
.B2(n_180),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_190),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_196),
.B(n_194),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_188),
.Y(n_196)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_183),
.Y(n_199)
);


endmodule