module real_aes_1265_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_503;
wire n_635;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_314;
wire n_283;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_0), .A2(n_235), .B1(n_386), .B2(n_419), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_1), .A2(n_227), .B1(n_426), .B2(n_427), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_2), .A2(n_196), .B1(n_336), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_3), .A2(n_80), .B1(n_341), .B2(n_345), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_4), .A2(n_140), .B1(n_426), .B2(n_427), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_5), .A2(n_206), .B1(n_501), .B2(n_503), .Y(n_500) );
AO22x2_ASAP7_75t_L g289 ( .A1(n_6), .A2(n_184), .B1(n_279), .B2(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g678 ( .A(n_6), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_7), .A2(n_102), .B1(n_346), .B2(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_8), .A2(n_69), .B1(n_539), .B2(n_540), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_9), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_10), .A2(n_70), .B1(n_328), .B2(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_11), .A2(n_198), .B1(n_304), .B2(n_308), .Y(n_303) );
AO22x2_ASAP7_75t_L g286 ( .A1(n_12), .A2(n_55), .B1(n_279), .B2(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_12), .B(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_13), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_14), .A2(n_173), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_15), .A2(n_138), .B1(n_304), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_16), .A2(n_207), .B1(n_423), .B2(n_424), .Y(n_422) );
AO222x2_ASAP7_75t_SL g601 ( .A1(n_17), .A2(n_36), .B1(n_150), .B2(n_397), .C1(n_398), .C2(n_401), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_18), .A2(n_183), .B1(n_700), .B2(n_701), .Y(n_699) );
AO222x2_ASAP7_75t_SL g718 ( .A1(n_19), .A2(n_155), .B1(n_236), .B2(n_370), .C1(n_623), .C2(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_20), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_21), .A2(n_115), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_22), .A2(n_250), .B1(n_368), .B2(n_528), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_23), .A2(n_158), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_24), .A2(n_143), .B1(n_410), .B2(n_413), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_25), .A2(n_255), .B1(n_264), .B2(n_670), .C(n_680), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_26), .B(n_565), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_27), .A2(n_226), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_28), .A2(n_238), .B1(n_644), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_29), .A2(n_144), .B1(n_419), .B2(n_420), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_30), .A2(n_114), .B1(n_454), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_31), .A2(n_179), .B1(n_304), .B2(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_32), .A2(n_126), .B1(n_426), .B2(n_427), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_33), .A2(n_197), .B1(n_451), .B2(n_462), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_34), .A2(n_128), .B1(n_423), .B2(n_424), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_35), .A2(n_125), .B1(n_304), .B2(n_454), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_37), .A2(n_172), .B1(n_423), .B2(n_424), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_38), .A2(n_181), .B1(n_348), .B2(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_39), .A2(n_71), .B1(n_427), .B2(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_40), .A2(n_142), .B1(n_348), .B2(n_351), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_41), .A2(n_165), .B1(n_308), .B2(n_531), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_42), .A2(n_60), .B1(n_383), .B2(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_43), .A2(n_214), .B1(n_313), .B2(n_318), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_44), .A2(n_232), .B1(n_325), .B2(n_328), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_45), .A2(n_100), .B1(n_410), .B2(n_451), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_46), .A2(n_87), .B1(n_464), .B2(n_465), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_47), .A2(n_229), .B1(n_381), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_48), .A2(n_153), .B1(n_328), .B2(n_341), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g292 ( .A1(n_49), .A2(n_252), .B1(n_293), .B2(n_297), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_50), .A2(n_221), .B1(n_336), .B2(n_382), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_51), .A2(n_160), .B1(n_424), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_52), .A2(n_119), .B1(n_464), .B2(n_465), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_53), .A2(n_141), .B1(n_397), .B2(n_398), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_54), .A2(n_244), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_56), .A2(n_86), .B1(n_329), .B2(n_543), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_57), .A2(n_239), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_58), .A2(n_98), .B1(n_413), .B2(n_462), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_59), .A2(n_253), .B1(n_325), .B2(n_722), .Y(n_721) );
AO222x2_ASAP7_75t_SL g656 ( .A1(n_61), .A2(n_175), .B1(n_194), .B2(n_397), .C1(n_398), .C2(n_401), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_62), .A2(n_149), .B1(n_385), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_63), .A2(n_139), .B1(n_575), .B2(n_630), .Y(n_694) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_64), .A2(n_392), .B1(n_393), .B2(n_428), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_64), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_65), .A2(n_108), .B1(n_336), .B2(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g279 ( .A(n_66), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_67), .A2(n_93), .B1(n_482), .B2(n_547), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_68), .A2(n_248), .B1(n_501), .B2(n_701), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_72), .A2(n_233), .B1(n_397), .B2(n_398), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_73), .A2(n_135), .B1(n_424), .B2(n_520), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_74), .A2(n_217), .B1(n_397), .B2(n_398), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_75), .A2(n_189), .B1(n_420), .B2(n_612), .Y(n_664) );
AOI22x1_ASAP7_75t_L g581 ( .A1(n_76), .A2(n_582), .B1(n_583), .B2(n_596), .Y(n_581) );
INVx1_ASAP7_75t_L g596 ( .A(n_76), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_77), .A2(n_148), .B1(n_533), .B2(n_534), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_78), .A2(n_123), .B1(n_641), .B2(n_642), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_79), .A2(n_101), .B1(n_479), .B2(n_482), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_81), .A2(n_224), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_82), .A2(n_90), .B1(n_417), .B2(n_420), .Y(n_443) );
INVx1_ASAP7_75t_SL g280 ( .A(n_83), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_83), .B(n_122), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_84), .A2(n_106), .B1(n_410), .B2(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_85), .A2(n_230), .B1(n_381), .B2(n_383), .Y(n_380) );
XOR2xp5_ASAP7_75t_L g686 ( .A(n_88), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g260 ( .A(n_89), .Y(n_260) );
XOR2x2_ASAP7_75t_L g357 ( .A(n_91), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_92), .B(n_273), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_94), .A2(n_211), .B1(n_569), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_95), .A2(n_133), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_96), .A2(n_202), .B1(n_464), .B2(n_660), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_97), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_99), .A2(n_185), .B1(n_637), .B2(n_638), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_103), .A2(n_222), .B1(n_293), .B2(n_368), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_104), .A2(n_113), .B1(n_342), .B2(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_105), .B(n_364), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_107), .A2(n_186), .B1(n_419), .B2(n_420), .Y(n_467) );
XNOR2x1_ASAP7_75t_SL g268 ( .A(n_109), .B(n_269), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_110), .A2(n_129), .B1(n_629), .B2(n_630), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_111), .A2(n_240), .B1(n_378), .B2(n_379), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_112), .A2(n_213), .B1(n_314), .B2(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_116), .A2(n_242), .B1(n_367), .B2(n_369), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_117), .A2(n_187), .B1(n_341), .B2(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g504 ( .A(n_118), .Y(n_504) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_120), .A2(n_618), .B(n_647), .Y(n_617) );
INVx1_ASAP7_75t_L g649 ( .A(n_120), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_121), .A2(n_176), .B1(n_625), .B2(n_703), .Y(n_702) );
AO22x2_ASAP7_75t_L g282 ( .A1(n_122), .A2(n_195), .B1(n_279), .B2(n_283), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_124), .A2(n_146), .B1(n_369), .B2(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g621 ( .A(n_127), .B(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_130), .A2(n_249), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_131), .A2(n_231), .B1(n_708), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_132), .A2(n_208), .B1(n_419), .B2(n_420), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_134), .A2(n_241), .B1(n_696), .B2(n_697), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_136), .A2(n_152), .B1(n_441), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_137), .A2(n_157), .B1(n_413), .B2(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g281 ( .A(n_145), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_147), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_151), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_154), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_156), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_159), .A2(n_177), .B1(n_496), .B2(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_161), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_162), .A2(n_209), .B1(n_361), .B2(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_163), .B(n_273), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_164), .B(n_365), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_166), .B(n_365), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_167), .A2(n_237), .B1(n_498), .B2(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_168), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g685 ( .A(n_169), .Y(n_685) );
AO22x2_ASAP7_75t_L g712 ( .A1(n_169), .A2(n_685), .B1(n_713), .B2(n_730), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_170), .A2(n_180), .B1(n_336), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_171), .A2(n_191), .B1(n_424), .B2(n_520), .Y(n_573) );
AO22x1_ASAP7_75t_L g624 ( .A1(n_174), .A2(n_223), .B1(n_495), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_178), .A2(n_200), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_182), .A2(n_234), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_188), .A2(n_192), .B1(n_419), .B2(n_613), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_190), .A2(n_204), .B1(n_346), .B2(n_445), .Y(n_444) );
OA22x2_ASAP7_75t_L g558 ( .A1(n_193), .A2(n_559), .B1(n_577), .B2(n_578), .Y(n_558) );
INVx1_ASAP7_75t_L g577 ( .A(n_193), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_199), .A2(n_218), .B1(n_332), .B2(n_336), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_201), .B(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_203), .A2(n_246), .B1(n_417), .B2(n_420), .Y(n_517) );
AND2x4_ASAP7_75t_L g262 ( .A(n_205), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g674 ( .A(n_205), .Y(n_674) );
AO21x1_ASAP7_75t_L g683 ( .A1(n_205), .A2(n_258), .B(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_210), .A2(n_216), .B1(n_386), .B2(n_417), .Y(n_470) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
AND2x2_ASAP7_75t_R g710 ( .A(n_212), .B(n_674), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_215), .B(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_219), .A2(n_245), .B1(n_297), .B2(n_528), .Y(n_587) );
INVxp67_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_225), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_228), .A2(n_247), .B1(n_424), .B2(n_520), .Y(n_667) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_243), .B(n_523), .Y(n_522) );
AOI22x1_ASAP7_75t_L g653 ( .A1(n_251), .A2(n_654), .B1(n_668), .B2(n_669), .Y(n_653) );
INVx1_ASAP7_75t_L g669 ( .A(n_251), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_263), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g684 ( .A(n_263), .Y(n_684) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_433), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_265), .A2(n_433), .B(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_354), .B2(n_432), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_322), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_302), .Y(n_270) );
OAI21xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_291), .B(n_292), .Y(n_271) );
OAI21xp5_ASAP7_75t_SL g525 ( .A1(n_272), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx4_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx4_ASAP7_75t_SL g365 ( .A(n_274), .Y(n_365) );
BUFx2_ASAP7_75t_L g493 ( .A(n_274), .Y(n_493) );
INVx3_ASAP7_75t_SL g565 ( .A(n_274), .Y(n_565) );
INVx3_ASAP7_75t_L g623 ( .A(n_274), .Y(n_623) );
INVx6_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_284), .Y(n_275) );
AND2x4_ASAP7_75t_L g309 ( .A(n_276), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g320 ( .A(n_276), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g401 ( .A(n_276), .B(n_284), .Y(n_401) );
AND2x2_ASAP7_75t_L g413 ( .A(n_276), .B(n_321), .Y(n_413) );
AND2x2_ASAP7_75t_L g451 ( .A(n_276), .B(n_321), .Y(n_451) );
AND2x2_ASAP7_75t_L g465 ( .A(n_276), .B(n_310), .Y(n_465) );
AND2x2_ASAP7_75t_L g660 ( .A(n_276), .B(n_310), .Y(n_660) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_282), .Y(n_276) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g300 ( .A(n_277), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g317 ( .A(n_277), .Y(n_317) );
OAI22x1_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B1(n_280), .B2(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
INVx2_ASAP7_75t_L g287 ( .A(n_279), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_279), .Y(n_290) );
INVx2_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
AND2x2_ASAP7_75t_L g316 ( .A(n_282), .B(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g338 ( .A(n_282), .Y(n_338) );
AND2x4_ASAP7_75t_L g327 ( .A(n_284), .B(n_300), .Y(n_327) );
AND2x4_ASAP7_75t_L g344 ( .A(n_284), .B(n_330), .Y(n_344) );
AND2x2_ASAP7_75t_L g350 ( .A(n_284), .B(n_316), .Y(n_350) );
AND2x6_ASAP7_75t_L g419 ( .A(n_284), .B(n_316), .Y(n_419) );
AND2x2_ASAP7_75t_L g423 ( .A(n_284), .B(n_300), .Y(n_423) );
AND2x2_ASAP7_75t_L g520 ( .A(n_284), .B(n_300), .Y(n_520) );
AND2x2_ASAP7_75t_L g612 ( .A(n_284), .B(n_330), .Y(n_612) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_286), .B(n_289), .Y(n_295) );
AND2x4_ASAP7_75t_L g299 ( .A(n_286), .B(n_288), .Y(n_299) );
INVx1_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVxp67_ASAP7_75t_L g321 ( .A(n_288), .Y(n_321) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_289), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g626 ( .A(n_293), .Y(n_626) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g371 ( .A(n_294), .Y(n_371) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x4_ASAP7_75t_L g329 ( .A(n_295), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g337 ( .A(n_295), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_SL g398 ( .A(n_295), .B(n_296), .Y(n_398) );
AND2x4_ASAP7_75t_L g424 ( .A(n_295), .B(n_330), .Y(n_424) );
AND2x4_ASAP7_75t_L g427 ( .A(n_295), .B(n_338), .Y(n_427) );
BUFx5_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
BUFx3_ASAP7_75t_L g496 ( .A(n_298), .Y(n_496) );
INVx2_ASAP7_75t_L g705 ( .A(n_298), .Y(n_705) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g315 ( .A(n_299), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g346 ( .A(n_299), .B(n_330), .Y(n_346) );
AND2x4_ASAP7_75t_L g397 ( .A(n_299), .B(n_300), .Y(n_397) );
AND2x2_ASAP7_75t_L g410 ( .A(n_299), .B(n_316), .Y(n_410) );
AND2x2_ASAP7_75t_L g462 ( .A(n_299), .B(n_316), .Y(n_462) );
AND2x2_ASAP7_75t_L g613 ( .A(n_299), .B(n_330), .Y(n_613) );
AND2x2_ASAP7_75t_L g305 ( .A(n_300), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g464 ( .A(n_300), .B(n_306), .Y(n_464) );
AND2x4_ASAP7_75t_L g330 ( .A(n_301), .B(n_317), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_312), .Y(n_302) );
INVx1_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
BUFx6f_ASAP7_75t_SL g700 ( .A(n_304), .Y(n_700) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g502 ( .A(n_305), .Y(n_502) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_305), .Y(n_645) );
AND2x2_ASAP7_75t_L g335 ( .A(n_306), .B(n_316), .Y(n_335) );
AND2x4_ASAP7_75t_L g353 ( .A(n_306), .B(n_330), .Y(n_353) );
AND2x6_ASAP7_75t_L g420 ( .A(n_306), .B(n_330), .Y(n_420) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_306), .B(n_316), .Y(n_426) );
AND2x2_ASAP7_75t_L g516 ( .A(n_306), .B(n_316), .Y(n_516) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_307), .Y(n_311) );
BUFx4f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
INVx1_ASAP7_75t_L g406 ( .A(n_309), .Y(n_406) );
BUFx6f_ASAP7_75t_SL g454 ( .A(n_309), .Y(n_454) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx4f_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
BUFx2_ASAP7_75t_L g498 ( .A(n_314), .Y(n_498) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g533 ( .A(n_315), .Y(n_533) );
BUFx2_ASAP7_75t_L g641 ( .A(n_315), .Y(n_641) );
BUFx3_ASAP7_75t_L g717 ( .A(n_315), .Y(n_717) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx2_ASAP7_75t_L g499 ( .A(n_319), .Y(n_499) );
INVx2_ASAP7_75t_L g534 ( .A(n_319), .Y(n_534) );
INVx2_ASAP7_75t_SL g642 ( .A(n_319), .Y(n_642) );
INVx2_ASAP7_75t_SL g708 ( .A(n_319), .Y(n_708) );
INVx6_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_339), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_331), .Y(n_323) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
INVx1_ASAP7_75t_SL g489 ( .A(n_326), .Y(n_489) );
INVx2_ASAP7_75t_L g637 ( .A(n_326), .Y(n_637) );
INVx6_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g543 ( .A(n_327), .Y(n_543) );
BUFx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_SL g379 ( .A(n_329), .Y(n_379) );
INVx2_ASAP7_75t_L g545 ( .A(n_329), .Y(n_545) );
BUFx3_ASAP7_75t_L g638 ( .A(n_329), .Y(n_638) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
INVx1_ASAP7_75t_L g572 ( .A(n_334), .Y(n_572) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_335), .Y(n_441) );
BUFx3_ASAP7_75t_L g592 ( .A(n_335), .Y(n_592) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
BUFx3_ASAP7_75t_L g442 ( .A(n_337), .Y(n_442) );
INVx5_ASAP7_75t_SL g485 ( .A(n_337), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_347), .Y(n_339) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g417 ( .A(n_343), .Y(n_417) );
INVx2_ASAP7_75t_L g487 ( .A(n_343), .Y(n_487) );
INVx2_ASAP7_75t_SL g547 ( .A(n_343), .Y(n_547) );
INVx3_ASAP7_75t_SL g575 ( .A(n_343), .Y(n_575) );
INVx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_346), .Y(n_548) );
INVx2_ASAP7_75t_L g570 ( .A(n_346), .Y(n_570) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g539 ( .A(n_349), .Y(n_539) );
INVx2_ASAP7_75t_L g594 ( .A(n_349), .Y(n_594) );
INVx2_ASAP7_75t_SL g728 ( .A(n_349), .Y(n_728) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g481 ( .A(n_350), .Y(n_481) );
BUFx2_ASAP7_75t_L g696 ( .A(n_350), .Y(n_696) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
INVx2_ASAP7_75t_L g482 ( .A(n_352), .Y(n_482) );
INVx2_ASAP7_75t_L g540 ( .A(n_352), .Y(n_540) );
INVx2_ASAP7_75t_SL g576 ( .A(n_352), .Y(n_576) );
INVx2_ASAP7_75t_L g630 ( .A(n_352), .Y(n_630) );
INVx1_ASAP7_75t_SL g729 ( .A(n_352), .Y(n_729) );
INVx8_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g432 ( .A(n_354), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_389), .B2(n_429), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx5_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_376), .Y(n_358) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .C(n_366), .D(n_372), .Y(n_359) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g528 ( .A(n_371), .Y(n_528) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g701 ( .A(n_375), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .C(n_384), .D(n_387), .Y(n_376) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g633 ( .A(n_386), .Y(n_633) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
INVx1_ASAP7_75t_L g428 ( .A(n_393), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_414), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_402), .C(n_407), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_399), .Y(n_395) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_402) );
INVx2_ASAP7_75t_SL g503 ( .A(n_406), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_412), .Y(n_407) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_421), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g446 ( .A(n_419), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
XOR2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_553), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_473), .B1(n_550), .B2(n_552), .Y(n_434) );
INVx2_ASAP7_75t_L g551 ( .A(n_435), .Y(n_551) );
AO22x2_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_455), .B1(n_471), .B2(n_472), .Y(n_435) );
INVx1_ASAP7_75t_SL g471 ( .A(n_436), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_448), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .C(n_444), .D(n_447), .Y(n_439) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_441), .Y(n_693) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g568 ( .A(n_446), .Y(n_568) );
NAND4xp25_ASAP7_75t_SL g448 ( .A(n_449), .B(n_450), .C(n_452), .D(n_453), .Y(n_448) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_454), .Y(n_646) );
INVx2_ASAP7_75t_SL g472 ( .A(n_455), .Y(n_472) );
XNOR2x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .C(n_461), .D(n_463), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .C(n_469), .D(n_470), .Y(n_466) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g552 ( .A(n_474), .Y(n_552) );
OA22x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_505), .B1(n_506), .B2(n_549), .Y(n_474) );
INVx1_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
XOR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_504), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_490), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .C(n_486), .D(n_488), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g724 ( .A(n_485), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .C(n_497), .D(n_500), .Y(n_490) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g531 ( .A(n_502), .Y(n_531) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
XNOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_522), .Y(n_506) );
XNOR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .C(n_512), .D(n_513), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .C(n_518), .D(n_519), .Y(n_514) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_548), .Y(n_697) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
XOR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_651), .Y(n_553) );
AOI22xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_556), .B1(n_616), .B2(n_650), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_579), .B1(n_580), .B2(n_615), .Y(n_556) );
INVx2_ASAP7_75t_L g615 ( .A(n_557), .Y(n_615) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g578 ( .A(n_559), .Y(n_578) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .D(n_564), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .C(n_573), .D(n_574), .Y(n_566) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g722 ( .A(n_570), .Y(n_722) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
XNOR2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_597), .Y(n_580) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .C(n_587), .D(n_588), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .C(n_593), .D(n_595), .Y(n_589) );
BUFx2_ASAP7_75t_L g635 ( .A(n_592), .Y(n_635) );
BUFx2_ASAP7_75t_L g629 ( .A(n_594), .Y(n_629) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
XOR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
NAND2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_617), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_618), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_639), .Y(n_619) );
NOR3xp33_ASAP7_75t_SL g620 ( .A(n_621), .B(n_624), .C(n_627), .Y(n_620) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .C(n_634), .D(n_636), .Y(n_627) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .Y(n_639) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g668 ( .A(n_654), .Y(n_668) );
NAND2x1_ASAP7_75t_SL g654 ( .A(n_655), .B(n_661), .Y(n_654) );
NOR2xp67_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx3_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_673), .B(n_676), .Y(n_731) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_686), .B2(n_709), .C1(n_711), .C2(n_731), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp33_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_690), .B(n_698), .Y(n_689) );
NAND4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_694), .D(n_695), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .C(n_706), .D(n_707), .Y(n_698) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g719 ( .A(n_705), .Y(n_719) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g730 ( .A(n_713), .Y(n_730) );
NOR4xp75_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .C(n_720), .D(n_725), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
endmodule