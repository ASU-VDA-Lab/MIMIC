module fake_jpeg_24354_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_23),
.B1(n_11),
.B2(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_18),
.B(n_19),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_19),
.B(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_18),
.CI(n_23),
.CON(n_42),
.SN(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.C(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_21),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_25),
.B(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_54),
.B1(n_57),
.B2(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_11),
.B1(n_24),
.B2(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_44),
.B1(n_58),
.B2(n_48),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_25),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_37),
.C(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_69),
.C(n_47),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_37),
.C(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_55),
.B1(n_39),
.B2(n_43),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_9),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_72),
.B1(n_78),
.B2(n_26),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_50),
.B1(n_49),
.B2(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_67),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_61),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_70),
.C(n_64),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_82),
.B(n_85),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_68),
.B1(n_62),
.B2(n_69),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_86),
.B(n_15),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_78),
.C(n_29),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_22),
.B(n_16),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_74),
.C(n_71),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_28),
.C(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_86),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_5),
.B(n_1),
.C(n_2),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_6),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_96),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_7),
.C(n_10),
.D(n_0),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_94),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_0),
.Y(n_104)
);


endmodule