module real_aes_733_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g584 ( .A(n_0), .B(n_265), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_1), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g142 ( .A(n_2), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_3), .B(n_507), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g533 ( .A(n_4), .B(n_154), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_5), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_6), .B(n_161), .Y(n_257) );
INVx1_ASAP7_75t_L g526 ( .A(n_7), .Y(n_526) );
INVx1_ASAP7_75t_L g170 ( .A(n_8), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_9), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_10), .Y(n_187) );
AND2x2_ASAP7_75t_L g537 ( .A(n_11), .B(n_214), .Y(n_537) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g266 ( .A(n_14), .Y(n_266) );
AOI221x1_ASAP7_75t_L g529 ( .A1(n_15), .A2(n_128), .B1(n_506), .B2(n_530), .C(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_16), .B(n_507), .Y(n_515) );
INVx1_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
INVx1_ASAP7_75t_L g263 ( .A(n_18), .Y(n_263) );
INVx1_ASAP7_75t_SL g228 ( .A(n_19), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_20), .B(n_148), .Y(n_249) );
AOI33xp33_ASAP7_75t_L g199 ( .A1(n_21), .A2(n_52), .A3(n_137), .B1(n_146), .B2(n_200), .B3(n_201), .Y(n_199) );
AOI221xp5_ASAP7_75t_SL g505 ( .A1(n_22), .A2(n_40), .B1(n_506), .B2(n_507), .C(n_508), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_23), .A2(n_506), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_24), .B(n_265), .Y(n_542) );
INVx1_ASAP7_75t_L g179 ( .A(n_25), .Y(n_179) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_26), .A2(n_91), .B(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g162 ( .A(n_26), .B(n_91), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_27), .B(n_268), .Y(n_519) );
INVxp67_ASAP7_75t_L g528 ( .A(n_28), .Y(n_528) );
AND2x2_ASAP7_75t_L g573 ( .A(n_29), .B(n_213), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_30), .B(n_156), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_31), .A2(n_506), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_32), .B(n_268), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_33), .A2(n_43), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_33), .Y(n_787) );
INVx1_ASAP7_75t_L g136 ( .A(n_34), .Y(n_136) );
AND2x2_ASAP7_75t_L g154 ( .A(n_34), .B(n_142), .Y(n_154) );
AND2x2_ASAP7_75t_L g160 ( .A(n_34), .B(n_139), .Y(n_160) );
OR2x6_ASAP7_75t_L g110 ( .A(n_35), .B(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_36), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_37), .B(n_156), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_38), .A2(n_129), .B1(n_161), .B2(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_39), .B(n_251), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_41), .A2(n_82), .B1(n_134), .B2(n_506), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_42), .B(n_148), .Y(n_229) );
INVx1_ASAP7_75t_L g788 ( .A(n_43), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_44), .B(n_265), .Y(n_571) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_45), .A2(n_78), .B1(n_117), .B2(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_45), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_46), .B(n_167), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_47), .B(n_148), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_48), .Y(n_246) );
AND2x2_ASAP7_75t_L g587 ( .A(n_49), .B(n_213), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_50), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_51), .B(n_213), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_53), .B(n_148), .Y(n_211) );
INVx1_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
INVx1_ASAP7_75t_L g150 ( .A(n_54), .Y(n_150) );
AND2x2_ASAP7_75t_L g212 ( .A(n_55), .B(n_213), .Y(n_212) );
AOI221xp5_ASAP7_75t_L g168 ( .A1(n_56), .A2(n_74), .B1(n_134), .B2(n_156), .C(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_57), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_58), .B(n_507), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_59), .B(n_129), .Y(n_189) );
AOI21xp5_ASAP7_75t_SL g133 ( .A1(n_60), .A2(n_134), .B(n_143), .Y(n_133) );
AND2x2_ASAP7_75t_L g552 ( .A(n_61), .B(n_213), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_62), .B(n_268), .Y(n_585) );
INVx1_ASAP7_75t_L g260 ( .A(n_63), .Y(n_260) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_64), .B(n_214), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_65), .B(n_265), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_66), .A2(n_506), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g210 ( .A(n_67), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_68), .B(n_268), .Y(n_543) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_69), .B(n_167), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_70), .A2(n_90), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_70), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_71), .A2(n_134), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g152 ( .A(n_72), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_73), .B(n_156), .Y(n_202) );
AND2x2_ASAP7_75t_L g230 ( .A(n_75), .B(n_128), .Y(n_230) );
INVx1_ASAP7_75t_L g261 ( .A(n_76), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_77), .A2(n_134), .B(n_227), .Y(n_226) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_78), .A2(n_104), .B1(n_471), .B2(n_478), .C1(n_796), .C2(n_801), .Y(n_103) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_79), .A2(n_134), .B(n_194), .C(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_80), .B(n_507), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_81), .A2(n_85), .B1(n_156), .B2(n_507), .Y(n_556) );
INVx1_ASAP7_75t_L g113 ( .A(n_83), .Y(n_113) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_84), .B(n_128), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_86), .A2(n_134), .B1(n_197), .B2(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_87), .B(n_265), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_88), .B(n_265), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_89), .A2(n_506), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g466 ( .A(n_90), .Y(n_466) );
NOR2xp33_ASAP7_75t_SL g489 ( .A(n_90), .B(n_490), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_90), .A2(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_90), .A2(n_490), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
XNOR2xp5_ASAP7_75t_L g785 ( .A(n_93), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_94), .B(n_268), .Y(n_549) );
AND2x2_ASAP7_75t_L g203 ( .A(n_95), .B(n_128), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_96), .A2(n_177), .B(n_178), .C(n_181), .Y(n_176) );
INVxp67_ASAP7_75t_L g531 ( .A(n_97), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_98), .B(n_507), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_99), .B(n_268), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_100), .A2(n_506), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g477 ( .A(n_101), .Y(n_477) );
BUFx2_ASAP7_75t_SL g805 ( .A(n_101), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_102), .B(n_148), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B(n_468), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g470 ( .A(n_107), .Y(n_470) );
BUFx2_ASAP7_75t_L g807 ( .A(n_107), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x6_ASAP7_75t_SL g485 ( .A(n_108), .B(n_110), .Y(n_485) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_108), .B(n_109), .Y(n_784) );
OR2x2_ASAP7_75t_L g795 ( .A(n_108), .B(n_110), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B1(n_119), .B2(n_467), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g467 ( .A(n_119), .Y(n_467) );
XOR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_463), .Y(n_119) );
NAND3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_353), .C(n_418), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_307), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_252), .B(n_280), .Y(n_122) );
AOI21xp33_ASAP7_75t_SL g491 ( .A1(n_123), .A2(n_252), .B(n_280), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_215), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_163), .Y(n_124) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_125), .A2(n_355), .B(n_366), .Y(n_354) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_125), .B(n_296), .Y(n_389) );
AND2x2_ASAP7_75t_L g404 ( .A(n_125), .B(n_405), .Y(n_404) );
OR2x6_ASAP7_75t_L g414 ( .A(n_125), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g416 ( .A(n_125), .B(n_406), .Y(n_416) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g290 ( .A(n_126), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_126), .B(n_304), .Y(n_303) );
INVx4_ASAP7_75t_L g322 ( .A(n_126), .Y(n_322) );
AND2x2_ASAP7_75t_L g325 ( .A(n_126), .B(n_241), .Y(n_325) );
NOR2x1_ASAP7_75t_SL g328 ( .A(n_126), .B(n_256), .Y(n_328) );
AND2x4_ASAP7_75t_L g340 ( .A(n_126), .B(n_338), .Y(n_340) );
OR2x2_ASAP7_75t_L g350 ( .A(n_126), .B(n_222), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_126), .B(n_362), .Y(n_367) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_128), .A2(n_176), .B1(n_182), .B2(n_183), .Y(n_175) );
INVx3_ASAP7_75t_L g183 ( .A(n_128), .Y(n_183) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_129), .B(n_186), .Y(n_185) );
AOI21x1_ASAP7_75t_L g580 ( .A1(n_129), .A2(n_581), .B(n_587), .Y(n_580) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
AND2x4_ASAP7_75t_L g161 ( .A(n_131), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_131), .B(n_162), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_155), .B(n_161), .Y(n_132) );
INVxp67_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_134), .A2(n_156), .B1(n_525), .B2(n_527), .Y(n_524) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
NOR2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x6_ASAP7_75t_L g145 ( .A(n_138), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g265 ( .A(n_139), .B(n_149), .Y(n_265) );
AND2x6_ASAP7_75t_L g506 ( .A(n_140), .B(n_160), .Y(n_506) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
INVx2_ASAP7_75t_L g146 ( .A(n_141), .Y(n_146) );
AND2x4_ASAP7_75t_L g268 ( .A(n_141), .B(n_151), .Y(n_268) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_147), .C(n_153), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_145), .A2(n_153), .B(n_170), .C(n_171), .Y(n_169) );
INVxp67_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_145), .A2(n_153), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g227 ( .A1(n_145), .A2(n_153), .B(n_228), .C(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g251 ( .A(n_145), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_145), .A2(n_180), .B1(n_260), .B2(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g157 ( .A(n_146), .B(n_158), .Y(n_157) );
INVxp33_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AND2x4_ASAP7_75t_L g507 ( .A(n_148), .B(n_154), .Y(n_507) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_153), .A2(n_249), .B(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_153), .B(n_161), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_153), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_153), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_153), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_153), .A2(n_549), .B(n_550), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_153), .A2(n_570), .B(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_153), .A2(n_584), .B(n_585), .Y(n_583) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g244 ( .A(n_157), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_161), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_161), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_161), .B(n_531), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_161), .B(n_180), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_539), .B(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_163), .A2(n_296), .B1(n_391), .B2(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g434 ( .A(n_163), .Y(n_434) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_191), .Y(n_163) );
INVx2_ASAP7_75t_L g365 ( .A(n_164), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_164), .B(n_311), .Y(n_437) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_173), .Y(n_164) );
BUFx3_ASAP7_75t_L g283 ( .A(n_165), .Y(n_283) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g276 ( .A(n_166), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_166), .B(n_193), .Y(n_298) );
AND2x4_ASAP7_75t_L g315 ( .A(n_166), .B(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_L g331 ( .A(n_166), .Y(n_331) );
INVx2_ASAP7_75t_L g388 ( .A(n_166), .Y(n_388) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_172), .Y(n_166) );
INVx2_ASAP7_75t_SL g194 ( .A(n_167), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_167), .A2(n_515), .B(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g306 ( .A(n_173), .B(n_272), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_173), .B(n_275), .Y(n_352) );
AND2x2_ASAP7_75t_L g371 ( .A(n_173), .B(n_275), .Y(n_371) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g233 ( .A(n_174), .Y(n_233) );
INVx1_ASAP7_75t_L g314 ( .A(n_174), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_174), .B(n_205), .Y(n_333) );
AND2x4_ASAP7_75t_L g387 ( .A(n_174), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_184), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_183), .A2(n_206), .B(n_212), .Y(n_205) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_183), .A2(n_206), .B(n_212), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g346 ( .A(n_191), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_191), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_204), .Y(n_191) );
AND2x2_ASAP7_75t_L g330 ( .A(n_192), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g370 ( .A(n_192), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_192), .B(n_275), .Y(n_375) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_193), .B(n_205), .Y(n_235) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_203), .Y(n_193) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_194), .A2(n_195), .B(n_203), .Y(n_272) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_194), .A2(n_555), .B(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_196), .B(n_202), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g311 ( .A(n_204), .Y(n_311) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_204), .B(n_283), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_204), .B(n_233), .Y(n_450) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_205), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_213), .Y(n_223) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_213), .A2(n_505), .B(n_511), .Y(n_504) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OAI21xp33_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_231), .B(n_236), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_218), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
AND2x2_ASAP7_75t_L g302 ( .A(n_219), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g336 ( .A(n_219), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g402 ( .A(n_219), .B(n_320), .Y(n_402) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_219), .B(n_449), .C(n_450), .Y(n_448) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_220), .Y(n_279) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g295 ( .A(n_222), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_222), .B(n_256), .Y(n_301) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_222), .Y(n_312) );
AND2x2_ASAP7_75t_L g357 ( .A(n_222), .B(n_255), .Y(n_357) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_222), .Y(n_380) );
INVx1_ASAP7_75t_L g397 ( .A(n_222), .Y(n_397) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_230), .Y(n_222) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_223), .A2(n_546), .B(n_552), .Y(n_545) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_223), .A2(n_567), .B(n_573), .Y(n_566) );
AO21x2_ASAP7_75t_L g630 ( .A1(n_223), .A2(n_567), .B(n_573), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g439 ( .A(n_231), .Y(n_439) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_232), .B(n_310), .Y(n_411) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g273 ( .A(n_233), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI211x1_ASAP7_75t_L g307 ( .A1(n_237), .A2(n_308), .B(n_317), .C(n_334), .Y(n_307) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_238), .B(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g360 ( .A(n_238), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g296 ( .A(n_240), .B(n_255), .Y(n_296) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_L g254 ( .A(n_241), .B(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_241), .Y(n_321) );
INVx1_ASAP7_75t_L g338 ( .A(n_241), .Y(n_338) );
AND2x2_ASAP7_75t_L g406 ( .A(n_241), .B(n_256), .Y(n_406) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
NOR3xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .C(n_246), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_270), .B(n_277), .Y(n_252) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_253), .B(n_322), .Y(n_425) );
INVx2_ASAP7_75t_L g457 ( .A(n_253), .Y(n_457) );
INVx4_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g362 ( .A(n_255), .Y(n_362) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g304 ( .A(n_256), .Y(n_304) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B(n_269), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_266), .B2(n_267), .Y(n_262) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
OR2x2_ASAP7_75t_L g364 ( .A(n_271), .B(n_365), .Y(n_364) );
NAND2x1_ASAP7_75t_SL g386 ( .A(n_271), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g286 ( .A(n_272), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g316 ( .A(n_272), .Y(n_316) );
INVx1_ASAP7_75t_L g440 ( .A(n_273), .Y(n_440) );
AND2x2_ASAP7_75t_L g305 ( .A(n_274), .B(n_306), .Y(n_305) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
INVxp33_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g344 ( .A(n_279), .B(n_337), .Y(n_344) );
OAI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B(n_291), .C(n_299), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g368 ( .A(n_282), .B(n_369), .Y(n_368) );
NOR2xp67_ASAP7_75t_SL g373 ( .A(n_282), .B(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_283), .B(n_370), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_289), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x2_ASAP7_75t_L g417 ( .A(n_286), .B(n_387), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_289), .A2(n_436), .B1(n_438), .B2(n_441), .C1(n_442), .C2(n_445), .Y(n_435) );
INVx1_ASAP7_75t_L g399 ( .A(n_290), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_295), .Y(n_326) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_295), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g415 ( .A(n_296), .Y(n_415) );
AND2x2_ASAP7_75t_L g460 ( .A(n_296), .B(n_312), .Y(n_460) );
AND2x2_ASAP7_75t_L g341 ( .A(n_297), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g454 ( .A(n_298), .B(n_333), .Y(n_454) );
OAI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_305), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_300), .A2(n_320), .B(n_361), .Y(n_421) );
AND2x2_ASAP7_75t_L g445 ( .A(n_301), .B(n_322), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g455 ( .A(n_301), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g393 ( .A(n_304), .Y(n_393) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_304), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g428 ( .A(n_306), .Y(n_428) );
INVx1_ASAP7_75t_L g490 ( .A(n_307), .Y(n_490) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g431 ( .A(n_311), .B(n_315), .Y(n_431) );
BUFx2_ASAP7_75t_L g319 ( .A(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
INVx2_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
AND2x2_ASAP7_75t_L g384 ( .A(n_314), .B(n_375), .Y(n_384) );
AND2x4_ASAP7_75t_L g351 ( .A(n_315), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g391 ( .A(n_315), .B(n_348), .Y(n_391) );
AND2x2_ASAP7_75t_L g442 ( .A(n_315), .B(n_443), .Y(n_442) );
AOI31xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_323), .A3(n_327), .B(n_329), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g339 ( .A(n_319), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x4_ASAP7_75t_L g337 ( .A(n_322), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_325), .A2(n_377), .B1(n_408), .B2(n_411), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_325), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g462 ( .A(n_325), .B(n_378), .Y(n_462) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_378), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g400 ( .A(n_330), .B(n_371), .Y(n_400) );
INVx1_ASAP7_75t_L g410 ( .A(n_332), .Y(n_410) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_343), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B(n_341), .Y(n_335) );
INVx1_ASAP7_75t_L g433 ( .A(n_336), .Y(n_433) );
AND2x2_ASAP7_75t_L g441 ( .A(n_337), .B(n_393), .Y(n_441) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_337), .Y(n_447) );
AND2x2_ASAP7_75t_L g392 ( .A(n_340), .B(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_345), .B1(n_349), .B2(n_351), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_346), .A2(n_365), .B1(n_459), .B2(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g358 ( .A(n_351), .Y(n_358) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_353), .B(n_418), .C(n_489), .D(n_491), .Y(n_488) );
INVxp67_ASAP7_75t_L g493 ( .A(n_353), .Y(n_493) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_381), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_357), .A2(n_360), .B(n_363), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g383 ( .A1(n_360), .A2(n_384), .B1(n_385), .B2(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_372), .B2(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_382), .B(n_394), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .Y(n_382) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NAND2xp33_ASAP7_75t_SL g436 ( .A(n_386), .B(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g409 ( .A(n_387), .Y(n_409) );
INVx3_ASAP7_75t_L g423 ( .A(n_391), .Y(n_423) );
INVxp67_ASAP7_75t_L g452 ( .A(n_392), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_403), .C(n_407), .D(n_412), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g405 ( .A(n_397), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
NAND2xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_416), .B(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
AND3x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_435), .C(n_446), .Y(n_418) );
AOI221x1_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_432), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp33_ASAP7_75t_SL g426 ( .A(n_427), .B(n_430), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
NAND2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI211xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_451), .C(n_458), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_451) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g797 ( .A(n_470), .B(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_SL g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g800 ( .A(n_475), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_475), .A2(n_803), .B(n_806), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g799 ( .A(n_477), .B(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_785), .B(n_789), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_486), .B(n_497), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_482), .A2(n_487), .B1(n_498), .B2(n_791), .Y(n_790) );
CKINVDCx6p67_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .C(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g494 ( .A(n_491), .Y(n_494) );
NAND2x1_ASAP7_75t_SL g497 ( .A(n_498), .B(n_780), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_693), .Y(n_499) );
NAND3xp33_ASAP7_75t_SL g500 ( .A(n_501), .B(n_603), .C(n_643), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_521), .B(n_534), .C(n_559), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_502), .B(n_608), .Y(n_642) );
NOR2x1p5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
INVx2_ASAP7_75t_L g594 ( .A(n_504), .Y(n_594) );
OR2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_513), .Y(n_606) );
AND2x2_ASAP7_75t_L g620 ( .A(n_504), .B(n_579), .Y(n_620) );
INVx1_ASAP7_75t_L g648 ( .A(n_504), .Y(n_648) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_504), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_504), .B(n_513), .Y(n_754) );
OR2x2_ASAP7_75t_L g575 ( .A(n_512), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_512), .Y(n_710) );
AND2x2_ASAP7_75t_L g715 ( .A(n_512), .B(n_577), .Y(n_715) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g521 ( .A(n_513), .B(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g574 ( .A(n_513), .B(n_523), .Y(n_574) );
OR2x2_ASAP7_75t_L g593 ( .A(n_513), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g622 ( .A(n_513), .Y(n_622) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_513), .B(n_523), .Y(n_661) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_513), .Y(n_665) );
OR2x2_ASAP7_75t_L g682 ( .A(n_513), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g692 ( .A(n_513), .B(n_599), .Y(n_692) );
INVx1_ASAP7_75t_L g721 ( .A(n_513), .Y(n_721) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_521), .B(n_650), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_522), .B(n_579), .Y(n_596) );
AND2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_593), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_522), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g599 ( .A(n_523), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g621 ( .A(n_523), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g656 ( .A(n_523), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_523), .B(n_579), .Y(n_680) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_535), .B(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g629 ( .A(n_535), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_535), .B(n_545), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_535), .B(n_650), .C(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g697 ( .A(n_535), .B(n_602), .Y(n_697) );
INVx5_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g564 ( .A(n_536), .B(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_536), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g617 ( .A(n_536), .Y(n_617) );
OR2x2_ASAP7_75t_L g640 ( .A(n_536), .B(n_630), .Y(n_640) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_536), .Y(n_657) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_536), .B(n_563), .Y(n_675) );
AND2x4_ASAP7_75t_L g690 ( .A(n_536), .B(n_566), .Y(n_690) );
AND2x2_ASAP7_75t_L g704 ( .A(n_536), .B(n_545), .Y(n_704) );
OR2x2_ASAP7_75t_L g725 ( .A(n_536), .B(n_553), .Y(n_725) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g779 ( .A(n_544), .B(n_657), .Y(n_779) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
AND2x4_ASAP7_75t_L g602 ( .A(n_545), .B(n_565), .Y(n_602) );
INVx2_ASAP7_75t_L g613 ( .A(n_545), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_545), .B(n_563), .Y(n_618) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_545), .Y(n_651) );
OR2x2_ASAP7_75t_L g674 ( .A(n_545), .B(n_566), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_545), .B(n_566), .Y(n_677) );
INVx1_ASAP7_75t_L g686 ( .A(n_545), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
AND2x2_ASAP7_75t_L g589 ( .A(n_553), .B(n_566), .Y(n_589) );
BUFx2_ASAP7_75t_L g638 ( .A(n_553), .Y(n_638) );
AND2x2_ASAP7_75t_L g733 ( .A(n_553), .B(n_613), .Y(n_733) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_554), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_574), .B1(n_575), .B2(n_588), .C(n_590), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_562), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_562), .B(n_629), .Y(n_669) );
OR2x2_ASAP7_75t_L g681 ( .A(n_562), .B(n_677), .Y(n_681) );
OR2x2_ASAP7_75t_L g684 ( .A(n_562), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g773 ( .A(n_562), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g612 ( .A(n_563), .B(n_613), .Y(n_612) );
OA33x2_ASAP7_75t_L g645 ( .A1(n_563), .A2(n_606), .A3(n_646), .B1(n_649), .B2(n_652), .B3(n_655), .Y(n_645) );
OR2x2_ASAP7_75t_L g676 ( .A(n_563), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g700 ( .A(n_563), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g708 ( .A(n_563), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g728 ( .A(n_563), .B(n_602), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_563), .B(n_617), .Y(n_766) );
INVx2_ASAP7_75t_L g636 ( .A(n_564), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g706 ( .A1(n_564), .A2(n_619), .A3(n_707), .B1(n_710), .B2(n_711), .C1(n_713), .C2(n_715), .Y(n_706) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_566), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
OR2x2_ASAP7_75t_L g688 ( .A(n_574), .B(n_667), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_574), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g761 ( .A(n_574), .Y(n_761) );
INVx1_ASAP7_75t_SL g627 ( .A(n_575), .Y(n_627) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g660 ( .A(n_577), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
INVx1_ASAP7_75t_L g609 ( .A(n_579), .Y(n_609) );
INVx1_ASAP7_75t_L g650 ( .A(n_579), .Y(n_650) );
OR2x2_ASAP7_75t_L g667 ( .A(n_579), .B(n_594), .Y(n_667) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_579), .Y(n_742) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_589), .B(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_597), .B(n_601), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_591), .A2(n_665), .B(n_666), .C(n_668), .Y(n_664) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_594), .Y(n_598) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g753 ( .A(n_596), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_SL g722 ( .A(n_599), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_599), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_599), .B(n_721), .Y(n_738) );
INVx3_ASAP7_75t_SL g663 ( .A(n_602), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_610), .B1(n_614), .B2(n_619), .C(n_623), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_609), .Y(n_654) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_612), .A2(n_639), .B(n_711), .Y(n_717) );
AND2x2_ASAP7_75t_L g743 ( .A(n_612), .B(n_690), .Y(n_743) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_613), .Y(n_631) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_617), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g752 ( .A(n_617), .B(n_674), .Y(n_752) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g701 ( .A(n_620), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_628), .B(n_632), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx2_ASAP7_75t_L g774 ( .A(n_629), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_630), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g703 ( .A(n_630), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_631), .B(n_653), .Y(n_652) );
OAI31xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_635), .A3(n_637), .B(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_636), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g714 ( .A(n_638), .B(n_640), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_638), .B(n_690), .Y(n_769) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR5xp2_ASAP7_75t_L g643 ( .A(n_644), .B(n_658), .C(n_670), .D(n_679), .E(n_687), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_648), .B(n_650), .Y(n_683) );
INVx1_ASAP7_75t_L g723 ( .A(n_648), .Y(n_723) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_648), .Y(n_760) );
INVx1_ASAP7_75t_L g712 ( .A(n_651), .Y(n_712) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OAI321xp33_ASAP7_75t_L g695 ( .A1(n_656), .A2(n_696), .A3(n_698), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_695) );
INVx1_ASAP7_75t_L g749 ( .A(n_657), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_660), .A2(n_733), .B1(n_740), .B2(n_743), .Y(n_739) );
AND2x2_ASAP7_75t_L g768 ( .A(n_661), .B(n_742), .Y(n_768) );
INVx1_ASAP7_75t_L g678 ( .A(n_666), .Y(n_678) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_676), .B(n_678), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_677), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g750 ( .A(n_677), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B1(n_682), .B2(n_684), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_686), .B(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_688), .A2(n_765), .B1(n_767), .B2(n_769), .C(n_770), .Y(n_764) );
INVx1_ASAP7_75t_L g771 ( .A(n_688), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_689), .A2(n_746), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_691), .A2(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_744), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_716), .C(n_734), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_697), .Y(n_763) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g762 ( .A(n_705), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_707), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g755 ( .A(n_715), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_724), .B(n_726), .Y(n_718) );
INVxp67_ASAP7_75t_L g776 ( .A(n_719), .Y(n_776) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g731 ( .A(n_722), .Y(n_731) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_739), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g777 ( .A(n_740), .Y(n_777) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_764), .C(n_775), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI21xp5_ASAP7_75t_SL g756 ( .A1(n_757), .A2(n_762), .B(n_763), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_768), .A2(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_778), .Y(n_775) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
BUFx4f_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g791 ( .A(n_783), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
AOI21xp33_ASAP7_75t_SL g789 ( .A1(n_785), .A2(n_790), .B(n_792), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx4f_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
CKINVDCx8_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
endmodule