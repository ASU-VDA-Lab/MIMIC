module fake_jpeg_24463_n_29 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.C(n_1),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_18),
.B(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_19),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

AOI32xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_1),
.A3(n_3),
.B1(n_5),
.B2(n_10),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_5),
.B(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI321xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.A3(n_25),
.B1(n_21),
.B2(n_22),
.C(n_16),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_18),
.C(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_25),
.Y(n_29)
);


endmodule