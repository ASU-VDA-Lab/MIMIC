module fake_jpeg_17890_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_12),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_58),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_42),
.B1(n_46),
.B2(n_44),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_42),
.B1(n_41),
.B2(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_46),
.B1(n_51),
.B2(n_37),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_37),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

AO21x2_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_70),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_45),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_68),
.B(n_5),
.C(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_3),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_92),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_85),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_4),
.B(n_8),
.C(n_10),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_98),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_16),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_94),
.B(n_95),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_92),
.B(n_79),
.C(n_84),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_107),
.B(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_92),
.B1(n_74),
.B2(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_114),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_102),
.C(n_100),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_106),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_115),
.B(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_17),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_21),
.B(n_23),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_26),
.B(n_29),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_30),
.Y(n_126)
);


endmodule