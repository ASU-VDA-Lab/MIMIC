module fake_jpeg_8322_n_224 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_3),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_28),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_22),
.C(n_32),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_58),
.C(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_19),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_18),
.B1(n_34),
.B2(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_51),
.Y(n_107)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_86),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_38),
.B1(n_23),
.B2(n_33),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_88),
.B(n_52),
.Y(n_98)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_90),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_41),
.B1(n_43),
.B2(n_19),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_79),
.B(n_77),
.C(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_13),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_33),
.B1(n_29),
.B2(n_19),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_19),
.B1(n_29),
.B2(n_41),
.Y(n_112)
);

NOR2x1p5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_48),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_98),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_48),
.B1(n_57),
.B2(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_110),
.B1(n_112),
.B2(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_51),
.B(n_55),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_49),
.B1(n_55),
.B2(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_29),
.B1(n_43),
.B2(n_28),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_43),
.C(n_4),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_84),
.C(n_4),
.Y(n_124)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_85),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_130),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_112),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_138),
.B(n_117),
.Y(n_145)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_89),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_129),
.C(n_141),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_135),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_101),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_13),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_16),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_86),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_82),
.C(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_74),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_108),
.B1(n_104),
.B2(n_111),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_140),
.B(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_132),
.B(n_135),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_116),
.B1(n_114),
.B2(n_105),
.C(n_110),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.C(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_98),
.C(n_116),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_137),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_103),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_103),
.B1(n_108),
.B2(n_73),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_131),
.B1(n_130),
.B2(n_136),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_111),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_165),
.B(n_169),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_138),
.B(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_177),
.C(n_155),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_132),
.B(n_120),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_170),
.A2(n_173),
.B(n_153),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_129),
.C(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_175),
.C(n_152),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_148),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_124),
.C(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_184),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_185),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_156),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_188),
.B(n_190),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_143),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_146),
.B1(n_157),
.B2(n_154),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_191),
.A2(n_172),
.B1(n_175),
.B2(n_177),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_165),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_162),
.B1(n_179),
.B2(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_196),
.B1(n_201),
.B2(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_167),
.B1(n_174),
.B2(n_168),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_146),
.B1(n_154),
.B2(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_206),
.Y(n_211)
);

HB1xp67_ASAP7_75t_SL g213 ( 
.A(n_203),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_205),
.B(n_207),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_183),
.B1(n_181),
.B2(n_191),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_16),
.B1(n_15),
.B2(n_6),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_3),
.C(n_5),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_197),
.B(n_7),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_199),
.C(n_196),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_194),
.B(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_6),
.B(n_7),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_203),
.Y(n_214)
);

AOI211xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_216),
.B(n_217),
.C(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_208),
.B1(n_202),
.B2(n_200),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NOR4xp25_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.C(n_12),
.D(n_8),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_193),
.B1(n_8),
.B2(n_9),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.C(n_11),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_7),
.B(n_9),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_11),
.Y(n_224)
);


endmodule