module real_aes_8682_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_555;
wire n_766;
wire n_1113;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1123;
wire n_549;
wire n_571;
wire n_491;
wire n_694;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_976;
wire n_1110;
wire n_752;
wire n_448;
wire n_1137;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_938;
wire n_384;
wire n_744;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_1049;
wire n_466;
wire n_559;
wire n_636;
wire n_1053;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_1017;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_598;
wire n_713;
wire n_1073;
wire n_404;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_1136;
wire n_1003;
wire n_533;
wire n_699;
wire n_1000;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_385;
wire n_649;
wire n_1056;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_1127;
wire n_968;
wire n_435;
wire n_972;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1114;
wire n_1045;
wire n_465;
wire n_566;
wire n_473;
wire n_837;
wire n_719;
wire n_871;
wire n_967;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_601;
wire n_500;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_0), .A2(n_194), .B1(n_474), .B2(n_702), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_1), .B(n_907), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g808 ( .A1(n_2), .A2(n_247), .B1(n_626), .B2(n_809), .Y(n_808) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_3), .A2(n_185), .B1(n_334), .B2(n_424), .C1(n_600), .C2(n_601), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_4), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_5), .A2(n_110), .B1(n_707), .B2(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_6), .A2(n_166), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_7), .A2(n_100), .B1(n_536), .B2(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_8), .B(n_554), .Y(n_553) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_9), .A2(n_232), .B1(n_407), .B2(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g1085 ( .A(n_9), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_10), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_11), .A2(n_177), .B1(n_478), .B2(n_572), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_12), .A2(n_360), .B1(n_433), .B2(n_597), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_13), .A2(n_174), .B1(n_483), .B2(n_701), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_14), .A2(n_163), .B1(n_575), .B2(n_676), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_15), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1136 ( .A(n_16), .Y(n_1136) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_17), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_18), .A2(n_202), .B1(n_551), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_19), .A2(n_114), .B1(n_532), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_20), .A2(n_258), .B1(n_676), .B2(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_21), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_22), .A2(n_322), .B1(n_483), .B2(n_532), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_23), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_24), .A2(n_308), .B1(n_734), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_25), .A2(n_239), .B1(n_490), .B2(n_494), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g1105 ( .A1(n_26), .A2(n_309), .B1(n_467), .B2(n_487), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_27), .Y(n_638) );
AOI22xp5_ASAP7_75t_SL g878 ( .A1(n_28), .A2(n_255), .B1(n_575), .B2(n_747), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_29), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_30), .A2(n_307), .B1(n_734), .B2(n_1030), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_31), .A2(n_262), .B1(n_478), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_32), .A2(n_366), .B1(n_569), .B2(n_935), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_33), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_34), .A2(n_253), .B1(n_539), .B2(n_572), .Y(n_773) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_35), .A2(n_129), .B1(n_407), .B2(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_36), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_37), .A2(n_180), .B1(n_488), .B2(n_495), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_38), .A2(n_941), .B1(n_960), .B2(n_961), .Y(n_940) );
INVx1_ASAP7_75t_L g961 ( .A(n_38), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_39), .A2(n_64), .B1(n_461), .B2(n_539), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_40), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_41), .A2(n_68), .B1(n_478), .B2(n_491), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_42), .A2(n_72), .B1(n_568), .B2(n_870), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_43), .A2(n_292), .B1(n_601), .B2(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_44), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_45), .A2(n_69), .B1(n_480), .B2(n_585), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_46), .A2(n_170), .B1(n_572), .B2(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_47), .B(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_48), .A2(n_302), .B1(n_626), .B2(n_707), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_49), .A2(n_132), .B1(n_631), .B2(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_50), .B(n_551), .Y(n_1063) );
INVx1_ASAP7_75t_L g725 ( .A(n_51), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_52), .A2(n_368), .B1(n_598), .B2(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_53), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g1088 ( .A(n_54), .B(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_55), .A2(n_323), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_56), .A2(n_298), .B1(n_595), .B2(n_721), .Y(n_754) );
AOI22xp5_ASAP7_75t_SL g877 ( .A1(n_57), .A2(n_316), .B1(n_574), .B2(n_672), .Y(n_877) );
AOI222xp33_ASAP7_75t_L g1040 ( .A1(n_58), .A2(n_299), .B1(n_321), .B2(n_615), .C1(n_691), .C2(n_854), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1131 ( .A(n_59), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_60), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_61), .Y(n_602) );
AOI22xp5_ASAP7_75t_SL g819 ( .A1(n_62), .A2(n_230), .B1(n_672), .B2(n_676), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1096 ( .A1(n_63), .A2(n_82), .B1(n_431), .B2(n_617), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_65), .Y(n_1004) );
CKINVDCx16_ASAP7_75t_R g996 ( .A(n_66), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_67), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_70), .B(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_71), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_73), .A2(n_260), .B1(n_734), .B2(n_1123), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_74), .A2(n_99), .B1(n_560), .B2(n_601), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_75), .Y(n_636) );
INVx1_ASAP7_75t_L g439 ( .A(n_76), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_77), .A2(n_137), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_78), .A2(n_351), .B1(n_474), .B2(n_478), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_79), .A2(n_156), .B1(n_487), .B2(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_80), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_81), .A2(n_211), .B1(n_628), .B2(n_752), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_83), .A2(n_226), .B1(n_552), .B2(n_770), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_84), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_85), .A2(n_236), .B1(n_526), .B2(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g797 ( .A(n_86), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_87), .A2(n_104), .B1(n_812), .B2(n_862), .Y(n_861) );
AOI22xp5_ASAP7_75t_SL g822 ( .A1(n_88), .A2(n_106), .B1(n_539), .B2(n_823), .Y(n_822) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_89), .A2(n_266), .B1(n_407), .B2(n_408), .Y(n_414) );
INVx1_ASAP7_75t_L g1082 ( .A(n_89), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_90), .A2(n_91), .B1(n_711), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_92), .A2(n_354), .B1(n_925), .B2(n_926), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_93), .A2(n_352), .B1(n_591), .B2(n_730), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_94), .A2(n_372), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_95), .A2(n_294), .B1(n_907), .B2(n_948), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_96), .A2(n_376), .B1(n_536), .B2(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_97), .A2(n_223), .B1(n_693), .B2(n_854), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_98), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_101), .A2(n_288), .B1(n_490), .B2(n_494), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_102), .A2(n_312), .B1(n_566), .B2(n_585), .Y(n_936) );
OA22x2_ASAP7_75t_L g1025 ( .A1(n_103), .A2(n_1026), .B1(n_1027), .B2(n_1041), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_103), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_105), .A2(n_213), .B1(n_626), .B2(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_107), .A2(n_122), .B1(n_539), .B2(n_564), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_108), .A2(n_116), .B1(n_597), .B2(n_615), .Y(n_768) );
INVx1_ASAP7_75t_L g816 ( .A(n_109), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_111), .A2(n_244), .B1(n_674), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_112), .A2(n_136), .B1(n_538), .B2(n_640), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_113), .A2(n_345), .B1(n_598), .B2(n_975), .Y(n_1066) );
INVx1_ASAP7_75t_L g1137 ( .A(n_115), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g976 ( .A1(n_117), .A2(n_220), .B1(n_977), .B2(n_978), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_118), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_119), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_120), .B(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_121), .A2(n_148), .B1(n_483), .B2(n_486), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_123), .A2(n_284), .B1(n_671), .B2(n_672), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_124), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_125), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_126), .A2(n_283), .B1(n_626), .B2(n_805), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_127), .Y(n_991) );
INVx1_ASAP7_75t_L g666 ( .A(n_128), .Y(n_666) );
INVx1_ASAP7_75t_L g1086 ( .A(n_129), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_130), .A2(n_153), .B1(n_494), .B2(n_1033), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_131), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_133), .A2(n_209), .B1(n_558), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_134), .A2(n_138), .B1(n_626), .B2(n_674), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_135), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_135), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_139), .Y(n_829) );
XNOR2x2_ASAP7_75t_L g894 ( .A(n_140), .B(n_895), .Y(n_894) );
AOI211xp5_ASAP7_75t_L g998 ( .A1(n_141), .A2(n_691), .B(n_999), .C(n_1003), .Y(n_998) );
INVx1_ASAP7_75t_L g679 ( .A(n_142), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_143), .A2(n_203), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g736 ( .A(n_144), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_145), .A2(n_200), .B1(n_628), .B2(n_752), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_146), .A2(n_179), .B1(n_564), .B2(n_586), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_147), .A2(n_336), .B1(n_624), .B2(n_678), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_149), .A2(n_264), .B1(n_598), .B2(n_617), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_150), .A2(n_249), .B1(n_461), .B2(n_467), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g983 ( .A1(n_151), .A2(n_229), .B1(n_591), .B2(n_984), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g993 ( .A(n_152), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_154), .A2(n_362), .B1(n_433), .B2(n_597), .Y(n_723) );
AOI211xp5_ASAP7_75t_L g985 ( .A1(n_155), .A2(n_640), .B(n_986), .C(n_992), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_157), .A2(n_270), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_158), .A2(n_191), .B1(n_491), .B2(n_495), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_159), .A2(n_361), .B1(n_950), .B2(n_975), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_160), .A2(n_279), .B1(n_561), .B2(n_975), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_161), .A2(n_241), .B1(n_490), .B2(n_959), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_162), .Y(n_609) );
AND2x6_ASAP7_75t_L g387 ( .A(n_164), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_164), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_165), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_167), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_168), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_169), .A2(n_265), .B1(n_441), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_171), .A2(n_356), .B1(n_491), .B2(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_172), .A2(n_246), .B1(n_561), .B2(n_601), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_173), .A2(n_374), .B1(n_539), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_175), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g758 ( .A1(n_176), .A2(n_195), .B1(n_215), .B2(n_600), .C1(n_617), .C2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_178), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_181), .A2(n_378), .B1(n_442), .B2(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g685 ( .A(n_182), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_183), .Y(n_641) );
INVx1_ASAP7_75t_L g801 ( .A(n_184), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_186), .A2(n_192), .B1(n_487), .B2(n_674), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_187), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_188), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_189), .A2(n_272), .B1(n_483), .B2(n_635), .Y(n_1104) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_190), .A2(n_256), .B1(n_407), .B2(n_411), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g1083 ( .A(n_190), .B(n_1084), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_193), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_196), .A2(n_271), .B1(n_574), .B2(n_575), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_197), .A2(n_259), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI222xp33_ASAP7_75t_L g909 ( .A1(n_198), .A2(n_231), .B1(n_293), .B2(n_433), .C1(n_617), .C2(n_759), .Y(n_909) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_199), .A2(n_348), .B1(n_586), .B2(n_676), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_201), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_204), .A2(n_381), .B1(n_433), .B2(n_617), .Y(n_798) );
INVx1_ASAP7_75t_L g793 ( .A(n_205), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_206), .Y(n_972) );
INVx1_ASAP7_75t_L g800 ( .A(n_207), .Y(n_800) );
AOI22xp5_ASAP7_75t_SL g880 ( .A1(n_208), .A2(n_281), .B1(n_825), .B2(n_881), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_210), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_212), .A2(n_324), .B1(n_490), .B2(n_494), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_214), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_216), .B(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_217), .A2(n_353), .B1(n_560), .B2(n_975), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_218), .B(n_441), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1128 ( .A(n_219), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1100 ( .A1(n_221), .A2(n_257), .B1(n_950), .B2(n_975), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_222), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_224), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_225), .A2(n_269), .B1(n_591), .B2(n_823), .Y(n_1120) );
INVx1_ASAP7_75t_L g429 ( .A(n_227), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_228), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_233), .A2(n_504), .B1(n_540), .B2(n_541), .Y(n_503) );
INVx1_ASAP7_75t_L g540 ( .A(n_233), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_234), .A2(n_357), .B1(n_624), .B2(n_678), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_235), .B(n_551), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_237), .A2(n_297), .B1(n_756), .B2(n_950), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_238), .A2(n_371), .B1(n_487), .B2(n_591), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_240), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_242), .A2(n_296), .B1(n_469), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_243), .Y(n_1060) );
AOI22xp5_ASAP7_75t_SL g397 ( .A1(n_245), .A2(n_398), .B1(n_498), .B2(n_499), .Y(n_397) );
INVx1_ASAP7_75t_L g499 ( .A(n_245), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_248), .A2(n_377), .B1(n_628), .B2(n_631), .Y(n_627) );
INVx2_ASAP7_75t_L g391 ( .A(n_250), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_251), .A2(n_330), .B1(n_433), .B2(n_443), .Y(n_548) );
INVx1_ASAP7_75t_L g1114 ( .A(n_252), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1115 ( .A1(n_252), .A2(n_1114), .B1(n_1116), .B2(n_1138), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_254), .Y(n_968) );
INVx1_ASAP7_75t_L g401 ( .A(n_261), .Y(n_401) );
INVx1_ASAP7_75t_L g451 ( .A(n_263), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_267), .A2(n_314), .B1(n_568), .B2(n_959), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_268), .A2(n_363), .B1(n_709), .B2(n_711), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_273), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_274), .A2(n_380), .B1(n_631), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_275), .A2(n_350), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_276), .A2(n_310), .B1(n_750), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_277), .A2(n_320), .B1(n_948), .B2(n_977), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_278), .A2(n_291), .B1(n_469), .B2(n_566), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_280), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_282), .A2(n_319), .B1(n_467), .B2(n_1049), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_285), .Y(n_830) );
INVx1_ASAP7_75t_L g407 ( .A(n_286), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_286), .Y(n_409) );
INVx1_ASAP7_75t_L g794 ( .A(n_287), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_289), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_290), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_295), .A2(n_340), .B1(n_564), .B2(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_300), .Y(n_837) );
INVx1_ASAP7_75t_L g687 ( .A(n_301), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_303), .A2(n_383), .B(n_392), .C(n_1087), .Y(n_382) );
INVx1_ASAP7_75t_L g1127 ( .A(n_304), .Y(n_1127) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_305), .A2(n_349), .B1(n_558), .B2(n_560), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_306), .B(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_311), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_313), .A2(n_341), .B1(n_597), .B2(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g1099 ( .A(n_315), .B(n_770), .Y(n_1099) );
AO22x2_ASAP7_75t_L g916 ( .A1(n_317), .A2(n_917), .B1(n_938), .B2(n_939), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_317), .Y(n_939) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_318), .A2(n_343), .B1(n_431), .B2(n_616), .Y(n_1061) );
INVx1_ASAP7_75t_L g390 ( .A(n_325), .Y(n_390) );
AOI22xp5_ASAP7_75t_SL g681 ( .A1(n_326), .A2(n_682), .B1(n_712), .B2(n_713), .Y(n_681) );
INVx1_ASAP7_75t_L g713 ( .A(n_326), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_327), .A2(n_335), .B1(n_484), .B2(n_711), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g1053 ( .A(n_328), .Y(n_1053) );
INVx1_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_331), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_332), .B(n_595), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_333), .B(n_978), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_337), .Y(n_514) );
AOI22xp5_ASAP7_75t_SL g605 ( .A1(n_338), .A2(n_606), .B1(n_645), .B2(n_646), .Y(n_605) );
INVx1_ASAP7_75t_L g646 ( .A(n_338), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_339), .B(n_907), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_342), .A2(n_358), .B1(n_756), .B2(n_766), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_344), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_346), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_347), .Y(n_593) );
INVx1_ASAP7_75t_L g1019 ( .A(n_355), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_359), .B(n_595), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_364), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_365), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_367), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_369), .A2(n_1044), .B1(n_1045), .B2(n_1067), .Y(n_1043) );
INVx1_ASAP7_75t_L g1067 ( .A(n_369), .Y(n_1067) );
INVx1_ASAP7_75t_L g446 ( .A(n_370), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g964 ( .A(n_373), .B(n_965), .Y(n_964) );
OA22x2_ASAP7_75t_L g840 ( .A1(n_375), .A2(n_841), .B1(n_842), .B2(n_871), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_375), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_379), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_388), .Y(n_1078) );
OAI21xp5_ASAP7_75t_L g1112 ( .A1(n_389), .A2(n_1077), .B(n_1113), .Y(n_1112) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_651), .B1(n_1072), .B2(n_1073), .C(n_1074), .Y(n_392) );
INVx1_ASAP7_75t_L g1073 ( .A(n_393), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_500), .B2(n_501), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g498 ( .A(n_398), .Y(n_498) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_458), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_422), .C(n_445), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_417), .B2(n_418), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g831 ( .A1(n_402), .A2(n_832), .B(n_833), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_402), .A2(n_511), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g509 ( .A(n_403), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g608 ( .A1(n_403), .A2(n_511), .B1(n_609), .B2(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_412), .Y(n_403) );
INVx2_ASAP7_75t_L g477 ( .A(n_404), .Y(n_477) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_410), .Y(n_404) );
AND2x2_ASAP7_75t_L g421 ( .A(n_405), .B(n_410), .Y(n_421) );
AND2x2_ASAP7_75t_L g466 ( .A(n_405), .B(n_437), .Y(n_466) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g426 ( .A(n_406), .B(n_410), .Y(n_426) );
AND2x2_ASAP7_75t_L g438 ( .A(n_406), .B(n_416), .Y(n_438) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_409), .Y(n_411) );
INVx2_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVx1_ASAP7_75t_L g497 ( .A(n_410), .Y(n_497) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_413), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g488 ( .A(n_413), .B(n_466), .Y(n_488) );
AND2x6_ASAP7_75t_L g552 ( .A(n_413), .B(n_421), .Y(n_552) );
AND2x4_ASAP7_75t_L g556 ( .A(n_413), .B(n_477), .Y(n_556) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
INVx1_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_414), .B(n_416), .Y(n_472) );
AND2x2_ASAP7_75t_L g427 ( .A(n_415), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g465 ( .A(n_416), .B(n_457), .Y(n_465) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g828 ( .A(n_419), .Y(n_828) );
INVx1_ASAP7_75t_L g905 ( .A(n_419), .Y(n_905) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g511 ( .A(n_420), .Y(n_511) );
AND2x4_ASAP7_75t_L g480 ( .A(n_421), .B(n_427), .Y(n_480) );
AND2x2_ASAP7_75t_L g493 ( .A(n_421), .B(n_465), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g988 ( .A(n_421), .B(n_465), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_429), .B1(n_430), .B2(n_439), .C(n_440), .Y(n_422) );
OAI222xp33_ASAP7_75t_L g512 ( .A1(n_423), .A2(n_432), .B1(n_513), .B2(n_514), .C1(n_515), .C2(n_516), .Y(n_512) );
OAI21xp33_ASAP7_75t_SL g796 ( .A1(n_423), .A2(n_797), .B(n_798), .Y(n_796) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g1094 ( .A(n_424), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g546 ( .A(n_425), .Y(n_546) );
INVx4_ASAP7_75t_L g612 ( .A(n_425), .Y(n_612) );
BUFx3_ASAP7_75t_L g691 ( .A(n_425), .Y(n_691) );
INVx2_ASAP7_75t_L g887 ( .A(n_425), .Y(n_887) );
AND2x6_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g454 ( .A(n_426), .Y(n_454) );
AND2x4_ASAP7_75t_L g561 ( .A(n_426), .B(n_456), .Y(n_561) );
AND2x6_ASAP7_75t_L g476 ( .A(n_427), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g485 ( .A(n_427), .B(n_466), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_430), .A2(n_850), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_849) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g836 ( .A(n_433), .Y(n_836) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_434), .Y(n_600) );
BUFx4f_ASAP7_75t_SL g615 ( .A(n_434), .Y(n_615) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_434), .Y(n_664) );
BUFx2_ASAP7_75t_L g925 ( .A(n_434), .Y(n_925) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g444 ( .A(n_436), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_437), .Y(n_450) );
AND2x4_ASAP7_75t_L g443 ( .A(n_438), .B(n_444), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_438), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g558 ( .A(n_438), .B(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g515 ( .A(n_442), .Y(n_515) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx12f_ASAP7_75t_L g601 ( .A(n_443), .Y(n_601) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_443), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_451), .B2(n_452), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g618 ( .A1(n_447), .A2(n_452), .B1(n_619), .B2(n_620), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g827 ( .A1(n_447), .A2(n_828), .B1(n_829), .B2(n_830), .Y(n_827) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g930 ( .A(n_448), .Y(n_930) );
INVx4_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_449), .Y(n_519) );
BUFx3_ASAP7_75t_L g696 ( .A(n_449), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_449), .A2(n_452), .B1(n_800), .B2(n_801), .Y(n_799) );
AND2x2_ASAP7_75t_L g825 ( .A(n_450), .B(n_471), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_452), .A2(n_696), .B1(n_856), .B2(n_857), .Y(n_855) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_453), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_453), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_481), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_473), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx4f_ASAP7_75t_SL g711 ( .A(n_463), .Y(n_711) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g538 ( .A(n_464), .Y(n_538) );
BUFx3_ASAP7_75t_L g572 ( .A(n_464), .Y(n_572) );
BUFx3_ASAP7_75t_L g676 ( .A(n_464), .Y(n_676) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_465), .B(n_466), .Y(n_644) );
AND2x4_ASAP7_75t_L g470 ( .A(n_466), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
BUFx3_ASAP7_75t_L g591 ( .A(n_470), .Y(n_591) );
BUFx2_ASAP7_75t_L g678 ( .A(n_470), .Y(n_678) );
BUFx2_ASAP7_75t_SL g702 ( .A(n_470), .Y(n_702) );
BUFx2_ASAP7_75t_SL g805 ( .A(n_470), .Y(n_805) );
BUFx3_ASAP7_75t_L g881 ( .A(n_470), .Y(n_881) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x6_ASAP7_75t_L g496 ( .A(n_472), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx5_ASAP7_75t_SL g586 ( .A(n_475), .Y(n_586) );
INVx4_ASAP7_75t_L g635 ( .A(n_475), .Y(n_635) );
INVx2_ASAP7_75t_SL g730 ( .A(n_475), .Y(n_730) );
INVx1_ASAP7_75t_L g898 ( .A(n_475), .Y(n_898) );
INVx11_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx11_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g534 ( .A(n_479), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_479), .A2(n_633), .B1(n_634), .B2(n_636), .Y(n_632) );
INVx2_ASAP7_75t_L g671 ( .A(n_479), .Y(n_671) );
INVx2_ASAP7_75t_L g707 ( .A(n_479), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_479), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1012) );
INVx6_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g575 ( .A(n_480), .Y(n_575) );
BUFx3_ASAP7_75t_L g734 ( .A(n_480), .Y(n_734) );
BUFx3_ASAP7_75t_L g750 ( .A(n_480), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_489), .Y(n_481) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g526 ( .A(n_484), .Y(n_526) );
INVx3_ASAP7_75t_L g710 ( .A(n_484), .Y(n_710) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_484), .Y(n_812) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g565 ( .A(n_485), .Y(n_565) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_485), .Y(n_640) );
BUFx2_ASAP7_75t_SL g747 ( .A(n_485), .Y(n_747) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g528 ( .A(n_488), .Y(n_528) );
BUFx3_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_488), .Y(n_626) );
BUFx3_ASAP7_75t_L g883 ( .A(n_488), .Y(n_883) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g869 ( .A(n_491), .Y(n_869) );
INVx5_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g568 ( .A(n_492), .Y(n_568) );
INVx4_ASAP7_75t_L g630 ( .A(n_492), .Y(n_630) );
INVx3_ASAP7_75t_L g672 ( .A(n_492), .Y(n_672) );
BUFx3_ASAP7_75t_L g705 ( .A(n_492), .Y(n_705) );
INVx2_ASAP7_75t_L g935 ( .A(n_492), .Y(n_935) );
INVx8_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx4f_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
BUFx2_ASAP7_75t_L g631 ( .A(n_495), .Y(n_631) );
BUFx2_ASAP7_75t_L g752 ( .A(n_495), .Y(n_752) );
INVx6_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g674 ( .A(n_496), .Y(n_674) );
INVx1_ASAP7_75t_L g870 ( .A(n_496), .Y(n_870) );
INVx1_ASAP7_75t_SL g959 ( .A(n_496), .Y(n_959) );
INVx1_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_579), .B1(n_649), .B2(n_650), .Y(n_501) );
INVx1_ASAP7_75t_L g649 ( .A(n_502), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_542), .B1(n_577), .B2(n_578), .Y(n_502) );
INVx1_ASAP7_75t_L g577 ( .A(n_503), .Y(n_577) );
INVx1_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_523), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .C(n_517), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_510), .B2(n_511), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_508), .A2(n_828), .B1(n_920), .B2(n_921), .Y(n_919) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g686 ( .A(n_509), .Y(n_686) );
OA211x2_ASAP7_75t_L g592 ( .A1(n_511), .A2(n_593), .B(n_594), .C(n_596), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_511), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
BUFx3_ASAP7_75t_L g795 ( .A(n_511), .Y(n_795) );
INVx2_ASAP7_75t_L g848 ( .A(n_511), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_519), .A2(n_698), .B1(n_1136), .B2(n_1137), .Y(n_1135) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g698 ( .A(n_522), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_530), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g701 ( .A(n_528), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_535), .Y(n_530) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g574 ( .A(n_533), .Y(n_574) );
INVx4_ASAP7_75t_L g743 ( .A(n_533), .Y(n_743) );
INVx4_ASAP7_75t_L g823 ( .A(n_533), .Y(n_823) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx4_ASAP7_75t_SL g578 ( .A(n_542), .Y(n_578) );
AO22x2_ASAP7_75t_SL g604 ( .A1(n_542), .A2(n_578), .B1(n_605), .B2(n_647), .Y(n_604) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_576), .Y(n_542) );
NAND3x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_562), .C(n_570), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_546), .A2(n_666), .B(n_667), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_546), .A2(n_725), .B(n_726), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_546), .A2(n_764), .B(n_765), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g943 ( .A1(n_546), .A2(n_944), .B(n_945), .Y(n_943) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .C(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g979 ( .A(n_551), .Y(n_979) );
BUFx4f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g721 ( .A(n_552), .Y(n_721) );
BUFx2_ASAP7_75t_L g948 ( .A(n_552), .Y(n_948) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g595 ( .A(n_555), .Y(n_595) );
INVx5_ASAP7_75t_L g770 ( .A(n_555), .Y(n_770) );
INVx2_ASAP7_75t_L g907 ( .A(n_555), .Y(n_907) );
INVx4_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g597 ( .A(n_558), .Y(n_597) );
INVx1_ASAP7_75t_L g757 ( .A(n_558), .Y(n_757) );
BUFx2_ASAP7_75t_L g975 ( .A(n_558), .Y(n_975) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_561), .Y(n_598) );
BUFx2_ASAP7_75t_SL g668 ( .A(n_561), .Y(n_668) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_561), .Y(n_766) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
BUFx3_ASAP7_75t_L g1123 ( .A(n_572), .Y(n_1123) );
INVx1_ASAP7_75t_L g1014 ( .A(n_574), .Y(n_1014) );
INVx1_ASAP7_75t_L g650 ( .A(n_579), .Y(n_650) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AO22x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_603), .B1(n_604), .B2(n_648), .Y(n_580) );
INVx2_ASAP7_75t_SL g648 ( .A(n_581), .Y(n_648) );
XOR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_602), .Y(n_581) );
NAND4xp75_ASAP7_75t_L g582 ( .A(n_583), .B(n_588), .C(n_592), .D(n_599), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g810 ( .A(n_586), .Y(n_810) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_SL g951 ( .A(n_598), .Y(n_951) );
BUFx4f_ASAP7_75t_SL g854 ( .A(n_601), .Y(n_854) );
INVx2_ASAP7_75t_L g927 ( .A(n_601), .Y(n_927) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g647 ( .A(n_605), .Y(n_647) );
INVx1_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_621), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .C(n_618), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_613), .B(n_614), .Y(n_611) );
INVx4_ASAP7_75t_L g759 ( .A(n_612), .Y(n_759) );
OAI22xp5_ASAP7_75t_SL g834 ( .A1(n_612), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
BUFx2_ASAP7_75t_L g850 ( .A(n_612), .Y(n_850) );
OAI21xp5_ASAP7_75t_SL g1059 ( .A1(n_612), .A2(n_1060), .B(n_1061), .Y(n_1059) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g971 ( .A(n_617), .Y(n_971) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_632), .C(n_637), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx4_ASAP7_75t_L g1049 ( .A(n_625), .Y(n_1049) );
INVx4_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_630), .Y(n_1033) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_630), .Y(n_1051) );
INVx1_ASAP7_75t_L g990 ( .A(n_631), .Y(n_990) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_641), .B2(n_642), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_639), .A2(n_642), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_642), .A2(n_1017), .B1(n_1018), .B2(n_1019), .Y(n_1016) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g1072 ( .A(n_651), .Y(n_1072) );
XOR2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_914), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_784), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_714), .B1(n_782), .B2(n_783), .Y(n_653) );
INVx1_ASAP7_75t_L g782 ( .A(n_654), .Y(n_782) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_657), .B1(n_680), .B2(n_681), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
XOR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_679), .Y(n_657) );
NAND4xp75_ASAP7_75t_SL g658 ( .A(n_659), .B(n_669), .C(n_675), .D(n_677), .Y(n_658) );
NOR2xp67_ASAP7_75t_SL g659 ( .A(n_660), .B(n_665), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .C(n_663), .Y(n_660) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_664), .Y(n_693) );
INVx1_ASAP7_75t_L g1005 ( .A(n_664), .Y(n_1005) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
BUFx2_ASAP7_75t_L g982 ( .A(n_676), .Y(n_982) );
INVx1_ASAP7_75t_L g1031 ( .A(n_676), .Y(n_1031) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g712 ( .A(n_682), .Y(n_712) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_683), .B(n_699), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .C(n_694), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_686), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_686), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_844) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_692), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g922 ( .A1(n_690), .A2(n_923), .B(n_924), .Y(n_922) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g969 ( .A(n_693), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
AND4x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .C(n_706), .D(n_708), .Y(n_699) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g783 ( .A(n_714), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_737), .B1(n_738), .B2(n_781), .Y(n_714) );
INVx1_ASAP7_75t_SL g781 ( .A(n_715), .Y(n_781) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
XOR2x2_ASAP7_75t_SL g716 ( .A(n_717), .B(n_736), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g717 ( .A(n_718), .B(n_727), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_724), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .C(n_723), .Y(n_719) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_732), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g867 ( .A(n_730), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g863 ( .A(n_734), .Y(n_863) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AO22x1_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_760), .B1(n_779), .B2(n_780), .Y(n_738) );
INVx1_ASAP7_75t_L g779 ( .A(n_739), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .C(n_753), .D(n_758), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_751), .Y(n_745) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_SL g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g1130 ( .A(n_759), .Y(n_1130) );
INVx3_ASAP7_75t_SL g780 ( .A(n_760), .Y(n_780) );
XOR2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_778), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_762), .B(n_771), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_770), .Y(n_977) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_770), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_813), .B1(n_912), .B2(n_913), .Y(n_784) );
INVx1_ASAP7_75t_L g912 ( .A(n_785), .Y(n_912) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_802), .Y(n_790) );
NOR3xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_796), .C(n_799), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_807), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_811), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_810), .A2(n_863), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
INVx1_ASAP7_75t_SL g1018 ( .A(n_812), .Y(n_1018) );
INVx1_ASAP7_75t_L g913 ( .A(n_813), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_838), .B1(n_910), .B2(n_911), .Y(n_813) );
INVx1_ASAP7_75t_SL g910 ( .A(n_814), .Y(n_910) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NAND3x1_ASAP7_75t_SL g817 ( .A(n_818), .B(n_821), .C(n_826), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVx1_ASAP7_75t_L g994 ( .A(n_823), .Y(n_994) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .C(n_834), .Y(n_826) );
INVx1_ASAP7_75t_L g911 ( .A(n_838), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_872), .B2(n_873), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g871 ( .A(n_842), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_858), .Y(n_842) );
NOR3xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_849), .C(n_855), .Y(n_843) );
OAI211xp5_ASAP7_75t_L g999 ( .A1(n_847), .A2(n_1000), .B(n_1001), .C(n_1002), .Y(n_999) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NOR2xp67_ASAP7_75t_L g858 ( .A(n_859), .B(n_864), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B1(n_893), .B2(n_894), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
XOR2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_892), .Y(n_875) );
NAND4xp75_ASAP7_75t_SL g876 ( .A(n_877), .B(n_878), .C(n_879), .D(n_884), .Y(n_876) );
AND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_883), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_889), .Y(n_884) );
OAI21xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B(n_888), .Y(n_885) );
OAI222xp33_ASAP7_75t_L g967 ( .A1(n_887), .A2(n_968), .B1(n_969), .B2(n_970), .C1(n_971), .C2(n_972), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NAND4xp75_ASAP7_75t_L g895 ( .A(n_896), .B(n_900), .C(n_903), .D(n_909), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .Y(n_896) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
OA211x2_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B(n_906), .C(n_908), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_962), .B1(n_1070), .B2(n_1071), .Y(n_914) );
INVx2_ASAP7_75t_L g1070 ( .A(n_915), .Y(n_1070) );
XNOR2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_940), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g1042 ( .A(n_916), .B(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_SL g938 ( .A(n_917), .Y(n_938) );
AND2x2_ASAP7_75t_SL g917 ( .A(n_918), .B(n_932), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_922), .C(n_928), .Y(n_918) );
INVx1_ASAP7_75t_L g1132 ( .A(n_925), .Y(n_1132) );
INVx1_ASAP7_75t_L g1007 ( .A(n_926), .Y(n_1007) );
INVx3_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
AND4x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .C(n_936), .D(n_937), .Y(n_932) );
INVx2_ASAP7_75t_SL g960 ( .A(n_941), .Y(n_960) );
AND2x2_ASAP7_75t_L g941 ( .A(n_942), .B(n_952), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .Y(n_942) );
NAND2xp5_ASAP7_75t_SL g946 ( .A(n_947), .B(n_949), .Y(n_946) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_953), .B(n_956), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .Y(n_956) );
INVx1_ASAP7_75t_SL g1071 ( .A(n_962), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_1022), .B1(n_1023), .B2(n_1069), .Y(n_962) );
INVx1_ASAP7_75t_L g1069 ( .A(n_963), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_995), .B1(n_1020), .B2(n_1021), .Y(n_963) );
INVx1_ASAP7_75t_L g1021 ( .A(n_964), .Y(n_1021) );
NAND3x1_ASAP7_75t_L g965 ( .A(n_966), .B(n_980), .C(n_985), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_973), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_976), .Y(n_973) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
AND2x2_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .Y(n_980) );
OAI22xp5_ASAP7_75t_SL g986 ( .A1(n_987), .A2(n_989), .B1(n_990), .B2(n_991), .Y(n_986) );
BUFx2_ASAP7_75t_R g987 ( .A(n_988), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g1020 ( .A(n_995), .Y(n_1020) );
XNOR2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
AND2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1008), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1006), .B2(n_1007), .Y(n_1003) );
NOR3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .C(n_1016), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
INVx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
AO22x1_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1042), .B2(n_1068), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_SL g1041 ( .A(n_1027), .Y(n_1041) );
NAND4xp75_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1034), .C(n_1037), .D(n_1040), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1032), .Y(n_1028) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
AND2x2_ASAP7_75t_SL g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1042), .Y(n_1068) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AND2x2_ASAP7_75t_SL g1045 ( .A(n_1046), .B(n_1058), .Y(n_1045) );
NOR3xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1052), .C(n_1055), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1050), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1062), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .C(n_1066), .Y(n_1062) );
INVx1_ASAP7_75t_SL g1074 ( .A(n_1075), .Y(n_1074) );
NOR2x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1080), .Y(n_1075) );
OR2x2_ASAP7_75t_SL g1141 ( .A(n_1076), .B(n_1081), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1079), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_1077), .Y(n_1107) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1078), .B(n_1110), .Y(n_1113) );
CKINVDCx16_ASAP7_75t_R g1110 ( .A(n_1079), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_1081), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
OAI322xp33_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1106), .A3(n_1108), .B1(n_1111), .B2(n_1114), .C1(n_1115), .C2(n_1139), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_1090), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
NAND4xp75_ASAP7_75t_SL g1091 ( .A(n_1092), .B(n_1101), .C(n_1104), .D(n_1105), .Y(n_1091) );
NOR2xp67_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1097), .Y(n_1092) );
OAI21xp5_ASAP7_75t_SL g1093 ( .A1(n_1094), .A2(n_1095), .B(n_1096), .Y(n_1093) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .C(n_1100), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1103), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
CKINVDCx16_ASAP7_75t_R g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1116), .Y(n_1138) );
AND2x2_ASAP7_75t_SL g1116 ( .A(n_1117), .B(n_1125), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1121), .Y(n_1117) );
NAND2xp33_ASAP7_75t_SL g1118 ( .A(n_1119), .B(n_1120), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1124), .Y(n_1121) );
NOR3xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1129), .C(n_1135), .Y(n_1125) );
OAI221xp5_ASAP7_75t_SL g1129 ( .A1(n_1130), .A2(n_1131), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_1129) );
CKINVDCx20_ASAP7_75t_R g1139 ( .A(n_1140), .Y(n_1139) );
CKINVDCx20_ASAP7_75t_R g1140 ( .A(n_1141), .Y(n_1140) );
endmodule