module fake_jpeg_11076_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_3),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_16),
.C(n_19),
.Y(n_20)
);

NOR2x1_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_17),
.B(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_5),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_5),
.B2(n_8),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_6),
.Y(n_18)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_11),
.C(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_15),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_15),
.B1(n_18),
.B2(n_9),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_20),
.B(n_19),
.C(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_14),
.C(n_23),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_13),
.Y(n_31)
);


endmodule