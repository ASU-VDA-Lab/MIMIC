module real_aes_7937_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_706, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_706;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_169), .C(n_173), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_1), .B(n_162), .Y(n_175) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_3), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_4), .A2(n_136), .B(n_153), .C(n_459), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_5), .A2(n_156), .B(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_6), .A2(n_156), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_7), .B(n_162), .Y(n_486) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_128), .B(n_215), .Y(n_214) );
AND2x6_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_10), .A2(n_136), .B(n_153), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g451 ( .A(n_11), .Y(n_451) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_12), .B(n_41), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_13), .B(n_172), .Y(n_461) );
INVx1_ASAP7_75t_L g133 ( .A(n_14), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_15), .B(n_147), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_16), .A2(n_148), .B(n_470), .C(n_472), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_17), .B(n_162), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_18), .A2(n_65), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_18), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_19), .B(n_205), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_20), .A2(n_136), .B(n_199), .C(n_204), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_21), .A2(n_171), .B(n_223), .C(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_22), .B(n_172), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_23), .B(n_172), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_24), .Y(n_489) );
INVx1_ASAP7_75t_L g501 ( .A(n_25), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_26), .A2(n_136), .B(n_204), .C(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_28), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_29), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g518 ( .A(n_30), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_31), .A2(n_156), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_33), .A2(n_151), .B(n_183), .C(n_184), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_34), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_35), .A2(n_171), .B(n_483), .C(n_485), .Y(n_482) );
INVxp67_ASAP7_75t_L g519 ( .A(n_36), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_37), .B(n_220), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g481 ( .A(n_38), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_39), .A2(n_136), .B(n_204), .C(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_40), .A2(n_102), .B1(n_111), .B2(n_704), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_41), .B(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_42), .A2(n_173), .B(n_449), .C(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_43), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_44), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_45), .B(n_147), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_46), .B(n_156), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_47), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_48), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_49), .A2(n_151), .B(n_183), .C(n_244), .Y(n_243) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_50), .A2(n_422), .B1(n_691), .B2(n_692), .C1(n_695), .C2(n_698), .Y(n_421) );
INVx1_ASAP7_75t_L g170 ( .A(n_51), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_52), .A2(n_82), .B1(n_693), .B2(n_694), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_52), .Y(n_694) );
INVx1_ASAP7_75t_L g245 ( .A(n_53), .Y(n_245) );
INVx1_ASAP7_75t_L g439 ( .A(n_54), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_55), .B(n_156), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_56), .Y(n_208) );
CKINVDCx14_ASAP7_75t_R g447 ( .A(n_57), .Y(n_447) );
INVx1_ASAP7_75t_L g154 ( .A(n_58), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_59), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_60), .B(n_162), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_61), .A2(n_143), .B(n_203), .C(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
INVx1_ASAP7_75t_SL g484 ( .A(n_63), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_66), .B(n_147), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_67), .B(n_162), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_68), .B(n_148), .Y(n_234) );
INVx1_ASAP7_75t_L g492 ( .A(n_69), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_70), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_71), .B(n_187), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_72), .A2(n_136), .B(n_141), .C(n_151), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_73), .Y(n_259) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_75), .A2(n_156), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_76), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_77), .A2(n_156), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_78), .A2(n_197), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g468 ( .A(n_79), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_80), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_81), .B(n_186), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_82), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_83), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_84), .A2(n_156), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g471 ( .A(n_85), .Y(n_471) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx1_ASAP7_75t_L g460 ( .A(n_87), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_88), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_89), .B(n_172), .Y(n_235) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_90), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g414 ( .A(n_90), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g425 ( .A(n_90), .B(n_416), .Y(n_425) );
INVx2_ASAP7_75t_L g429 ( .A(n_90), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_91), .A2(n_136), .B(n_151), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_92), .B(n_156), .Y(n_181) );
INVx1_ASAP7_75t_L g185 ( .A(n_93), .Y(n_185) );
INVxp67_ASAP7_75t_L g262 ( .A(n_94), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_95), .B(n_128), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
INVx1_ASAP7_75t_L g230 ( .A(n_98), .Y(n_230) );
INVx2_ASAP7_75t_L g442 ( .A(n_99), .Y(n_442) );
AND2x2_ASAP7_75t_L g247 ( .A(n_100), .B(n_190), .Y(n_247) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g704 ( .A(n_103), .Y(n_704) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g416 ( .A(n_107), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_420), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g703 ( .A(n_115), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_412), .B(n_418), .Y(n_116) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx2_ASAP7_75t_L g426 ( .A(n_121), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_121), .A2(n_424), .B1(n_700), .B2(n_701), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_355), .Y(n_121) );
AND4x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_295), .C(n_310), .D(n_335), .Y(n_122) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_268), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_176), .B(n_248), .Y(n_124) );
AND2x2_ASAP7_75t_L g298 ( .A(n_125), .B(n_194), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_125), .B(n_193), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_125), .B(n_177), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_125), .Y(n_365) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
INVx2_ASAP7_75t_L g282 ( .A(n_126), .Y(n_282) );
BUFx2_ASAP7_75t_L g309 ( .A(n_126), .Y(n_309) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_159), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_127), .B(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_127), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_127), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_127), .A2(n_229), .B(n_236), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_127), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_127), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_127), .B(n_504), .Y(n_503) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_128), .A2(n_216), .B(n_217), .Y(n_215) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_128), .Y(n_256) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g238 ( .A(n_129), .Y(n_238) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_130), .B(n_131), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_155), .Y(n_134) );
INVx5_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx3_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g224 ( .A(n_138), .Y(n_224) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
AND2x2_ASAP7_75t_L g157 ( .A(n_140), .B(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_144), .B(n_442), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_144), .B(n_471), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_144), .A2(n_147), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx2_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_147), .B(n_262), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_147), .A2(n_202), .B(n_501), .C(n_502), .Y(n_500) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_148), .B(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g485 ( .A(n_150), .Y(n_485) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_152), .A2(n_165), .B(n_166), .C(n_167), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_152), .A2(n_166), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g438 ( .A1(n_152), .A2(n_166), .B(n_439), .C(n_440), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_152), .A2(n_166), .B(n_447), .C(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_152), .A2(n_166), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_152), .A2(n_166), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_152), .A2(n_166), .B(n_515), .C(n_516), .Y(n_514) );
INVx4_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g156 ( .A(n_153), .B(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_153), .B(n_157), .Y(n_231) );
BUFx2_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx1_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
AND2x2_ASAP7_75t_L g249 ( .A(n_161), .B(n_194), .Y(n_249) );
INVx2_ASAP7_75t_L g265 ( .A(n_161), .Y(n_265) );
AND2x2_ASAP7_75t_L g274 ( .A(n_161), .B(n_193), .Y(n_274) );
AND2x2_ASAP7_75t_L g353 ( .A(n_161), .B(n_282), .Y(n_353) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_175), .Y(n_161) );
INVx2_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_171), .B(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g449 ( .A(n_172), .Y(n_449) );
INVx2_ASAP7_75t_L g462 ( .A(n_173), .Y(n_462) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
INVx1_ASAP7_75t_L g472 ( .A(n_174), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_210), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_177), .B(n_280), .Y(n_318) );
INVx1_ASAP7_75t_L g406 ( .A(n_177), .Y(n_406) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
AND2x2_ASAP7_75t_L g264 ( .A(n_178), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g278 ( .A(n_178), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_178), .Y(n_307) );
OR2x2_ASAP7_75t_L g339 ( .A(n_178), .B(n_281), .Y(n_339) );
AND2x2_ASAP7_75t_L g347 ( .A(n_178), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g380 ( .A(n_178), .B(n_349), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_178), .B(n_249), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_178), .B(n_309), .Y(n_405) );
AND2x2_ASAP7_75t_L g411 ( .A(n_178), .B(n_298), .Y(n_411) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g271 ( .A(n_179), .Y(n_271) );
AND2x2_ASAP7_75t_L g301 ( .A(n_179), .B(n_281), .Y(n_301) );
AND2x2_ASAP7_75t_L g334 ( .A(n_179), .B(n_294), .Y(n_334) );
AND2x2_ASAP7_75t_L g354 ( .A(n_179), .B(n_194), .Y(n_354) );
AND2x2_ASAP7_75t_L g388 ( .A(n_179), .B(n_254), .Y(n_388) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_191), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_190), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_186), .A2(n_189), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g459 ( .A1(n_186), .A2(n_460), .B(n_461), .C(n_462), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_186), .A2(n_462), .B(n_492), .C(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
INVx1_ASAP7_75t_L g209 ( .A(n_190), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_190), .A2(n_242), .B(n_243), .Y(n_241) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_190), .A2(n_445), .B(n_452), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_190), .A2(n_231), .B(n_498), .C(n_499), .Y(n_497) );
AND2x4_ASAP7_75t_L g294 ( .A(n_193), .B(n_265), .Y(n_294) );
AND2x2_ASAP7_75t_L g305 ( .A(n_193), .B(n_301), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_193), .B(n_281), .Y(n_344) );
INVx2_ASAP7_75t_L g359 ( .A(n_193), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_193), .B(n_293), .Y(n_382) );
AND2x2_ASAP7_75t_L g401 ( .A(n_193), .B(n_353), .Y(n_401) );
INVx5_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
AND2x2_ASAP7_75t_L g308 ( .A(n_194), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g349 ( .A(n_194), .B(n_265), .Y(n_349) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
AOI21xp5_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_198), .B(n_205), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .Y(n_199) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_203), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_206), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_209), .A2(n_456), .B(n_463), .Y(n_455) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
AND2x2_ASAP7_75t_L g272 ( .A(n_212), .B(n_255), .Y(n_272) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_213), .B(n_228), .Y(n_252) );
OR2x2_ASAP7_75t_L g285 ( .A(n_213), .B(n_255), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_213), .B(n_255), .Y(n_290) );
AND2x2_ASAP7_75t_L g317 ( .A(n_213), .B(n_254), .Y(n_317) );
AND2x2_ASAP7_75t_L g369 ( .A(n_213), .B(n_227), .Y(n_369) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_214), .B(n_239), .Y(n_277) );
AND2x2_ASAP7_75t_L g313 ( .A(n_214), .B(n_228), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_221), .B(n_222), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_222), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_225), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g303 ( .A(n_226), .B(n_285), .Y(n_303) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_239), .Y(n_226) );
OAI322xp33_ASAP7_75t_L g268 ( .A1(n_227), .A2(n_269), .A3(n_273), .B1(n_275), .B2(n_278), .C1(n_283), .C2(n_291), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_227), .B(n_254), .Y(n_276) );
OR2x2_ASAP7_75t_L g286 ( .A(n_227), .B(n_240), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_227), .B(n_240), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_227), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_227), .B(n_255), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_227), .B(n_384), .Y(n_383) );
INVx5_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_228), .B(n_272), .Y(n_398) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_231), .A2(n_457), .B(n_458), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_231), .A2(n_489), .B(n_490), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g512 ( .A(n_238), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_239), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_239), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g328 ( .A(n_239), .B(n_255), .Y(n_328) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_239), .A2(n_357), .B(n_360), .C(n_372), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_239), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g394 ( .A(n_239), .B(n_369), .Y(n_394) );
INVx5_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g322 ( .A(n_240), .B(n_255), .Y(n_322) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_240), .Y(n_331) );
AND2x2_ASAP7_75t_L g371 ( .A(n_240), .B(n_369), .Y(n_371) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_240), .B(n_272), .Y(n_402) );
AND2x2_ASAP7_75t_L g409 ( .A(n_240), .B(n_368), .Y(n_409) );
OR2x6_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B1(n_264), .B2(n_266), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_249), .B(n_271), .Y(n_319) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g267 ( .A(n_252), .Y(n_267) );
OR2x2_ASAP7_75t_L g327 ( .A(n_252), .B(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g375 ( .A1(n_252), .A2(n_376), .B1(n_378), .B2(n_379), .C(n_381), .Y(n_375) );
INVx2_ASAP7_75t_L g314 ( .A(n_253), .Y(n_314) );
AND2x2_ASAP7_75t_L g287 ( .A(n_254), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g377 ( .A(n_254), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_254), .B(n_369), .Y(n_390) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVxp67_ASAP7_75t_L g332 ( .A(n_255), .Y(n_332) );
AND2x2_ASAP7_75t_L g368 ( .A(n_255), .B(n_369), .Y(n_368) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_263), .Y(n_255) );
OA21x2_ASAP7_75t_L g436 ( .A1(n_256), .A2(n_437), .B(n_443), .Y(n_436) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_256), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_256), .A2(n_479), .B(n_486), .Y(n_478) );
AND2x2_ASAP7_75t_L g370 ( .A(n_264), .B(n_309), .Y(n_370) );
AND2x2_ASAP7_75t_L g280 ( .A(n_265), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_265), .B(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_267), .B(n_314), .Y(n_351) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g357 ( .A(n_270), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OR2x2_ASAP7_75t_L g343 ( .A(n_271), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g408 ( .A(n_271), .B(n_353), .Y(n_408) );
INVx2_ASAP7_75t_L g341 ( .A(n_272), .Y(n_341) );
NAND4xp25_ASAP7_75t_SL g404 ( .A(n_273), .B(n_405), .C(n_406), .D(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_274), .B(n_338), .Y(n_373) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_SL g410 ( .A(n_277), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_SL g372 ( .A1(n_278), .A2(n_341), .B(n_345), .C(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g367 ( .A(n_280), .B(n_359), .Y(n_367) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_281), .Y(n_293) );
INVx1_ASAP7_75t_L g348 ( .A(n_281), .Y(n_348) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
AOI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B(n_287), .C(n_289), .Y(n_283) );
AND2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_288), .Y(n_304) );
OAI322xp33_ASAP7_75t_SL g342 ( .A1(n_284), .A2(n_343), .A3(n_345), .B1(n_346), .B2(n_350), .C1(n_351), .C2(n_352), .Y(n_342) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g364 ( .A(n_286), .B(n_290), .Y(n_364) );
INVx1_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
INVx1_ASAP7_75t_SL g363 ( .A(n_290), .Y(n_363) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AOI222xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_302), .B1(n_304), .B2(n_305), .C1(n_306), .C2(n_706), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_297), .A2(n_359), .A3(n_364), .B1(n_386), .B2(n_387), .C1(n_389), .C2(n_390), .Y(n_385) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_298), .A2(n_312), .B1(n_336), .B2(n_340), .C(n_342), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI222xp33_ASAP7_75t_L g315 ( .A1(n_303), .A2(n_316), .B1(n_318), .B2(n_319), .C1(n_320), .C2(n_323), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_305), .A2(n_312), .B1(n_382), .B2(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_315), .C(n_326), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_312), .A2(n_349), .B(n_392), .C(n_395), .Y(n_391) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_313), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g384 ( .A(n_317), .Y(n_384) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_324), .B(n_349), .Y(n_378) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B(n_333), .Y(n_326) );
OAI221xp5_ASAP7_75t_SL g395 ( .A1(n_327), .A2(n_396), .B1(n_397), .B2(n_398), .C(n_399), .Y(n_395) );
INVxp33_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_331), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_338), .B(n_349), .Y(n_389) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g400 ( .A(n_353), .B(n_359), .Y(n_400) );
AND4x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_374), .C(n_391), .D(n_403), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B1(n_364), .B2(n_365), .C(n_366), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_370), .B2(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
INVx1_ASAP7_75t_SL g386 ( .A(n_371), .Y(n_386) );
NOR2xp33_ASAP7_75t_SL g374 ( .A(n_375), .B(n_385), .Y(n_374) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_387), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_394), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_409), .B1(n_410), .B2(n_411), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g419 ( .A(n_414), .Y(n_419) );
NOR2x2_ASAP7_75t_L g697 ( .A(n_415), .B(n_429), .Y(n_697) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g428 ( .A(n_416), .B(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_418), .A2(n_421), .B(n_702), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx6_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g700 ( .A(n_428), .Y(n_700) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g701 ( .A(n_431), .Y(n_701) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_617), .Y(n_431) );
NOR4xp25_ASAP7_75t_L g432 ( .A(n_433), .B(n_559), .C(n_589), .D(n_599), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_474), .B(n_522), .C(n_549), .Y(n_433) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_434), .A2(n_564), .B1(n_645), .B2(n_646), .C1(n_647), .C2(n_648), .Y(n_644) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_453), .Y(n_434) );
AOI33xp33_ASAP7_75t_L g570 ( .A1(n_435), .A2(n_557), .A3(n_558), .B1(n_571), .B2(n_576), .B3(n_578), .Y(n_570) );
OAI211xp5_ASAP7_75t_SL g627 ( .A1(n_435), .A2(n_628), .B(n_630), .C(n_632), .Y(n_627) );
OR2x2_ASAP7_75t_L g643 ( .A(n_435), .B(n_629), .Y(n_643) );
INVx1_ASAP7_75t_L g676 ( .A(n_435), .Y(n_676) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_444), .Y(n_435) );
INVx2_ASAP7_75t_L g553 ( .A(n_436), .Y(n_553) );
AND2x2_ASAP7_75t_L g569 ( .A(n_436), .B(n_465), .Y(n_569) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_436), .Y(n_604) );
AND2x2_ASAP7_75t_L g633 ( .A(n_436), .B(n_444), .Y(n_633) );
INVx2_ASAP7_75t_L g533 ( .A(n_444), .Y(n_533) );
BUFx3_ASAP7_75t_L g541 ( .A(n_444), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_444), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g552 ( .A(n_444), .B(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_444), .B(n_454), .Y(n_581) );
AND2x2_ASAP7_75t_L g650 ( .A(n_444), .B(n_584), .Y(n_650) );
INVx2_ASAP7_75t_SL g544 ( .A(n_453), .Y(n_544) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_465), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_454), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g586 ( .A(n_454), .Y(n_586) );
AND2x2_ASAP7_75t_L g597 ( .A(n_454), .B(n_553), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_454), .B(n_582), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_454), .B(n_584), .Y(n_629) );
AND2x2_ASAP7_75t_L g688 ( .A(n_454), .B(n_633), .Y(n_688) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g558 ( .A(n_455), .B(n_465), .Y(n_558) );
AND2x2_ASAP7_75t_L g568 ( .A(n_455), .B(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g590 ( .A(n_455), .Y(n_590) );
AND3x2_ASAP7_75t_L g649 ( .A(n_455), .B(n_650), .C(n_651), .Y(n_649) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_465), .Y(n_540) );
INVx1_ASAP7_75t_SL g584 ( .A(n_465), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_465), .B(n_533), .C(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_505), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_475), .A2(n_568), .B(n_620), .C(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_477), .B(n_496), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_477), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_SL g636 ( .A(n_477), .Y(n_636) );
AND2x2_ASAP7_75t_L g657 ( .A(n_477), .B(n_507), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_477), .B(n_566), .Y(n_685) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
AND2x2_ASAP7_75t_L g530 ( .A(n_478), .B(n_521), .Y(n_530) );
INVx2_ASAP7_75t_L g537 ( .A(n_478), .Y(n_537) );
AND2x2_ASAP7_75t_L g557 ( .A(n_478), .B(n_507), .Y(n_557) );
AND2x2_ASAP7_75t_L g607 ( .A(n_478), .B(n_496), .Y(n_607) );
INVx1_ASAP7_75t_L g611 ( .A(n_478), .Y(n_611) );
INVx2_ASAP7_75t_SL g521 ( .A(n_487), .Y(n_521) );
BUFx2_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
AND2x2_ASAP7_75t_L g674 ( .A(n_487), .B(n_496), .Y(n_674) );
INVx3_ASAP7_75t_SL g507 ( .A(n_496), .Y(n_507) );
AND2x2_ASAP7_75t_L g529 ( .A(n_496), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g536 ( .A(n_496), .B(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g566 ( .A(n_496), .B(n_526), .Y(n_566) );
OR2x2_ASAP7_75t_L g575 ( .A(n_496), .B(n_521), .Y(n_575) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_496), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_496), .B(n_551), .Y(n_598) );
AND2x2_ASAP7_75t_L g626 ( .A(n_496), .B(n_509), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_496), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g664 ( .A(n_496), .B(n_508), .Y(n_664) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g588 ( .A(n_507), .B(n_537), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_507), .B(n_530), .Y(n_616) );
AND2x2_ASAP7_75t_L g634 ( .A(n_507), .B(n_551), .Y(n_634) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
AND2x2_ASAP7_75t_L g535 ( .A(n_509), .B(n_521), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_509), .B(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
OR2x2_ASAP7_75t_L g621 ( .A(n_509), .B(n_541), .Y(n_621) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_513), .B(n_520), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_511), .A2(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g527 ( .A(n_513), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_520), .Y(n_528) );
AND2x2_ASAP7_75t_L g556 ( .A(n_521), .B(n_526), .Y(n_556) );
INVx1_ASAP7_75t_L g564 ( .A(n_521), .Y(n_564) );
AND2x2_ASAP7_75t_L g659 ( .A(n_521), .B(n_537), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_531), .B1(n_534), .B2(n_538), .C1(n_542), .C2(n_545), .Y(n_522) );
INVx1_ASAP7_75t_L g654 ( .A(n_523), .Y(n_654) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
AND2x2_ASAP7_75t_L g550 ( .A(n_524), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g561 ( .A(n_524), .B(n_530), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_524), .B(n_552), .Y(n_577) );
OAI222xp33_ASAP7_75t_L g599 ( .A1(n_524), .A2(n_600), .B1(n_605), .B2(n_606), .C1(n_614), .C2(n_616), .Y(n_599) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g587 ( .A(n_526), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_526), .B(n_607), .Y(n_647) );
AND2x2_ASAP7_75t_L g658 ( .A(n_526), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g666 ( .A(n_529), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_531), .B(n_582), .Y(n_645) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_533), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_533), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx3_ASAP7_75t_L g548 ( .A(n_536), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_536), .A2(n_639), .B(n_642), .C(n_644), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_536), .B(n_573), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_536), .B(n_556), .Y(n_678) );
AND2x2_ASAP7_75t_L g551 ( .A(n_537), .B(n_547), .Y(n_551) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_541), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g630 ( .A(n_541), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g669 ( .A(n_541), .B(n_569), .Y(n_669) );
INVx1_ASAP7_75t_L g681 ( .A(n_541), .Y(n_681) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_544), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g662 ( .A(n_547), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_552), .B(n_554), .C(n_558), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_550), .A2(n_580), .B1(n_595), .B2(n_598), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_551), .B(n_565), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_551), .B(n_573), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_552), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g615 ( .A(n_552), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_552), .B(n_602), .Y(n_622) );
INVx2_ASAP7_75t_L g583 ( .A(n_553), .Y(n_583) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NOR4xp25_ASAP7_75t_L g560 ( .A(n_557), .B(n_561), .C(n_562), .D(n_565), .Y(n_560) );
INVx1_ASAP7_75t_SL g631 ( .A(n_558), .Y(n_631) );
AND2x2_ASAP7_75t_L g675 ( .A(n_558), .B(n_676), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_567), .B(n_570), .C(n_579), .Y(n_559) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_566), .B(n_636), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_568), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_SL g641 ( .A(n_569), .Y(n_641) );
AND2x2_ASAP7_75t_L g680 ( .A(n_569), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_573), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_577), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_578), .B(n_603), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_585), .B(n_587), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g655 ( .A(n_582), .Y(n_655) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g683 ( .A(n_583), .Y(n_683) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_584), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_594), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_590), .Y(n_602) );
OR2x2_ASAP7_75t_L g640 ( .A(n_590), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI21xp33_ASAP7_75t_SL g635 ( .A1(n_593), .A2(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_597), .A2(n_624), .B1(n_627), .B2(n_634), .C(n_635), .Y(n_623) );
INVx1_ASAP7_75t_SL g667 ( .A(n_598), .Y(n_667) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OR2x2_ASAP7_75t_L g614 ( .A(n_602), .B(n_615), .Y(n_614) );
INVxp67_ASAP7_75t_L g651 ( .A(n_604), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_611), .B2(n_612), .Y(n_606) );
INVx1_ASAP7_75t_L g646 ( .A(n_607), .Y(n_646) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_610), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR4xp25_ASAP7_75t_L g617 ( .A(n_618), .B(n_652), .C(n_665), .D(n_677), .Y(n_617) );
NAND3xp33_ASAP7_75t_SL g618 ( .A(n_619), .B(n_623), .C(n_638), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_621), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_628), .B(n_633), .Y(n_637) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_640), .A2(n_666), .B1(n_667), .B2(n_668), .C(n_670), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_642), .A2(n_657), .B(n_658), .C(n_660), .Y(n_656) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_643), .A2(n_661), .B1(n_663), .B2(n_664), .Y(n_660) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_655), .C(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g671 ( .A(n_664), .Y(n_671) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_672), .B(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx3_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
endmodule