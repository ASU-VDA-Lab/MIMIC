module fake_jpeg_11146_n_298 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_45),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_59),
.Y(n_71)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_2),
.C(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_66),
.B(n_70),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_25),
.B1(n_30),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_99),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_43),
.B(n_39),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_74),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_33),
.B1(n_42),
.B2(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_30),
.B1(n_25),
.B2(n_43),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_30),
.B1(n_25),
.B2(n_39),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_36),
.B1(n_35),
.B2(n_24),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_104),
.A3(n_67),
.B1(n_54),
.B2(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_38),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_36),
.B1(n_35),
.B2(n_38),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_37),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_44),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_109),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_37),
.B1(n_34),
.B2(n_27),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_64),
.B(n_34),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_21),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_85),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_91),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_129),
.Y(n_167)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_138),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_45),
.B1(n_27),
.B2(n_21),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_149),
.B1(n_122),
.B2(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_56),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_133),
.Y(n_165)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_81),
.B(n_67),
.CON(n_131),
.SN(n_131)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_97),
.Y(n_170)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_4),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_147),
.Y(n_151)
);

OR2x2_ASAP7_75t_SL g137 ( 
.A(n_86),
.B(n_5),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_13),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_14),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_6),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_8),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_82),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_90),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_90),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_166),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_75),
.B1(n_88),
.B2(n_87),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_116),
.B1(n_148),
.B2(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_89),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_178),
.Y(n_199)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_172),
.B(n_136),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_10),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_173),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_83),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_97),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_117),
.B(n_83),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_114),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_105),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_91),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_137),
.A3(n_140),
.B1(n_123),
.B2(n_116),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_105),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_121),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_140),
.C(n_136),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_158),
.C(n_165),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_191),
.B(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_146),
.B(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_209),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_156),
.B1(n_181),
.B2(n_163),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_200),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_167),
.B1(n_151),
.B2(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_202),
.B1(n_205),
.B2(n_207),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_121),
.B1(n_139),
.B2(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_206),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_170),
.B1(n_162),
.B2(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_164),
.B1(n_159),
.B2(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_217),
.C(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_221),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_228),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_153),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_223),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_163),
.B(n_197),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_199),
.B1(n_184),
.B2(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_187),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_199),
.B1(n_192),
.B2(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_218),
.B(n_210),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_182),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_183),
.C(n_189),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_216),
.C(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_200),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_222),
.B1(n_214),
.B2(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_247),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_258),
.C(n_238),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_254),
.B(n_255),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_226),
.B1(n_210),
.B2(n_214),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_246),
.B1(n_235),
.B2(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_220),
.C(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_249),
.C(n_259),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_240),
.B1(n_244),
.B2(n_239),
.C(n_235),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_258),
.B1(n_261),
.B2(n_202),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_234),
.C(n_209),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_259),
.C(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_272),
.C(n_264),
.Y(n_282)
);

AOI211xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_261),
.B(n_255),
.C(n_233),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_219),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_232),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_278),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_274),
.B(n_279),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_282),
.B(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.C(n_289),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_275),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_294),
.B(n_243),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_201),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_203),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_297),
.Y(n_298)
);


endmodule