module fake_jpeg_21327_n_86 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_8),
.B1(n_10),
.B2(n_15),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_13),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_18),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_21),
.C(n_26),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_43),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_42),
.B(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_51),
.B1(n_41),
.B2(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_47),
.B1(n_33),
.B2(n_8),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_40),
.C(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.C(n_27),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_42),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_11),
.B(n_15),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_9),
.B(n_12),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_55),
.B(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_9),
.B1(n_36),
.B2(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_58),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_73),
.B(n_59),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_77),
.B1(n_16),
.B2(n_4),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_16),
.B(n_4),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_69),
.C(n_61),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_2),
.B(n_5),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.C(n_76),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_16),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_6),
.Y(n_86)
);


endmodule