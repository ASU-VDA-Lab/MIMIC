module real_jpeg_999_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_2),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_31),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_3),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_3),
.B(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_5),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_10),
.B(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_12),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_12),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_12),
.B(n_23),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_12),
.B(n_28),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_85),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_84),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_54),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_18),
.B(n_54),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.C(n_46),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_30),
.C(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_66),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_28),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_37),
.A2(n_38),
.B1(n_46),
.B2(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.C(n_42),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_39),
.B(n_41),
.CI(n_42),
.CON(n_91),
.SN(n_91)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_49),
.C(n_50),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_72),
.B2(n_73),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_56),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_64),
.CI(n_71),
.CON(n_56),
.SN(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_99),
.B(n_129),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_90),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.C(n_98),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_126),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_91),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_123),
.B(n_128),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_112),
.B(n_122),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_105),
.C(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B(n_121),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);


endmodule