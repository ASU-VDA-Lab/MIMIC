module fake_jpeg_11785_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_16),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_10),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_12),
.B1(n_15),
.B2(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_12),
.B1(n_29),
.B2(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_32),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_56),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_41),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_58),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_60),
.B(n_59),
.C(n_51),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_53),
.B(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_26),
.C(n_4),
.Y(n_67)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_67),
.B(n_4),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_1),
.B(n_6),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_46),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_47),
.B(n_42),
.Y(n_72)
);


endmodule