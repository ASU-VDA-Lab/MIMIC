module real_jpeg_31365_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

NAND2xp67_ASAP7_75t_SL g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_1),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_1),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_1),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_1),
.B(n_372),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_4),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_5),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_6),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_6),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_57),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g71 ( 
.A(n_7),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_7),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_121),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_7),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_8),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_8),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_8),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_8),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_8),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_9),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_9),
.B(n_326),
.Y(n_325)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_9),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_10),
.B(n_77),
.Y(n_76)
);

NAND2x2_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_10),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_10),
.B(n_132),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_13),
.B(n_61),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_13),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_13),
.B(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_16),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_16),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_16),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_17),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_17),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_17),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_17),
.B(n_352),
.Y(n_351)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_75),
.B(n_283),
.C(n_436),
.D(n_445),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_248),
.C(n_273),
.Y(n_24)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_199),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_27),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_162),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_28),
.B(n_162),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_98),
.C(n_134),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_29),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_67),
.C(n_81),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_31),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_45),
.C(n_54),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_32),
.B(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_34),
.A2(n_35),
.B1(n_239),
.B2(n_260),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_34),
.B(n_159),
.C(n_239),
.Y(n_445)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_42),
.C(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_38),
.A2(n_133),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_51),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_42),
.B(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_45),
.B(n_54),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_50),
.B(n_53),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_49),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_51),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_51),
.A2(n_222),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_51),
.B(n_300),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_52),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_53),
.B(n_320),
.C(n_325),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_56),
.A2(n_339),
.B1(n_340),
.B2(n_342),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_56),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_56),
.B(n_109),
.C(n_339),
.Y(n_375)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_60),
.B(n_63),
.C(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_68),
.A2(n_69),
.B1(n_82),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_79),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_76),
.C(n_79),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_71),
.A2(n_78),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_71),
.A2(n_78),
.B1(n_95),
.B2(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_71),
.B(n_171),
.C(n_172),
.Y(n_254)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_77),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_83),
.C(n_94),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_83),
.B(n_241),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_84),
.A2(n_151),
.B1(n_156),
.B2(n_157),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_84),
.B(n_157),
.C(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_84),
.A2(n_91),
.B1(n_156),
.B2(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_88),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_90),
.Y(n_311)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_91),
.Y(n_213)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_95),
.Y(n_242)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_97),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_99),
.A2(n_136),
.B1(n_198),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_115),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_116),
.C(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

AOI21x1_ASAP7_75t_SL g191 ( 
.A1(n_102),
.A2(n_192),
.B(n_195),
.Y(n_191)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_106),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_106),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_106),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_114),
.Y(n_107)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_108),
.B(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_109),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_111),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_109),
.B(n_179),
.C(n_187),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_128),
.C(n_133),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_128),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_111),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_111),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_111),
.B(n_291),
.C(n_293),
.Y(n_364)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_113),
.Y(n_238)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_113),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_117),
.A2(n_141),
.B1(n_239),
.B2(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_184),
.C(n_239),
.Y(n_278)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_120),
.B(n_179),
.C(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_SL g377 ( 
.A(n_120),
.Y(n_377)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_132),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_147),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.C(n_144),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_147),
.B(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_149),
.C(n_197),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_158),
.A2(n_159),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_196),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_164),
.B(n_165),
.C(n_196),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_166),
.B(n_190),
.C(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_176),
.A2(n_186),
.B1(n_187),
.B2(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_176),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_179),
.A2(n_184),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_179),
.A2(n_184),
.B1(n_215),
.B2(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_181),
.Y(n_349)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_194),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_244),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_200),
.B(n_244),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_209),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_201),
.B(n_205),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_209),
.B(n_434),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_223),
.B(n_243),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_210),
.B(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_211),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_214),
.A2(n_219),
.B1(n_220),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_214),
.Y(n_409)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_240),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_224),
.B(n_240),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_236),
.C(n_239),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_225),
.A2(n_226),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_227),
.B(n_229),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_232),
.Y(n_388)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_235),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_260),
.Y(n_402)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g437 ( 
.A1(n_249),
.A2(n_274),
.B(n_438),
.C(n_441),
.D(n_443),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_272),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_251),
.B(n_442),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_269),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_255),
.C(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B1(n_262),
.B2(n_268),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_272),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_275),
.B(n_276),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_278),
.B(n_444),
.Y(n_443)
);

CKINVDCx11_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_414),
.B(n_428),
.C(n_435),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_390),
.B(n_413),
.Y(n_285)
);

NAND2x1p5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_365),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_317),
.C(n_343),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_297),
.C(n_303),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_312),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_329),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_330),
.C(n_337),
.Y(n_382)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx12f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_334),
.B(n_336),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_334),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_405),
.C(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_360),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_361),
.C(n_363),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_353),
.C(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_353),
.B1(n_358),
.B2(n_359),
.Y(n_350)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_353),
.Y(n_358)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_381),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_382),
.C(n_383),
.Y(n_412)
);

XOR2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_380),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_376),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_380),
.C(n_393),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_375),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_371),
.C(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_412),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_412),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_416),
.C(n_417),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_407),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_395),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_404),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_400),
.B2(n_403),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_398),
.Y(n_421)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_407),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_418),
.B1(n_429),
.B2(n_433),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.Y(n_418)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_419),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.C(n_422),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_433),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.C(n_432),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);


endmodule