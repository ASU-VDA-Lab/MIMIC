module fake_jpeg_10184_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_6),
.B(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_35),
.B1(n_33),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_50),
.B1(n_47),
.B2(n_21),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_47),
.B1(n_45),
.B2(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_69),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_35),
.B1(n_33),
.B2(n_20),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_37),
.B1(n_21),
.B2(n_31),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_73),
.B1(n_95),
.B2(n_96),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_89),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_38),
.B1(n_25),
.B2(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_38),
.B1(n_37),
.B2(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_84),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_56),
.B1(n_34),
.B2(n_26),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_36),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_30),
.B(n_19),
.Y(n_112)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_91),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_41),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_30),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_25),
.B1(n_37),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_37),
.B1(n_44),
.B2(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_126),
.B1(n_80),
.B2(n_97),
.Y(n_144)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_66),
.B1(n_65),
.B2(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_124),
.B1(n_83),
.B2(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_58),
.B(n_26),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_114),
.B(n_19),
.Y(n_147)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_107),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_34),
.B1(n_70),
.B2(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_121),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_41),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_52),
.B1(n_41),
.B2(n_42),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_75),
.B1(n_88),
.B2(n_84),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_139),
.B1(n_144),
.B2(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_121),
.C(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_145),
.C(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_116),
.B1(n_120),
.B2(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_148),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_70),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_99),
.B1(n_107),
.B2(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_151),
.B1(n_39),
.B2(n_40),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_149),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_87),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_124),
.B1(n_123),
.B2(n_114),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_80),
.B1(n_81),
.B2(n_18),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_119),
.B1(n_28),
.B2(n_32),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_147),
.B(n_150),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_179),
.B(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_162),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_114),
.C(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_111),
.B1(n_116),
.B2(n_118),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_167),
.B1(n_184),
.B2(n_23),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_41),
.Y(n_165)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_30),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_40),
.C(n_39),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_81),
.B1(n_91),
.B2(n_103),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_180),
.B1(n_134),
.B2(n_137),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_149),
.B1(n_129),
.B2(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_175),
.B(n_176),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_119),
.B1(n_103),
.B2(n_40),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_42),
.C(n_40),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_53),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_140),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_12),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_189),
.B1(n_192),
.B2(n_206),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_141),
.B1(n_129),
.B2(n_134),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_177),
.B(n_137),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_208),
.B1(n_168),
.B2(n_179),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_173),
.B1(n_169),
.B2(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_195),
.B(n_203),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_49),
.B(n_53),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_204),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_53),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_32),
.B1(n_23),
.B2(n_22),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_42),
.B1(n_32),
.B2(n_23),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_188),
.C(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_30),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_22),
.B1(n_30),
.B2(n_10),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_160),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_165),
.C(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_183),
.C(n_175),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_234),
.C(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_228),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_201),
.B1(n_193),
.B2(n_197),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_206),
.B1(n_196),
.B2(n_2),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_158),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_162),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_204),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_176),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_203),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_22),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_191),
.B1(n_199),
.B2(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_195),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_261),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_260),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_220),
.B1(n_218),
.B2(n_240),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_0),
.B(n_1),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_9),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_220),
.CI(n_219),
.CON(n_264),
.SN(n_264)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_276),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_216),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_270),
.C(n_272),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_217),
.C(n_215),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_232),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_243),
.C(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_281),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_9),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_7),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_262),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_0),
.C(n_1),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_256),
.B(n_251),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_275),
.B(n_280),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_253),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_248),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_241),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_258),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_254),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_268),
.C(n_277),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_13),
.C(n_2),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_278),
.B1(n_250),
.B2(n_265),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_290),
.B1(n_285),
.B2(n_291),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_283),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_264),
.B(n_247),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_305),
.B(n_304),
.Y(n_318)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_247),
.A3(n_10),
.B1(n_11),
.B2(n_16),
.C(n_15),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_3),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_299),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_317),
.B1(n_0),
.B2(n_2),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_283),
.C(n_1),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_318),
.C(n_319),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_327),
.C(n_3),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_308),
.B(n_298),
.Y(n_322)
);

AOI321xp33_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_323),
.A3(n_324),
.B1(n_325),
.B2(n_3),
.C(n_4),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_300),
.B(n_13),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_311),
.B(n_4),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_330),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_320),
.B(n_4),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_3),
.B(n_4),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_6),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_6),
.B(n_322),
.Y(n_338)
);


endmodule