module fake_jpeg_5147_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_39),
.Y(n_43)
);

OR2x4_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_25),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_28),
.B(n_21),
.C(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_51),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_19),
.B1(n_39),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_53),
.B1(n_46),
.B2(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_32),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_56),
.B1(n_55),
.B2(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_32),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_59),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_17),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_72),
.B(n_49),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_75),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_50),
.B1(n_46),
.B2(n_57),
.Y(n_65)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_25),
.B1(n_32),
.B2(n_40),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_81),
.B1(n_18),
.B2(n_42),
.Y(n_96)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_74),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_42),
.B1(n_57),
.B2(n_26),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_26),
.B1(n_20),
.B2(n_31),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_37),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_37),
.CI(n_44),
.CON(n_104),
.SN(n_104)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_26),
.B1(n_40),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_44),
.B1(n_54),
.B2(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_54),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_43),
.B(n_52),
.Y(n_92)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_0),
.B1(n_31),
.B2(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_44),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_1),
.B(n_2),
.Y(n_128)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_96),
.B1(n_68),
.B2(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_77),
.C(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_64),
.A3(n_79),
.B1(n_76),
.B2(n_68),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_59),
.B(n_72),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_112),
.B1(n_123),
.B2(n_129),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_127),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_68),
.B1(n_69),
.B2(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_121),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_60),
.B(n_70),
.C(n_42),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_8),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_125),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_82),
.B1(n_18),
.B2(n_74),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_91),
.C(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_128),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_93),
.B(n_88),
.C(n_105),
.D(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_74),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_83),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_86),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_85),
.B1(n_83),
.B2(n_87),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_118),
.B1(n_109),
.B2(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_5),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_5),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_8),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_9),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_157),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_162),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_125),
.B1(n_119),
.B2(n_122),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_114),
.B1(n_108),
.B2(n_130),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_169),
.B1(n_153),
.B2(n_140),
.Y(n_188)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_109),
.B(n_127),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_150),
.B(n_134),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

OAI22x1_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_128),
.B1(n_131),
.B2(n_11),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_9),
.C(n_10),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_144),
.C(n_155),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_12),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_146),
.B(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_197),
.B1(n_176),
.B2(n_163),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_171),
.B1(n_149),
.B2(n_139),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_133),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_151),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_133),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_135),
.C(n_164),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_206),
.C(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_161),
.C(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_208),
.B1(n_188),
.B2(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_172),
.B1(n_161),
.B2(n_145),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_187),
.C(n_181),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_218),
.C(n_221),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_210),
.B1(n_201),
.B2(n_198),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_185),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_220),
.B(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_165),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_186),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.C(n_184),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_200),
.B(n_209),
.C(n_198),
.D(n_182),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_230),
.Y(n_234)
);

OAI321xp33_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_194),
.A3(n_192),
.B1(n_180),
.B2(n_191),
.C(n_208),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_178),
.B1(n_177),
.B2(n_189),
.Y(n_235)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_217),
.C(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_233),
.C(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_203),
.B1(n_217),
.B2(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_213),
.C(n_178),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_224),
.C(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_197),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_174),
.B(n_158),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_237),
.B(n_173),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_158),
.B1(n_174),
.B2(n_237),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_244),
.A2(n_13),
.B(n_14),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_13),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_248),
.Y(n_249)
);


endmodule