module fake_jpeg_14875_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_17),
.B1(n_24),
.B2(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_19),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_28),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_18),
.B(n_21),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_70),
.A2(n_29),
.B1(n_23),
.B2(n_18),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_62),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_43),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_43),
.B1(n_40),
.B2(n_51),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_30),
.B1(n_24),
.B2(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_35),
.C(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_22),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_109),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_114),
.B1(n_63),
.B2(n_47),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_69),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_122),
.B(n_68),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_50),
.B1(n_66),
.B2(n_46),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_46),
.B1(n_59),
.B2(n_42),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_92),
.B1(n_90),
.B2(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_84),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_22),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_29),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_91),
.B1(n_80),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_114),
.B1(n_108),
.B2(n_97),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_23),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_67),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_30),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_96),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_90),
.B1(n_76),
.B2(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_44),
.A3(n_42),
.B1(n_38),
.B2(n_27),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_54),
.B(n_38),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_106),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_54),
.C(n_82),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_85),
.B(n_27),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_27),
.B(n_31),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_120),
.B1(n_116),
.B2(n_112),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_104),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_159),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_164),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_169),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_178),
.B(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

OR2x2_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_115),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_177),
.B(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_111),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_111),
.C(n_82),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_126),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_144),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_150),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_185),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_142),
.B1(n_130),
.B2(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_191),
.B1(n_192),
.B2(n_207),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_142),
.B1(n_174),
.B2(n_131),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_132),
.B1(n_136),
.B2(n_138),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_148),
.B1(n_135),
.B2(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_124),
.C(n_149),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_204),
.C(n_209),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_126),
.B(n_150),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_102),
.B(n_160),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_172),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_57),
.B1(n_47),
.B2(n_68),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_181),
.C(n_170),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_161),
.CI(n_180),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_158),
.C(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_217),
.C(n_223),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_0),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_155),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_0),
.B(n_1),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_197),
.Y(n_217)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_164),
.B(n_162),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_228),
.B(n_193),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_162),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_227),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_159),
.C(n_73),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_169),
.B1(n_31),
.B2(n_32),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_235),
.B1(n_193),
.B2(n_187),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_73),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_195),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_225),
.Y(n_238)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_200),
.B1(n_202),
.B2(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_245),
.B1(n_248),
.B2(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_194),
.B(n_200),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_221),
.A2(n_194),
.B1(n_57),
.B2(n_111),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_16),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_215),
.B1(n_227),
.B2(n_210),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_211),
.B(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_1),
.B(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_1),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_212),
.C(n_210),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_266),
.C(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_231),
.C(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.C(n_273),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_228),
.C(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_247),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_236),
.B(n_214),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_4),
.C(n_5),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_237),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_255),
.C(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_283),
.C(n_268),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_255),
.C(n_256),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_259),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_239),
.C(n_256),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_242),
.B(n_249),
.Y(n_286)
);

XOR2x2_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_242),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_276),
.C(n_283),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_248),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_299),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_9),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_14),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_308),
.C(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_277),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_276),
.C(n_298),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_280),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_10),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_6),
.C(n_8),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

AOI31xp67_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_318),
.B(n_11),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_9),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_13),
.C(n_11),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_317),
.Y(n_324)
);

AOI321xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_321),
.A3(n_320),
.B1(n_313),
.B2(n_13),
.C(n_12),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.Y(n_327)
);


endmodule