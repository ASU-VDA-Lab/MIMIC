module fake_netlist_5_1106_n_3082 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_409, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_3082);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_3082;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_2771;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_3036;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_3010;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_3048;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2959;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_436;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_422;
wire n_1070;
wire n_777;
wire n_1547;
wire n_475;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_415;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_485;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_901;
wire n_553;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1556;
wire n_1384;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_2932;
wire n_2753;
wire n_464;
wire n_2980;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3025;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_586;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_2218;
wire n_2267;
wire n_1072;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_1276;
wire n_702;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_3042;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_1510;
wire n_1380;
wire n_624;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3003;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_3030;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3075;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_3031;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_457;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2729;
wire n_1820;
wire n_2261;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_513;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_2953;
wire n_824;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_1684;
wire n_921;
wire n_2658;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_3059;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_1630;
wire n_716;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_531;
wire n_3020;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_419;
wire n_1346;
wire n_3053;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_418;
wire n_968;
wire n_912;
wire n_451;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_515;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1631;
wire n_1203;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_2733;
wire n_455;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3041;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_3067;
wire n_1932;
wire n_2755;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_1594;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2393;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_2971;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_472;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_669;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_458;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_1499;
wire n_711;
wire n_3061;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_2988;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_3035;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_500;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_2692;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_416;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_620;
wire n_2430;
wire n_643;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_3070;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_508;
wire n_2186;
wire n_1320;
wire n_506;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_2748;
wire n_518;
wire n_505;
wire n_2057;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3081;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_428;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3017;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_3054;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_3050;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_2957;
wire n_839;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_2961;
wire n_413;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_2612;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_465;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_3004;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_453;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_3057;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_412;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_2938;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_2975;
wire n_438;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

BUFx3_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_155),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_50),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_160),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_175),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_79),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_52),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_286),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_310),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_130),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_206),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_191),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_186),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_84),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_67),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_348),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_149),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_121),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_326),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_15),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_324),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_197),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_46),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_156),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_336),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_205),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_300),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_2),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_215),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_183),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_91),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_275),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_357),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_145),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_226),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_266),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_235),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_118),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_279),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_292),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_271),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_52),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_238),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_289),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_40),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_48),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_62),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_364),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_78),
.Y(n_467)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_146),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_95),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_245),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_246),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_314),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_337),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_239),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_353),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_90),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_399),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_304),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_263),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_13),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_372),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_201),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_228),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_192),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_80),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_177),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_296),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_354),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_268),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_247),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_356),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_63),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_105),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_77),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_397),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_378),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_126),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_302),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_117),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_89),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_234),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_129),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_1),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_159),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_142),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_62),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_408),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g509 ( 
.A(n_28),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_44),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_233),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_377),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_317),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_398),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_251),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_57),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_178),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_313),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_120),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_135),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_26),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_164),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_132),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_71),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_213),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_184),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_148),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_359),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_57),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_207),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_95),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_55),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_391),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_127),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_403),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_5),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_406),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_298),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_89),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_209),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_64),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_250),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_217),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_38),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_31),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_311),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_241),
.Y(n_548)
);

BUFx2_ASAP7_75t_R g549 ( 
.A(n_322),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_396),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_131),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_59),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_158),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_144),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_193),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_74),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_151),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_389),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_351),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_154),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_393),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_38),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_5),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_200),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_129),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_280),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_19),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_77),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_16),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_407),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_249),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_63),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_196),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_94),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_194),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_227),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_375),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_306),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_273),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_190),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_366),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_257),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_285),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_260),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_299),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_157),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_139),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_140),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_320),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_150),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_182),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_86),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_138),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_203),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_363),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_46),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_171),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_256),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_39),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_60),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_288),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_404),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_136),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_297),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_360),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_100),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_109),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_222),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_19),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_242),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_409),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_58),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_365),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_381),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_290),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_64),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_338),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_333),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_316),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_305),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_390),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_73),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_42),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_34),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_42),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_98),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_143),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_291),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_167),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_115),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_283),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_17),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_49),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_332),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_162),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_4),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_120),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_94),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_172),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_189),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_410),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_72),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_405),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_259),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_6),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_0),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_84),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_328),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_61),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_301),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_79),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_23),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_220),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_400),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_86),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_214),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_202),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_368),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_80),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_240),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_319),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_373),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_161),
.Y(n_663)
);

CKINVDCx14_ASAP7_75t_R g664 ( 
.A(n_61),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_125),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_87),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_48),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_237),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_342),
.Y(n_669)
);

BUFx2_ASAP7_75t_R g670 ( 
.A(n_110),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_165),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_99),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_248),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_124),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_153),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_36),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_91),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_90),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_344),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_35),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_176),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_261),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_369),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_47),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_101),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_388),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_45),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_303),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_36),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_12),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_137),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_92),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_60),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_181),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_16),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_284),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_23),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_22),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_258),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_295),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_72),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_169),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_2),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_168),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_83),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_188),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_252),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_98),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_294),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_225),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_392),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_13),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_312),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_29),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_70),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_12),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_500),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_509),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_509),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_509),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_509),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_509),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_416),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_509),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_664),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_569),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_419),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_509),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_414),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_430),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_674),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

INVxp33_ASAP7_75t_SL g733 ( 
.A(n_596),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_468),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_521),
.Y(n_735)
);

CKINVDCx14_ASAP7_75t_R g736 ( 
.A(n_686),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_521),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_521),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_418),
.B(n_0),
.Y(n_739)
);

BUFx2_ASAP7_75t_SL g740 ( 
.A(n_429),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_414),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_521),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_525),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_525),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_532),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_525),
.Y(n_746)
);

INVxp33_ASAP7_75t_SL g747 ( 
.A(n_701),
.Y(n_747)
);

INVxp33_ASAP7_75t_L g748 ( 
.A(n_545),
.Y(n_748)
);

INVxp33_ASAP7_75t_SL g749 ( 
.A(n_435),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_525),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_562),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_562),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_562),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_562),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_651),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_468),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_676),
.Y(n_757)
);

CKINVDCx14_ASAP7_75t_R g758 ( 
.A(n_457),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_676),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_489),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_411),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_468),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_411),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_468),
.Y(n_764)
);

INVxp33_ASAP7_75t_SL g765 ( 
.A(n_435),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_694),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_422),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_676),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_676),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_420),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_421),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_532),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_546),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_708),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_426),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_429),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_445),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_492),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_448),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_463),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_465),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_423),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_546),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_467),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_477),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_441),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_501),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_504),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_507),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_687),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_468),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_687),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_623),
.Y(n_793)
);

INVxp33_ASAP7_75t_SL g794 ( 
.A(n_431),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_455),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_623),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_510),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_460),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_520),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_437),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_530),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_535),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_551),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_565),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_492),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_464),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_592),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_603),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_441),
.Y(n_809)
);

INVxp33_ASAP7_75t_L g810 ( 
.A(n_486),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_469),
.Y(n_811)
);

INVxp33_ASAP7_75t_SL g812 ( 
.A(n_481),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_603),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_607),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_632),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_493),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_494),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_473),
.Y(n_818)
);

BUFx2_ASAP7_75t_SL g819 ( 
.A(n_453),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_638),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_453),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_680),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_611),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_685),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_468),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_495),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_697),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_458),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_698),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_473),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_425),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_498),
.Y(n_833)
);

INVxp33_ASAP7_75t_SL g834 ( 
.A(n_503),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_468),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_473),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

INVxp33_ASAP7_75t_SL g838 ( 
.A(n_517),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_712),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_412),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_415),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_427),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_434),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_548),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_443),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_458),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_437),
.Y(n_847)
);

CKINVDCx16_ASAP7_75t_R g848 ( 
.A(n_462),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_454),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_459),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_461),
.Y(n_851)
);

INVxp33_ASAP7_75t_L g852 ( 
.A(n_486),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_527),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_428),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_612),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_813),
.Y(n_856)
);

BUFx8_ASAP7_75t_L g857 ( 
.A(n_798),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_726),
.Y(n_858)
);

AND3x2_ASAP7_75t_L g859 ( 
.A(n_739),
.B(n_625),
.C(n_612),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_733),
.A2(n_480),
.B1(n_534),
.B2(n_462),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_818),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_813),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_818),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_822),
.B(n_450),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_723),
.B(n_450),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_718),
.A2(n_720),
.B(n_719),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_818),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_831),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_809),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_831),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_721),
.A2(n_417),
.B(n_413),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_722),
.A2(n_728),
.B(n_724),
.Y(n_872)
);

CKINVDCx11_ASAP7_75t_R g873 ( 
.A(n_729),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_734),
.A2(n_417),
.B(n_413),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_831),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_831),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_725),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_761),
.B(n_440),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_735),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_726),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_836),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_725),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_766),
.B(n_452),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_734),
.A2(n_471),
.B(n_452),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_756),
.A2(n_491),
.B(n_471),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_737),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_836),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_738),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_740),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_742),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_763),
.B(n_440),
.Y(n_892)
);

OA21x2_ASAP7_75t_L g893 ( 
.A1(n_756),
.A2(n_554),
.B(n_491),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_822),
.B(n_547),
.Y(n_894)
);

OA21x2_ASAP7_75t_L g895 ( 
.A1(n_762),
.A2(n_598),
.B(n_554),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_743),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_744),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_733),
.A2(n_534),
.B1(n_561),
.B2(n_480),
.Y(n_898)
);

OA21x2_ASAP7_75t_L g899 ( 
.A1(n_762),
.A2(n_707),
.B(n_598),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_727),
.B(n_547),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_746),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_750),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_767),
.B(n_650),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_782),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_730),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_751),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_778),
.B(n_599),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_752),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_753),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_754),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_822),
.Y(n_911)
);

BUFx8_ASAP7_75t_SL g912 ( 
.A(n_729),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_758),
.B(n_650),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_824),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_730),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_757),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_805),
.B(n_599),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_759),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_808),
.B(n_707),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_824),
.B(n_710),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_768),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_764),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_747),
.A2(n_629),
.B1(n_658),
.B2(n_561),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_840),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_841),
.B(n_710),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_791),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_826),
.A2(n_835),
.B(n_843),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_853),
.B(n_484),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_826),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_835),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_832),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_845),
.B(n_488),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_849),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_850),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_747),
.A2(n_524),
.B1(n_533),
.B2(n_522),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_851),
.B(n_511),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_771),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_731),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_775),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_819),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_777),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_779),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_780),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_781),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_784),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_833),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_787),
.Y(n_951)
);

BUFx8_ASAP7_75t_SL g952 ( 
.A(n_741),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_788),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_810),
.B(n_606),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_758),
.A2(n_658),
.B1(n_660),
.B2(n_629),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_844),
.B(n_512),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_789),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_797),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_799),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_801),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_842),
.B(n_519),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_803),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_804),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_732),
.B(n_531),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_807),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_854),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_736),
.B(n_541),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_806),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_814),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_717),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_815),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_820),
.B(n_543),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_823),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_800),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_940),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_925),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_928),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_944),
.Y(n_979)
);

BUFx8_ASAP7_75t_L g980 ( 
.A(n_877),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_961),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_954),
.B(n_810),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_962),
.B(n_736),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_972),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_926),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_925),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_863),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_941),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_931),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_928),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_919),
.B(n_865),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_SL g992 ( 
.A(n_877),
.B(n_549),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_863),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_935),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_935),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_935),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_931),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_856),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_928),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_919),
.B(n_760),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_935),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_919),
.B(n_900),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_922),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_922),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_922),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_932),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_882),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_932),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_935),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_954),
.B(n_852),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_928),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_936),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_936),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_932),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_936),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_936),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_936),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_975),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_929),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_SL g1020 ( 
.A(n_883),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_929),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_965),
.B(n_825),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_863),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_890),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_939),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_929),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_928),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_939),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_939),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_889),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_889),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_939),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_901),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_939),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_942),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_883),
.B(n_473),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_867),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_942),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_867),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_901),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_909),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_874),
.A2(n_558),
.B(n_553),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_856),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_942),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_867),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_878),
.B(n_852),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_903),
.B(n_794),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_909),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_882),
.B(n_904),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_910),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_942),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_942),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_956),
.B(n_555),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_873),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_948),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_862),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_910),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_948),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_948),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_948),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_867),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_948),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_916),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_956),
.B(n_555),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_953),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_890),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_953),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_916),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_872),
.A2(n_560),
.B(n_559),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_924),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_876),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_876),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_924),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_956),
.B(n_794),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_868),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_953),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_878),
.B(n_855),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_876),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_953),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_911),
.B(n_555),
.Y(n_1080)
);

INVxp33_ASAP7_75t_L g1081 ( 
.A(n_913),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_872),
.A2(n_579),
.B(n_578),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_953),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_SL g1084 ( 
.A1(n_860),
.A2(n_829),
.B1(n_846),
.B2(n_809),
.Y(n_1084)
);

XNOR2xp5_ASAP7_75t_L g1085 ( 
.A(n_898),
.B(n_829),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_975),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_957),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_957),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_965),
.B(n_828),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_957),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_868),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_876),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_875),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_911),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_949),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_892),
.B(n_855),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_943),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_875),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_957),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_960),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_960),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_960),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_911),
.B(n_555),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_887),
.B(n_812),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_888),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_862),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_881),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_965),
.B(n_830),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_960),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_881),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_960),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_891),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_966),
.Y(n_1114)
);

XNOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_923),
.B(n_846),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_966),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_911),
.B(n_581),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_891),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_874),
.A2(n_594),
.B(n_591),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_891),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_891),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_888),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_966),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_966),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_914),
.Y(n_1125)
);

XOR2xp5_ASAP7_75t_L g1126 ( 
.A(n_955),
.B(n_741),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_892),
.B(n_811),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_966),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_891),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_914),
.B(n_837),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_973),
.B(n_839),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_943),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_970),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_970),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_911),
.B(n_581),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_970),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_897),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_970),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_970),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1003),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1081),
.B(n_1047),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1125),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_991),
.A2(n_774),
.B1(n_626),
.B2(n_646),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1019),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1046),
.B(n_933),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1003),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_976),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_982),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_979),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_1125),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1004),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1046),
.B(n_949),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1130),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1077),
.B(n_933),
.Y(n_1154)
);

AND2x6_ASAP7_75t_L g1155 ( 
.A(n_1019),
.B(n_864),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1004),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_981),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1130),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_982),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1021),
.B(n_866),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_998),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1005),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1077),
.B(n_1096),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1096),
.B(n_907),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1074),
.B(n_776),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1021),
.B(n_866),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1005),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1010),
.B(n_907),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1010),
.B(n_933),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1006),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1081),
.B(n_967),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1006),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1026),
.B(n_866),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1130),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1026),
.B(n_893),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1127),
.B(n_967),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1127),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1002),
.B(n_967),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1018),
.B(n_786),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1000),
.B(n_893),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1008),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_977),
.B(n_893),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1075),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_984),
.Y(n_1184)
);

NOR2x1p5_ASAP7_75t_L g1185 ( 
.A(n_1024),
.B(n_904),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1086),
.B(n_821),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_985),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1105),
.B(n_968),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1024),
.B(n_917),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1036),
.A2(n_626),
.B1(n_646),
.B2(n_606),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1066),
.B(n_917),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1131),
.B(n_1022),
.Y(n_1192)
);

INVxp33_ASAP7_75t_SL g1193 ( 
.A(n_1049),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1075),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1066),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_977),
.B(n_895),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_988),
.B(n_864),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_986),
.B(n_895),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_983),
.B(n_969),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_998),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_1097),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1043),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_986),
.B(n_895),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_L g1204 ( 
.A(n_1036),
.B(n_1095),
.C(n_1043),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1030),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1030),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1031),
.Y(n_1207)
);

NOR2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1097),
.B(n_853),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1132),
.B(n_905),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1056),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1014),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1126),
.A2(n_937),
.B1(n_677),
.B2(n_540),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_989),
.B(n_899),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1020),
.B(n_660),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_1132),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1107),
.B(n_848),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1031),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1033),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1033),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1040),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_989),
.B(n_899),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1040),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1020),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1041),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_980),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1041),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1020),
.B(n_812),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1014),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1048),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_980),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1131),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1084),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1022),
.Y(n_1233)
);

NOR2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1131),
.B(n_542),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_994),
.B(n_915),
.Y(n_1235)
);

AND2x2_ASAP7_75t_SL g1236 ( 
.A(n_992),
.B(n_858),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_980),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1022),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1091),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1089),
.B(n_827),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1089),
.B(n_858),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1048),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1089),
.B(n_816),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_997),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1053),
.B(n_871),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_978),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1109),
.A2(n_880),
.B1(n_938),
.B2(n_934),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1109),
.B(n_827),
.Y(n_1248)
);

BUFx8_ASAP7_75t_SL g1249 ( 
.A(n_1007),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1050),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1109),
.A2(n_880),
.B1(n_938),
.B2(n_934),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_993),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1053),
.A2(n_1064),
.B1(n_996),
.B2(n_1001),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1064),
.B(n_834),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1007),
.Y(n_1255)
);

BUFx4f_ASAP7_75t_L g1256 ( 
.A(n_1042),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1085),
.A2(n_677),
.B1(n_755),
.B2(n_748),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1085),
.B(n_817),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1050),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_995),
.A2(n_938),
.B1(n_934),
.B2(n_838),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1115),
.B(n_748),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1115),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1009),
.A2(n_871),
.B1(n_894),
.B2(n_864),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1012),
.B(n_834),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1013),
.B(n_838),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1091),
.Y(n_1267)
);

INVx8_ASAP7_75t_L g1268 ( 
.A(n_987),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1057),
.B(n_755),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1015),
.A2(n_871),
.B1(n_894),
.B2(n_973),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1054),
.B(n_670),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1016),
.B(n_749),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1007),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1063),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_993),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1063),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1068),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1126),
.B(n_971),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1093),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1068),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1070),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_L g1282 ( 
.A(n_1017),
.B(n_432),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_978),
.B(n_749),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_978),
.B(n_990),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1073),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_990),
.B(n_765),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1073),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_990),
.B(n_765),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1093),
.Y(n_1289)
);

AND2x2_ASAP7_75t_SL g1290 ( 
.A(n_1042),
.B(n_790),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1099),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1099),
.B(n_792),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1108),
.B(n_847),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1108),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1042),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1111),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1111),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1025),
.B(n_920),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1028),
.B(n_920),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_999),
.Y(n_1300)
);

AO22x2_ASAP7_75t_L g1301 ( 
.A1(n_1080),
.A2(n_616),
.B1(n_665),
.B2(n_537),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_999),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1029),
.B(n_920),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_999),
.B(n_894),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_993),
.Y(n_1305)
);

XNOR2x2_ASAP7_75t_L g1306 ( 
.A(n_1080),
.B(n_692),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_993),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1011),
.B(n_745),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1027),
.B(n_884),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1104),
.B(n_552),
.Y(n_1310)
);

INVx4_ASAP7_75t_SL g1311 ( 
.A(n_1094),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1032),
.A2(n_973),
.B1(n_927),
.B2(n_601),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1039),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1027),
.B(n_884),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1119),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1027),
.B(n_745),
.Y(n_1316)
);

NAND2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1104),
.B(n_556),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1119),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1119),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1034),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1035),
.B(n_930),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1038),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1044),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1069),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1113),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1051),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1177),
.B(n_693),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1144),
.B(n_1052),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1177),
.B(n_958),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1144),
.B(n_1055),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1299),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1141),
.B(n_772),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1171),
.B(n_772),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1303),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1178),
.B(n_1058),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1163),
.A2(n_1059),
.B1(n_1062),
.B2(n_1060),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1233),
.B(n_857),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1148),
.B(n_773),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1164),
.B(n_1065),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1281),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1195),
.B(n_1227),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1168),
.B(n_1067),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1233),
.B(n_857),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1148),
.B(n_1076),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1205),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1159),
.B(n_1079),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1161),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1183),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1206),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1194),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1159),
.B(n_1083),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1190),
.A2(n_1135),
.B(n_1117),
.C(n_974),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1252),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1207),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1200),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1214),
.A2(n_783),
.B1(n_793),
.B2(n_773),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_SL g1357 ( 
.A(n_1236),
.B(n_527),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1225),
.B(n_625),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1264),
.B(n_1087),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1233),
.B(n_857),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1217),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1290),
.A2(n_1088),
.B1(n_1098),
.B2(n_1090),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1270),
.B(n_1100),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1175),
.A2(n_1082),
.B(n_1069),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1200),
.B(n_783),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1283),
.B(n_1101),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1269),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_L g1368 ( 
.A(n_1197),
.B(n_1102),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1142),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1286),
.B(n_1103),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_L g1371 ( 
.A(n_1254),
.B(n_958),
.Y(n_1371)
);

AND2x6_ASAP7_75t_L g1372 ( 
.A(n_1315),
.B(n_1318),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1150),
.B(n_958),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1218),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1288),
.B(n_1293),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1231),
.B(n_433),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1152),
.A2(n_1204),
.B1(n_1155),
.B2(n_1190),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1292),
.B(n_1110),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1219),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1231),
.B(n_1153),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1160),
.B(n_1112),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1241),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1243),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1153),
.B(n_433),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1298),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1189),
.B(n_793),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1220),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1298),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1188),
.A2(n_1117),
.B(n_1135),
.C(n_974),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1194),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_L g1391 ( 
.A(n_1197),
.B(n_1114),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1202),
.B(n_796),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_L g1393 ( 
.A(n_1150),
.B(n_974),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1202),
.B(n_796),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1204),
.A2(n_1116),
.B1(n_1124),
.B2(n_1123),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1175),
.A2(n_1166),
.B(n_1160),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1153),
.B(n_436),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1166),
.B(n_1128),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1191),
.B(n_869),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1173),
.A2(n_1082),
.B(n_1133),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1165),
.B(n_945),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1239),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1249),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1199),
.B(n_869),
.Y(n_1404)
);

NOR2xp67_ASAP7_75t_L g1405 ( 
.A(n_1240),
.B(n_1134),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1179),
.B(n_945),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1142),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1173),
.B(n_1136),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1252),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1192),
.B(n_436),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1176),
.B(n_873),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1145),
.B(n_912),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1321),
.B(n_1138),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1239),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1192),
.B(n_438),
.Y(n_1415)
);

BUFx5_ASAP7_75t_L g1416 ( 
.A(n_1155),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1155),
.A2(n_1139),
.B1(n_927),
.B2(n_602),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1222),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1186),
.B(n_946),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1257),
.A2(n_568),
.B1(n_572),
.B2(n_567),
.C(n_563),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1238),
.B(n_438),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1154),
.B(n_912),
.Y(n_1422)
);

BUFx5_ASAP7_75t_L g1423 ( 
.A(n_1155),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1224),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1267),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1226),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_L g1427 ( 
.A(n_1197),
.B(n_1113),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1185),
.B(n_1234),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1210),
.B(n_859),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1267),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1279),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1158),
.B(n_439),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1216),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1169),
.B(n_1248),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1147),
.B(n_1039),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1158),
.B(n_439),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1229),
.Y(n_1437)
);

NOR3xp33_ASAP7_75t_L g1438 ( 
.A(n_1257),
.B(n_447),
.C(n_424),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1242),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1279),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1325),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1201),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1259),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1313),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1149),
.B(n_1039),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1250),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1142),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1174),
.B(n_442),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1274),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1157),
.B(n_1045),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1268),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1258),
.B(n_1262),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1252),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1143),
.A2(n_1180),
.B(n_1319),
.C(n_1295),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1308),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1184),
.B(n_1045),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1256),
.A2(n_885),
.B(n_605),
.C(n_610),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1214),
.B(n_952),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1187),
.B(n_1061),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1247),
.B(n_442),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1180),
.B(n_1061),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1304),
.B(n_1061),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1251),
.B(n_688),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1276),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1304),
.B(n_1071),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1277),
.B(n_1280),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1285),
.B(n_1287),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1143),
.A2(n_950),
.B1(n_951),
.B2(n_947),
.C(n_946),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1260),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1316),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1209),
.B(n_952),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1291),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1295),
.B(n_1071),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1320),
.B(n_688),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1375),
.B(n_1301),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1377),
.A2(n_1245),
.B1(n_1256),
.B2(n_1253),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1355),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1438),
.A2(n_1212),
.B1(n_1232),
.B2(n_1301),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1357),
.A2(n_1212),
.B1(n_1306),
.B2(n_1197),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1466),
.Y(n_1480)
);

NAND2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1451),
.B(n_1275),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1347),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1467),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1332),
.B(n_1263),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1348),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1434),
.B(n_1261),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1345),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1349),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1354),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1378),
.B(n_1235),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1377),
.B(n_1371),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1407),
.Y(n_1492)
);

AOI211xp5_ASAP7_75t_L g1493 ( 
.A1(n_1356),
.A2(n_1333),
.B(n_1452),
.C(n_1338),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1455),
.B(n_1263),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1451),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1357),
.A2(n_1278),
.B1(n_1323),
.B2(n_1322),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1367),
.B(n_1201),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1470),
.B(n_1193),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1361),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1331),
.B(n_1319),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1382),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1334),
.B(n_1244),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1458),
.A2(n_1271),
.B1(n_1225),
.B2(n_1223),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1453),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1374),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1383),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1369),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1339),
.A2(n_1326),
.B1(n_1245),
.B2(n_1317),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1346),
.B(n_1351),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_SL g1510 ( 
.A(n_1420),
.B(n_1272),
.C(n_1266),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1379),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1329),
.B(n_1312),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1350),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1406),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1396),
.B(n_1265),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1386),
.Y(n_1516)
);

A2O1A1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1454),
.A2(n_1310),
.B(n_1146),
.C(n_1151),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1327),
.B(n_1215),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1403),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_SL g1521 ( 
.A(n_1399),
.B(n_1271),
.C(n_571),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1404),
.A2(n_1208),
.B1(n_1282),
.B2(n_1215),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1390),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1380),
.B(n_1275),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1402),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1416),
.B(n_1423),
.Y(n_1526)
);

OR2x2_ASAP7_75t_SL g1527 ( 
.A(n_1401),
.B(n_1230),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1407),
.B(n_1223),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1365),
.A2(n_1237),
.B1(n_1273),
.B2(n_574),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1418),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1407),
.B(n_1311),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1416),
.B(n_1313),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1424),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1342),
.B(n_1140),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1426),
.Y(n_1535)
);

AND2x4_ASAP7_75t_SL g1536 ( 
.A(n_1447),
.B(n_1255),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1437),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1414),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1392),
.A2(n_437),
.B1(n_564),
.B2(n_527),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1344),
.B(n_1156),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1453),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1439),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1447),
.B(n_1311),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1447),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1443),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1453),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1372),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1341),
.B(n_1246),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1425),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1416),
.B(n_1162),
.Y(n_1550)
);

OAI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1394),
.A2(n_609),
.B(n_600),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1449),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1413),
.B(n_1167),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1430),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1340),
.B(n_1385),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1464),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1416),
.B(n_1170),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1472),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1419),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1433),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1509),
.B(n_1441),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1487),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1560),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1488),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1547),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1555),
.B(n_1531),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1480),
.B(n_1441),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1483),
.B(n_1405),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1547),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1547),
.Y(n_1572)
);

NAND2xp33_ASAP7_75t_L g1573 ( 
.A(n_1486),
.B(n_1416),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1489),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1555),
.B(n_1385),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1499),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1493),
.B(n_1411),
.C(n_1471),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1388),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1482),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1505),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1511),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1514),
.B(n_1366),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1490),
.B(n_1370),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1516),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1484),
.B(n_1474),
.Y(n_1586)
);

AND3x1_ASAP7_75t_SL g1587 ( 
.A(n_1478),
.B(n_1468),
.C(n_644),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_R g1588 ( 
.A(n_1520),
.B(n_1442),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1559),
.B(n_1388),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1518),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1484),
.B(n_1412),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1539),
.B(n_1422),
.C(n_1460),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1507),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1477),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1477),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1530),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1475),
.B(n_1381),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1543),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1494),
.B(n_1398),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1494),
.B(n_1410),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1533),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1501),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_L g1605 ( 
.A(n_1476),
.B(n_1423),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1535),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1491),
.A2(n_1335),
.B1(n_1363),
.B2(n_1359),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1544),
.Y(n_1608)
);

CKINVDCx8_ASAP7_75t_R g1609 ( 
.A(n_1546),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1546),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1541),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1537),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1566),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1607),
.A2(n_1491),
.B(n_1584),
.Y(n_1615)
);

A2O1A1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1592),
.A2(n_1479),
.B(n_1510),
.C(n_1539),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1591),
.B(n_1498),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1584),
.A2(n_1400),
.B(n_1364),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1601),
.B(n_1519),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1599),
.B(n_1515),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1570),
.A2(n_1526),
.B(n_1550),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1605),
.A2(n_1427),
.B(n_1391),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1565),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1605),
.A2(n_1368),
.B(n_1461),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1478),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1573),
.A2(n_1526),
.B(n_1268),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1570),
.A2(n_1557),
.B(n_1550),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1569),
.A2(n_1517),
.B(n_1457),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1573),
.A2(n_1508),
.B(n_1362),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1570),
.A2(n_1557),
.B(n_1532),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1572),
.A2(n_1532),
.B(n_1465),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1574),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1577),
.A2(n_1508),
.B(n_1610),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1561),
.A2(n_1268),
.B(n_1328),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1588),
.Y(n_1637)
);

OA22x2_ASAP7_75t_L g1638 ( 
.A1(n_1585),
.A2(n_1522),
.B1(n_1343),
.B2(n_1360),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1567),
.B(n_1563),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1568),
.A2(n_1330),
.B(n_1408),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1564),
.B(n_1527),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1580),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1576),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1586),
.A2(n_1362),
.B(n_1336),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1576),
.A2(n_1336),
.B(n_1462),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1572),
.A2(n_1324),
.B(n_1534),
.Y(n_1646)
);

AND3x1_ASAP7_75t_L g1647 ( 
.A(n_1594),
.B(n_1479),
.C(n_1496),
.Y(n_1647)
);

AND3x2_ASAP7_75t_L g1648 ( 
.A(n_1564),
.B(n_1429),
.C(n_1541),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1567),
.B(n_1496),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1572),
.A2(n_1324),
.B(n_1553),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1562),
.A2(n_1436),
.B(n_1432),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1590),
.A2(n_1510),
.B(n_1521),
.C(n_1551),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1590),
.A2(n_1503),
.B1(n_1558),
.B2(n_1545),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1603),
.A2(n_1503),
.B1(n_1556),
.B2(n_1552),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_SL g1655 ( 
.A(n_1566),
.B(n_1497),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1603),
.Y(n_1656)
);

AO31x2_ASAP7_75t_L g1657 ( 
.A1(n_1581),
.A2(n_1473),
.A3(n_1540),
.B(n_1314),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1582),
.A2(n_1314),
.B(n_1309),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1575),
.A2(n_1521),
.B1(n_1529),
.B2(n_1428),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1583),
.A2(n_1358),
.B1(n_1337),
.B2(n_1512),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1580),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1609),
.B(n_1255),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1598),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1642),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1637),
.Y(n_1665)
);

BUFx2_ASAP7_75t_R g1666 ( 
.A(n_1619),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1618),
.A2(n_1524),
.B(n_1309),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_R g1668 ( 
.A(n_1662),
.B(n_1609),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1639),
.B(n_1567),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1661),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1649),
.B(n_1612),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1620),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1657),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1614),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1595),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1621),
.B(n_1635),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1624),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1616),
.B(n_1384),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1614),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1662),
.B(n_1593),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1615),
.B(n_1566),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_1397),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1635),
.B(n_1566),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1623),
.A2(n_1571),
.B(n_1566),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1644),
.A2(n_564),
.B1(n_634),
.B2(n_631),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1652),
.A2(n_1415),
.B(n_1448),
.C(n_1421),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1625),
.A2(n_1571),
.B(n_1548),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1653),
.A2(n_1463),
.B(n_1376),
.C(n_1528),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1641),
.B(n_1606),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1628),
.A2(n_1633),
.B(n_1622),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1631),
.A2(n_1571),
.B(n_1597),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1644),
.B(n_1571),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1626),
.B(n_1596),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1631),
.A2(n_885),
.B(n_1395),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1634),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_SL g1699 ( 
.A(n_1653),
.B(n_1571),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1640),
.A2(n_1597),
.B(n_1417),
.Y(n_1700)
);

CKINVDCx11_ASAP7_75t_R g1701 ( 
.A(n_1656),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1643),
.B(n_1589),
.Y(n_1702)
);

INVx6_ASAP7_75t_SL g1703 ( 
.A(n_1648),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1663),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1657),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1638),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1621),
.B(n_1575),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1638),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1654),
.B(n_1575),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1654),
.B(n_1542),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1657),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1615),
.B(n_1655),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1645),
.B(n_1593),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1659),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1630),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1651),
.B(n_1579),
.Y(n_1716)
);

BUFx12f_ASAP7_75t_L g1717 ( 
.A(n_1636),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1646),
.B(n_1650),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1658),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1629),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1663),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1620),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1617),
.A2(n_1358),
.B1(n_1524),
.B2(n_1604),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1639),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1649),
.B(n_1579),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1649),
.B(n_1600),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1657),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1663),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1637),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1649),
.B(n_1600),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1639),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_SL g1734 ( 
.A(n_1637),
.B(n_1495),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1620),
.Y(n_1735)
);

BUFx8_ASAP7_75t_L g1736 ( 
.A(n_1642),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1663),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1623),
.A2(n_1597),
.B(n_1417),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1623),
.A2(n_1597),
.B(n_1495),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1657),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1663),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1641),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1620),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1619),
.B(n_1485),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1617),
.B(n_1600),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1620),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1616),
.A2(n_1358),
.B(n_1502),
.C(n_597),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1649),
.B(n_1513),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1678),
.B(n_654),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1675),
.B(n_1608),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_656),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1718),
.A2(n_1597),
.B(n_1409),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1688),
.A2(n_624),
.B1(n_630),
.B2(n_622),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1677),
.B(n_663),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1741),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1741),
.B(n_927),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1701),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1701),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1692),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1672),
.B(n_1578),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_SL g1762 ( 
.A1(n_1680),
.A2(n_950),
.B(n_951),
.C(n_947),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1688),
.A2(n_636),
.B1(n_637),
.B2(n_633),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

NOR2xp67_ASAP7_75t_L g1765 ( 
.A(n_1664),
.B(n_1506),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1742),
.B(n_673),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1736),
.Y(n_1767)
);

AOI21x1_ASAP7_75t_SL g1768 ( 
.A1(n_1683),
.A2(n_1445),
.B(n_1435),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1727),
.B(n_1578),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1723),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1714),
.A2(n_645),
.B1(n_647),
.B2(n_642),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1666),
.B(n_1563),
.Y(n_1772)
);

O2A1O1Ixp5_ASAP7_75t_L g1773 ( 
.A1(n_1680),
.A2(n_683),
.B(n_702),
.C(n_675),
.Y(n_1773)
);

A2O1A1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1685),
.A2(n_1352),
.B(n_1536),
.C(n_711),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1730),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_SL g1776 ( 
.A1(n_1685),
.A2(n_959),
.B(n_964),
.C(n_963),
.Y(n_1776)
);

NOR2xp67_ASAP7_75t_L g1777 ( 
.A(n_1670),
.B(n_1395),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1717),
.B(n_1523),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1748),
.B(n_706),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1744),
.B(n_649),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1737),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1747),
.A2(n_1689),
.B(n_1691),
.C(n_1713),
.Y(n_1782)
);

OR2x2_ASAP7_75t_SL g1783 ( 
.A(n_1712),
.B(n_959),
.Y(n_1783)
);

AOI221x1_ASAP7_75t_L g1784 ( 
.A1(n_1725),
.A2(n_621),
.B1(n_640),
.B2(n_590),
.C(n_581),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1693),
.A2(n_879),
.B(n_1294),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1716),
.Y(n_1786)
);

O2A1O1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1710),
.A2(n_608),
.B(n_502),
.C(n_1389),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1673),
.B(n_1578),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1673),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1702),
.B(n_652),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1696),
.B(n_655),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1719),
.Y(n_1792)
);

OR2x6_ASAP7_75t_SL g1793 ( 
.A(n_1665),
.B(n_659),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1718),
.A2(n_879),
.B(n_1296),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1695),
.B(n_963),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1728),
.B(n_1578),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1745),
.B(n_666),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1679),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1679),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1705),
.A2(n_1456),
.B(n_1450),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1745),
.B(n_667),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1698),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1698),
.Y(n_1803)
);

NOR2xp67_ASAP7_75t_L g1804 ( 
.A(n_1708),
.B(n_1525),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1724),
.B(n_1735),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1724),
.B(n_1578),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1708),
.A2(n_678),
.B1(n_684),
.B2(n_672),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1695),
.B(n_964),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1706),
.A2(n_690),
.B1(n_695),
.B2(n_689),
.Y(n_1809)
);

NOR2xp67_ASAP7_75t_L g1810 ( 
.A(n_1733),
.B(n_1538),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1705),
.A2(n_1459),
.B(n_1469),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1735),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1743),
.Y(n_1813)
);

INVxp33_ASAP7_75t_L g1814 ( 
.A(n_1734),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1684),
.Y(n_1815)
);

INVxp33_ASAP7_75t_L g1816 ( 
.A(n_1671),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1732),
.B(n_1611),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1682),
.A2(n_1700),
.B(n_1738),
.C(n_1694),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1743),
.B(n_1611),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1746),
.B(n_1611),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1703),
.A2(n_714),
.B1(n_715),
.B2(n_703),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1684),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1709),
.A2(n_1587),
.B(n_716),
.C(n_1393),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1746),
.B(n_1611),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1686),
.B(n_886),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1733),
.B(n_1611),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1676),
.Y(n_1827)
);

BUFx10_ASAP7_75t_L g1828 ( 
.A(n_1669),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1676),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1731),
.B(n_713),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1703),
.A2(n_1549),
.B1(n_1554),
.B2(n_713),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1684),
.B(n_1492),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1669),
.B(n_1504),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1671),
.B(n_1504),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1671),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1671),
.B(n_564),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1681),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1681),
.Y(n_1838)
);

O2A1O1Ixp5_ASAP7_75t_SL g1839 ( 
.A1(n_1722),
.A2(n_902),
.B(n_906),
.C(n_896),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1699),
.B(n_921),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_SL g1841 ( 
.A1(n_1687),
.A2(n_1446),
.B(n_870),
.C(n_861),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1726),
.B(n_631),
.Y(n_1842)
);

A2O1A1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1690),
.A2(n_1373),
.B(n_446),
.C(n_449),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1668),
.Y(n_1844)
);

INVx8_ASAP7_75t_L g1845 ( 
.A(n_1726),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1720),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1668),
.B(n_631),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1674),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1674),
.A2(n_1481),
.B1(n_590),
.B2(n_621),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1739),
.A2(n_1353),
.B(n_1481),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1726),
.B(n_634),
.Y(n_1851)
);

OA21x2_ASAP7_75t_L g1852 ( 
.A1(n_1721),
.A2(n_1284),
.B(n_1289),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1726),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1715),
.B(n_1),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1711),
.B(n_444),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1711),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1720),
.Y(n_1857)
);

OA21x2_ASAP7_75t_L g1858 ( 
.A1(n_1729),
.A2(n_1284),
.B(n_1297),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1715),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1729),
.A2(n_590),
.B1(n_621),
.B2(n_581),
.Y(n_1860)
);

O2A1O1Ixp5_ASAP7_75t_L g1861 ( 
.A1(n_1740),
.A2(n_1440),
.B(n_1431),
.C(n_1444),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1740),
.B(n_451),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1667),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1697),
.B(n_456),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_SL g1865 ( 
.A1(n_1697),
.A2(n_621),
.B1(n_640),
.B2(n_590),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1697),
.B(n_634),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1680),
.A2(n_470),
.B(n_472),
.C(n_466),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1672),
.B(n_662),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1671),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1665),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1678),
.B(n_474),
.Y(n_1871)
);

NOR2x2_ASAP7_75t_L g1872 ( 
.A(n_1684),
.B(n_662),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1704),
.Y(n_1873)
);

BUFx8_ASAP7_75t_L g1874 ( 
.A(n_1664),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1672),
.B(n_662),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1678),
.B(n_475),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1704),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1672),
.B(n_640),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1741),
.Y(n_1879)
);

NOR2xp67_ASAP7_75t_R g1880 ( 
.A(n_1717),
.B(n_1300),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1731),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1675),
.B(n_476),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1716),
.B(n_1172),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1678),
.B(n_478),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1704),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1704),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1678),
.B(n_479),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1704),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1741),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1672),
.B(n_3),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1704),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1741),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1672),
.B(n_3),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1675),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1672),
.B(n_4),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1704),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1678),
.B(n_1372),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1786),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1874),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1755),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1869),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1812),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1846),
.B(n_6),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1874),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1848),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1758),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1758),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1792),
.B(n_7),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1760),
.B(n_7),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1879),
.Y(n_1910)
);

AO31x2_ASAP7_75t_L g1911 ( 
.A1(n_1860),
.A2(n_1120),
.A3(n_1121),
.B(n_1118),
.Y(n_1911)
);

OAI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1784),
.A2(n_483),
.B1(n_485),
.B2(n_482),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1894),
.B(n_8),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1869),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1857),
.B(n_8),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1889),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1813),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1892),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1859),
.B(n_9),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1837),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1775),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1781),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1873),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1856),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1877),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1789),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1815),
.B(n_9),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1885),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1798),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1799),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1822),
.B(n_10),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1896),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1757),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1818),
.A2(n_490),
.B(n_487),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1770),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1886),
.Y(n_1936)
);

OA21x2_ASAP7_75t_L g1937 ( 
.A1(n_1864),
.A2(n_497),
.B(n_496),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1761),
.B(n_10),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1888),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1891),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1802),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1859),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1803),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1805),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1844),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1829),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1838),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1811),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_L g1949 ( 
.A1(n_1839),
.A2(n_1196),
.B(n_1182),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1782),
.A2(n_505),
.B(n_499),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1811),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1819),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1820),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1824),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1827),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1863),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1758),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1788),
.Y(n_1958)
);

OA21x2_ASAP7_75t_L g1959 ( 
.A1(n_1861),
.A2(n_508),
.B(n_506),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1788),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1806),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1806),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1796),
.B(n_11),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1858),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1858),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1835),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1852),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1795),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1808),
.Y(n_1969)
);

AO31x2_ASAP7_75t_L g1970 ( 
.A1(n_1849),
.A2(n_1137),
.A3(n_1129),
.B(n_1302),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1773),
.A2(n_514),
.B(n_513),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1756),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1756),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1825),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1852),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1783),
.B(n_11),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1800),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1825),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1817),
.B(n_14),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1800),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1759),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1759),
.Y(n_1982)
);

INVx4_ASAP7_75t_L g1983 ( 
.A(n_1759),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1883),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1855),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1785),
.Y(n_1986)
);

INVx3_ASAP7_75t_L g1987 ( 
.A(n_1883),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1785),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1862),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1794),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1750),
.B(n_1878),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1764),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1769),
.B(n_14),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1794),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1866),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1754),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1897),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1768),
.A2(n_1203),
.B(n_1198),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1749),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1779),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1804),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1897),
.B(n_15),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1751),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1766),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1854),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1840),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1826),
.B(n_17),
.Y(n_2007)
);

OAI221xp5_ASAP7_75t_L g2008 ( 
.A1(n_1847),
.A2(n_518),
.B1(n_523),
.B2(n_516),
.C(n_515),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1826),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1777),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1832),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1778),
.Y(n_2012)
);

NOR2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1870),
.B(n_526),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1816),
.B(n_18),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1845),
.Y(n_2015)
);

OAI21x1_ASAP7_75t_L g2016 ( 
.A1(n_1752),
.A2(n_1849),
.B(n_1850),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1810),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1832),
.Y(n_2018)
);

BUFx2_ASAP7_75t_L g2019 ( 
.A(n_1853),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1791),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1787),
.A2(n_1221),
.B(n_1213),
.Y(n_2021)
);

AOI22x1_ASAP7_75t_L g2022 ( 
.A1(n_1836),
.A2(n_529),
.B1(n_536),
.B2(n_528),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1771),
.A2(n_539),
.B1(n_544),
.B2(n_538),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1890),
.B(n_18),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1868),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1845),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1875),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1790),
.Y(n_2028)
);

AOI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1871),
.A2(n_1221),
.B(n_1213),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1893),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_1807),
.A2(n_566),
.B1(n_570),
.B2(n_557),
.C(n_550),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1895),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1842),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1851),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1865),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1865),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1845),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1828),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1828),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1780),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1767),
.B(n_20),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1833),
.B(n_20),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1872),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1834),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1876),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1765),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1884),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1887),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1880),
.Y(n_2049)
);

BUFx2_ASAP7_75t_SL g2050 ( 
.A(n_1831),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1841),
.A2(n_1211),
.B(n_1181),
.Y(n_2051)
);

BUFx3_ASAP7_75t_L g2052 ( 
.A(n_1793),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1831),
.A2(n_1228),
.B(n_1137),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1926),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1898),
.B(n_2044),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1954),
.B(n_1881),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1926),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1954),
.B(n_1814),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_2050),
.A2(n_1771),
.B1(n_1807),
.B2(n_1763),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1929),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1934),
.A2(n_1763),
.B1(n_1753),
.B2(n_1882),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1943),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1943),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1952),
.B(n_1772),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1929),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1905),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_1995),
.B(n_1797),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1930),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2010),
.B(n_1801),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1953),
.B(n_1830),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1930),
.Y(n_2071)
);

AO31x2_ASAP7_75t_L g2072 ( 
.A1(n_1964),
.A2(n_1867),
.A3(n_1774),
.B(n_1809),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2011),
.B(n_1809),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1906),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1941),
.Y(n_2075)
);

NOR2x1p5_ASAP7_75t_L g2076 ( 
.A(n_2043),
.B(n_1880),
.Y(n_2076)
);

BUFx2_ASAP7_75t_SL g2077 ( 
.A(n_1899),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1905),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1992),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2011),
.B(n_1821),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2018),
.B(n_1821),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1924),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1941),
.Y(n_2083)
);

OAI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_2043),
.A2(n_1823),
.B1(n_1843),
.B2(n_1753),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2018),
.B(n_21),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2045),
.B(n_1776),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1920),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1924),
.Y(n_2088)
);

INVx1_ASAP7_75t_SL g2089 ( 
.A(n_1945),
.Y(n_2089)
);

INVx5_ASAP7_75t_SL g2090 ( 
.A(n_1957),
.Y(n_2090)
);

NAND2x1p5_ASAP7_75t_L g2091 ( 
.A(n_1934),
.B(n_1762),
.Y(n_2091)
);

AND2x4_ASAP7_75t_SL g2092 ( 
.A(n_1992),
.B(n_897),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2009),
.B(n_21),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_1906),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1921),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_1900),
.B(n_22),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1910),
.B(n_24),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1922),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1902),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2009),
.B(n_24),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1902),
.Y(n_2101)
);

INVx3_ASAP7_75t_L g2102 ( 
.A(n_1992),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1923),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1925),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1917),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1916),
.B(n_25),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1992),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2035),
.A2(n_575),
.B1(n_576),
.B2(n_573),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1928),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1917),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1932),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1918),
.B(n_25),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1944),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_2039),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1933),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1944),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2045),
.B(n_26),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1948),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_1957),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2048),
.B(n_27),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_2039),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1948),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1935),
.Y(n_2123)
);

OR2x2_ASAP7_75t_L g2124 ( 
.A(n_1920),
.B(n_27),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1951),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1951),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_2005),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_1966),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_1997),
.B(n_28),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1958),
.B(n_29),
.Y(n_2130)
);

NAND2x1p5_ASAP7_75t_L g2131 ( 
.A(n_1934),
.B(n_1275),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_1956),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1936),
.Y(n_2133)
);

AND2x4_ASAP7_75t_SL g2134 ( 
.A(n_1957),
.B(n_897),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1899),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1960),
.B(n_30),
.Y(n_2136)
);

INVx4_ASAP7_75t_L g2137 ( 
.A(n_1957),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1939),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1904),
.Y(n_2139)
);

INVxp67_ASAP7_75t_L g2140 ( 
.A(n_2005),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1940),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1946),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1947),
.Y(n_2143)
);

AO31x2_ASAP7_75t_L g2144 ( 
.A1(n_1964),
.A2(n_1129),
.A3(n_32),
.B(n_30),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_1956),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1955),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_1997),
.B(n_31),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_2012),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2048),
.A2(n_2047),
.B1(n_1989),
.B2(n_1985),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1904),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2035),
.A2(n_580),
.B1(n_582),
.B2(n_577),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1961),
.B(n_32),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1962),
.B(n_33),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1982),
.B(n_33),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_1991),
.B(n_34),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1977),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1977),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1966),
.B(n_35),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2019),
.B(n_37),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2036),
.A2(n_584),
.B1(n_585),
.B2(n_583),
.Y(n_2160)
);

NOR2x1p5_ASAP7_75t_L g2161 ( 
.A(n_2052),
.B(n_586),
.Y(n_2161)
);

AOI21xp33_ASAP7_75t_L g2162 ( 
.A1(n_1937),
.A2(n_37),
.B(n_39),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1968),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1969),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1907),
.B(n_40),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2001),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1907),
.B(n_41),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1980),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2001),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2006),
.B(n_1972),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_1973),
.B(n_41),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1907),
.B(n_43),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1942),
.B(n_43),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1980),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1974),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1965),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1983),
.B(n_44),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_2012),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_1901),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1965),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1978),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1967),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_1983),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2017),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2017),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1983),
.B(n_45),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1901),
.Y(n_2187)
);

AO31x2_ASAP7_75t_L g2188 ( 
.A1(n_1967),
.A2(n_50),
.A3(n_47),
.B(n_49),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_1942),
.B(n_51),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1984),
.B(n_51),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1914),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1975),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2036),
.A2(n_588),
.B1(n_589),
.B2(n_587),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1999),
.B(n_2000),
.Y(n_2194)
);

AOI222xp33_ASAP7_75t_L g2195 ( 
.A1(n_2040),
.A2(n_593),
.B1(n_595),
.B2(n_604),
.C1(n_613),
.C2(n_614),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1914),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1975),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1984),
.B(n_53),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_SL g2199 ( 
.A1(n_1937),
.A2(n_617),
.B1(n_618),
.B2(n_615),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_2038),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2033),
.B(n_53),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2034),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1986),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1987),
.B(n_54),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_1903),
.Y(n_2205)
);

OR2x6_ASAP7_75t_L g2206 ( 
.A(n_2016),
.B(n_897),
.Y(n_2206)
);

INVxp67_ASAP7_75t_SL g2207 ( 
.A(n_1986),
.Y(n_2207)
);

OAI21xp33_ASAP7_75t_SL g2208 ( 
.A1(n_2049),
.A2(n_1981),
.B(n_1908),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1996),
.B(n_54),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1988),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2025),
.B(n_55),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2027),
.B(n_56),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1988),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2055),
.B(n_1987),
.Y(n_2214)
);

INVx5_ASAP7_75t_L g2215 ( 
.A(n_2206),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2066),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_2183),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2127),
.B(n_2030),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2088),
.B(n_2004),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2149),
.B(n_1937),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_2192),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2208),
.B(n_2046),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2058),
.B(n_2128),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2149),
.B(n_2003),
.Y(n_2224)
);

INVxp67_ASAP7_75t_SL g2225 ( 
.A(n_2192),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_2127),
.B(n_1942),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2140),
.B(n_2037),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2140),
.B(n_2037),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2066),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2056),
.B(n_2032),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2054),
.B(n_2028),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2176),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2148),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2079),
.B(n_2046),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2079),
.B(n_2020),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_SL g2236 ( 
.A1(n_2069),
.A2(n_1976),
.B1(n_2052),
.B2(n_2007),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2078),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2102),
.B(n_1903),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2102),
.B(n_1903),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2183),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_2094),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2107),
.B(n_1915),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_2135),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2166),
.B(n_2169),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2107),
.B(n_1915),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2078),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2057),
.B(n_1913),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2114),
.B(n_1915),
.Y(n_2248)
);

OR2x6_ASAP7_75t_L g2249 ( 
.A(n_2077),
.B(n_2016),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2082),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2148),
.B(n_2178),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2082),
.Y(n_2252)
);

NAND3xp33_ASAP7_75t_L g2253 ( 
.A(n_2059),
.B(n_1976),
.C(n_1950),
.Y(n_2253)
);

INVx2_ASAP7_75t_R g2254 ( 
.A(n_2197),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2060),
.B(n_1909),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2071),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_2137),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2086),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2133),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2178),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2062),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_2184),
.B(n_2002),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_2137),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2121),
.B(n_2064),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2133),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2095),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2205),
.B(n_1927),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2098),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2205),
.B(n_1931),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2175),
.B(n_1990),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2200),
.B(n_1938),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2181),
.B(n_1990),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2062),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2103),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2185),
.B(n_2015),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2176),
.Y(n_2276)
);

INVx1_ASAP7_75t_SL g2277 ( 
.A(n_2087),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_2119),
.B(n_2015),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2104),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_2132),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2109),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2111),
.Y(n_2282)
);

BUFx3_ASAP7_75t_L g2283 ( 
.A(n_2094),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2132),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2080),
.B(n_1963),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2115),
.Y(n_2286)
);

AO21x2_ASAP7_75t_L g2287 ( 
.A1(n_2207),
.A2(n_1912),
.B(n_1994),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2081),
.B(n_1979),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_2146),
.B(n_2024),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2187),
.B(n_2073),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2187),
.B(n_2026),
.Y(n_2291)
);

INVx5_ASAP7_75t_L g2292 ( 
.A(n_2206),
.Y(n_2292)
);

BUFx2_ASAP7_75t_SL g2293 ( 
.A(n_2135),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2087),
.B(n_2026),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_2139),
.Y(n_2295)
);

INVxp67_ASAP7_75t_SL g2296 ( 
.A(n_2207),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2063),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2123),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2063),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_SL g2300 ( 
.A(n_2162),
.B(n_1912),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2138),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2141),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_2139),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2179),
.B(n_1993),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2099),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2179),
.B(n_2041),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2202),
.B(n_2007),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2074),
.B(n_2007),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2074),
.B(n_1919),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2065),
.B(n_1911),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2191),
.B(n_1919),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2145),
.Y(n_2312)
);

BUFx2_ASAP7_75t_L g2313 ( 
.A(n_2150),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2142),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2142),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2143),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2196),
.B(n_1919),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2143),
.B(n_2042),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_2150),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2065),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2068),
.B(n_1911),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2068),
.B(n_1911),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2070),
.B(n_2014),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2163),
.B(n_2053),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2099),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2145),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2101),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2101),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2170),
.B(n_1970),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2180),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2075),
.B(n_1911),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2164),
.B(n_1970),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2075),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2083),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2083),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2124),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2113),
.B(n_2013),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_SL g2338 ( 
.A1(n_2069),
.A2(n_2021),
.B1(n_1959),
.B2(n_2008),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2313),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2286),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2298),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2258),
.B(n_2194),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_2295),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2301),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2217),
.B(n_2076),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2251),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2302),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2266),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2336),
.B(n_2067),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2290),
.Y(n_2350)
);

BUFx3_ASAP7_75t_L g2351 ( 
.A(n_2283),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2280),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2268),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2258),
.B(n_2118),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2217),
.B(n_2173),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2223),
.B(n_2090),
.Y(n_2356)
);

NOR2xp67_ASAP7_75t_L g2357 ( 
.A(n_2222),
.B(n_2113),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2224),
.B(n_2118),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2264),
.B(n_2090),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2274),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2238),
.B(n_2090),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2240),
.B(n_2173),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2279),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2281),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2239),
.B(n_2155),
.Y(n_2365)
);

NOR2xp67_ASAP7_75t_L g2366 ( 
.A(n_2222),
.B(n_2116),
.Y(n_2366)
);

BUFx3_ASAP7_75t_L g2367 ( 
.A(n_2283),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_2280),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2242),
.B(n_2116),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2282),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_2295),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2219),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2224),
.B(n_2122),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2219),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2234),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2220),
.B(n_2122),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2251),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2257),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2257),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2218),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2245),
.B(n_2106),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2309),
.B(n_2248),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2293),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2284),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2231),
.Y(n_2385)
);

AOI222xp33_ASAP7_75t_L g2386 ( 
.A1(n_2253),
.A2(n_2059),
.B1(n_2061),
.B2(n_2084),
.C1(n_2159),
.C2(n_2161),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2308),
.B(n_2112),
.Y(n_2387)
);

OAI21xp5_ASAP7_75t_SL g2388 ( 
.A1(n_2253),
.A2(n_2061),
.B(n_2199),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2285),
.B(n_2105),
.Y(n_2389)
);

INVx1_ASAP7_75t_SL g2390 ( 
.A(n_2277),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2231),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2263),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2241),
.B(n_2209),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2336),
.B(n_2129),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_2295),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2284),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2263),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2319),
.B(n_2117),
.Y(n_2398)
);

INVx5_ASAP7_75t_L g2399 ( 
.A(n_2249),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2220),
.B(n_2125),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2288),
.B(n_2105),
.Y(n_2401)
);

OR2x2_ASAP7_75t_L g2402 ( 
.A(n_2262),
.B(n_2147),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2247),
.B(n_2096),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2226),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2312),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2312),
.Y(n_2406)
);

INVxp67_ASAP7_75t_SL g2407 ( 
.A(n_2221),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2326),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2226),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2247),
.B(n_2097),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2240),
.B(n_2173),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2326),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2221),
.Y(n_2413)
);

INVx5_ASAP7_75t_L g2414 ( 
.A(n_2249),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2306),
.B(n_2110),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2256),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2227),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2311),
.B(n_2110),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2216),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2229),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2227),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2237),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2225),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2317),
.B(n_2085),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2319),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2228),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2246),
.B(n_2125),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2250),
.Y(n_2428)
);

BUFx2_ASAP7_75t_SL g2429 ( 
.A(n_2243),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2228),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2252),
.B(n_2126),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2320),
.B(n_2126),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2275),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2259),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2265),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2214),
.B(n_2089),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2333),
.B(n_2156),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2275),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2300),
.A2(n_2199),
.B1(n_2195),
.B2(n_2108),
.Y(n_2439)
);

AOI222xp33_ASAP7_75t_L g2440 ( 
.A1(n_2300),
.A2(n_2120),
.B1(n_2031),
.B2(n_2193),
.C1(n_2151),
.C2(n_2160),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2314),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2337),
.B(n_2093),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2319),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2334),
.B(n_2156),
.Y(n_2444)
);

NAND2x1p5_ASAP7_75t_L g2445 ( 
.A(n_2277),
.B(n_2189),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2315),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2335),
.B(n_2157),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2316),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2255),
.B(n_2171),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_L g2450 ( 
.A1(n_2338),
.A2(n_2131),
.B1(n_1971),
.B2(n_2091),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_2303),
.B(n_2189),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2352),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2383),
.B(n_2233),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2386),
.A2(n_2338),
.B1(n_2287),
.B2(n_2236),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2342),
.B(n_2225),
.Y(n_2455)
);

AOI21xp33_ASAP7_75t_L g2456 ( 
.A1(n_2388),
.A2(n_2287),
.B(n_2236),
.Y(n_2456)
);

OAI21x1_ASAP7_75t_L g2457 ( 
.A1(n_2346),
.A2(n_2296),
.B(n_2276),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2383),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2352),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2388),
.B(n_2023),
.C(n_2249),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2368),
.Y(n_2461)
);

OAI211xp5_ASAP7_75t_L g2462 ( 
.A1(n_2386),
.A2(n_2296),
.B(n_2165),
.C(n_2172),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2368),
.Y(n_2463)
);

OAI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2439),
.A2(n_2131),
.B1(n_2212),
.B2(n_2211),
.C(n_2091),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2346),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2439),
.A2(n_2450),
.B1(n_2440),
.B2(n_2350),
.Y(n_2466)
);

AOI222xp33_ASAP7_75t_L g2467 ( 
.A1(n_2393),
.A2(n_2154),
.B1(n_2186),
.B2(n_2177),
.C1(n_2167),
.C2(n_2255),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2429),
.B(n_2235),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2384),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2382),
.B(n_2291),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2351),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2367),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2349),
.B(n_2449),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2384),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2445),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2445),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2371),
.Y(n_2477)
);

OAI31xp33_ASAP7_75t_L g2478 ( 
.A1(n_2450),
.A2(n_2189),
.A3(n_2269),
.B(n_2267),
.Y(n_2478)
);

INVxp67_ASAP7_75t_SL g2479 ( 
.A(n_2423),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2345),
.B(n_2323),
.Y(n_2480)
);

INVxp67_ASAP7_75t_SL g2481 ( 
.A(n_2423),
.Y(n_2481)
);

OAI221xp5_ASAP7_75t_L g2482 ( 
.A1(n_2440),
.A2(n_2201),
.B1(n_2206),
.B2(n_2289),
.C(n_2022),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_2339),
.B(n_2260),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2345),
.B(n_2278),
.Y(n_2484)
);

OAI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2393),
.A2(n_2292),
.B1(n_2215),
.B2(n_2158),
.C(n_2198),
.Y(n_2485)
);

OA21x2_ASAP7_75t_L g2486 ( 
.A1(n_2407),
.A2(n_2276),
.B(n_2232),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2407),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2340),
.Y(n_2488)
);

INVx1_ASAP7_75t_SL g2489 ( 
.A(n_2390),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2342),
.B(n_2270),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2341),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2344),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2361),
.B(n_2294),
.Y(n_2493)
);

INVxp67_ASAP7_75t_SL g2494 ( 
.A(n_2357),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2355),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_2425),
.Y(n_2496)
);

AOI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_2376),
.A2(n_2292),
.B(n_2215),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2395),
.B(n_2307),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2390),
.Y(n_2499)
);

AND4x1_ASAP7_75t_L g2500 ( 
.A(n_2398),
.B(n_2204),
.C(n_2190),
.D(n_2100),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2347),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2355),
.B(n_2278),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2396),
.Y(n_2503)
);

OAI21x1_ASAP7_75t_L g2504 ( 
.A1(n_2378),
.A2(n_2330),
.B(n_2232),
.Y(n_2504)
);

AO21x2_ASAP7_75t_L g2505 ( 
.A1(n_2366),
.A2(n_2254),
.B(n_2310),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2362),
.Y(n_2506)
);

INVxp33_ASAP7_75t_L g2507 ( 
.A(n_2436),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2362),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2348),
.Y(n_2509)
);

INVx2_ASAP7_75t_SL g2510 ( 
.A(n_2411),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_2404),
.A2(n_2254),
.B1(n_2292),
.B2(n_2215),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2411),
.Y(n_2512)
);

OAI33xp33_ASAP7_75t_L g2513 ( 
.A1(n_2405),
.A2(n_2310),
.A3(n_2331),
.B1(n_2321),
.B2(n_2322),
.B3(n_2329),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2353),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2398),
.A2(n_2318),
.B1(n_2324),
.B2(n_2304),
.Y(n_2515)
);

OAI33xp33_ASAP7_75t_L g2516 ( 
.A1(n_2406),
.A2(n_2331),
.A3(n_2321),
.B1(n_2322),
.B2(n_2270),
.B3(n_2272),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2360),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2451),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2359),
.B(n_2271),
.Y(n_2519)
);

HB1xp67_ASAP7_75t_L g2520 ( 
.A(n_2408),
.Y(n_2520)
);

AOI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2409),
.A2(n_2324),
.B1(n_2230),
.B2(n_2292),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2451),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2363),
.Y(n_2523)
);

OAI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2399),
.A2(n_2215),
.B1(n_2244),
.B2(n_2332),
.Y(n_2524)
);

AOI221xp5_ASAP7_75t_L g2525 ( 
.A1(n_2376),
.A2(n_2152),
.B1(n_2153),
.B2(n_2136),
.C(n_2130),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2364),
.Y(n_2526)
);

OAI21xp5_ASAP7_75t_SL g2527 ( 
.A1(n_2442),
.A2(n_2092),
.B(n_2134),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2370),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2403),
.B(n_2272),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_2400),
.B(n_2330),
.C(n_2327),
.Y(n_2530)
);

BUFx3_ASAP7_75t_L g2531 ( 
.A(n_2443),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2372),
.B(n_2374),
.Y(n_2532)
);

AOI22xp33_ASAP7_75t_L g2533 ( 
.A1(n_2375),
.A2(n_2053),
.B1(n_2305),
.B2(n_2328),
.Y(n_2533)
);

HB1xp67_ASAP7_75t_L g2534 ( 
.A(n_2412),
.Y(n_2534)
);

INVx1_ASAP7_75t_SL g2535 ( 
.A(n_2343),
.Y(n_2535)
);

INVx1_ASAP7_75t_SL g2536 ( 
.A(n_2394),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2387),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2416),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2413),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2499),
.Y(n_2540)
);

NOR2xp67_ASAP7_75t_L g2541 ( 
.A(n_2485),
.B(n_2399),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2461),
.Y(n_2542)
);

INVx3_ASAP7_75t_L g2543 ( 
.A(n_2472),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2474),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2479),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2481),
.Y(n_2546)
);

NAND2x1_ASAP7_75t_L g2547 ( 
.A(n_2484),
.B(n_2377),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2489),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_2458),
.Y(n_2549)
);

HB1xp67_ASAP7_75t_L g2550 ( 
.A(n_2489),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2484),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2508),
.B(n_2379),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2536),
.B(n_2380),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2536),
.B(n_2385),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2468),
.B(n_2433),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2452),
.B(n_2391),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2502),
.Y(n_2557)
);

INVx1_ASAP7_75t_SL g2558 ( 
.A(n_2477),
.Y(n_2558)
);

OR2x2_ASAP7_75t_L g2559 ( 
.A(n_2473),
.B(n_2410),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2487),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2496),
.B(n_2402),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2471),
.B(n_2498),
.Y(n_2562)
);

NAND2x1_ASAP7_75t_L g2563 ( 
.A(n_2502),
.B(n_2438),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2519),
.B(n_2356),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2459),
.B(n_2419),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2455),
.B(n_2420),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2463),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2469),
.B(n_2422),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2537),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2455),
.B(n_2428),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2510),
.B(n_2392),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2503),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2520),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2534),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2493),
.B(n_2417),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2470),
.B(n_2421),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2506),
.B(n_2426),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2506),
.B(n_2430),
.Y(n_2578)
);

INVx4_ASAP7_75t_L g2579 ( 
.A(n_2531),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2507),
.B(n_2397),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2518),
.B(n_2365),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2462),
.B(n_2381),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2466),
.B(n_2358),
.Y(n_2583)
);

NAND2x1_ASAP7_75t_L g2584 ( 
.A(n_2453),
.B(n_2434),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2488),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2495),
.B(n_2399),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2512),
.B(n_2399),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2453),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2491),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2462),
.B(n_2358),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2529),
.B(n_2373),
.Y(n_2591)
);

OR2x2_ASAP7_75t_L g2592 ( 
.A(n_2535),
.B(n_2373),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2522),
.B(n_2414),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2535),
.B(n_2389),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2465),
.B(n_2401),
.Y(n_2595)
);

AND2x4_ASAP7_75t_SL g2596 ( 
.A(n_2483),
.B(n_2424),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2475),
.B(n_2418),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2490),
.B(n_2354),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2490),
.B(n_2354),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2480),
.B(n_2414),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2492),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2501),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_2476),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2483),
.B(n_2369),
.Y(n_2604)
);

OR2x2_ASAP7_75t_L g2605 ( 
.A(n_2539),
.B(n_2400),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2515),
.B(n_2494),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2500),
.B(n_2415),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2454),
.B(n_2435),
.Y(n_2608)
);

INVx1_ASAP7_75t_SL g2609 ( 
.A(n_2497),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2457),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2521),
.B(n_2441),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2509),
.B(n_2446),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2467),
.B(n_2448),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2532),
.B(n_2427),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2467),
.B(n_2414),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2514),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2478),
.B(n_2414),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2527),
.B(n_2427),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2486),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2511),
.B(n_2517),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2523),
.B(n_2431),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2548),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2548),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2579),
.Y(n_2624)
);

OR2x2_ASAP7_75t_L g2625 ( 
.A(n_2550),
.B(n_2573),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2579),
.Y(n_2626)
);

NAND2x1_ASAP7_75t_L g2627 ( 
.A(n_2600),
.B(n_2486),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2550),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2619),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2543),
.B(n_2456),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2619),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2573),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2540),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2540),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2558),
.B(n_2456),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2543),
.B(n_2526),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2558),
.B(n_2600),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2545),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2549),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2546),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2561),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2553),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2542),
.Y(n_2643)
);

BUFx2_ASAP7_75t_L g2644 ( 
.A(n_2588),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2582),
.B(n_2460),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2547),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2544),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2572),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2582),
.B(n_2528),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2574),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2560),
.Y(n_2651)
);

BUFx2_ASAP7_75t_L g2652 ( 
.A(n_2552),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2592),
.B(n_2532),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2564),
.B(n_2538),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2607),
.B(n_2525),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2596),
.B(n_2497),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2594),
.B(n_2504),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2580),
.B(n_2525),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2577),
.B(n_2482),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2565),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2565),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2551),
.B(n_2505),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2606),
.B(n_2505),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2568),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2604),
.B(n_2524),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2568),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2555),
.B(n_2557),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2617),
.B(n_2524),
.Y(n_2668)
);

AND2x4_ASAP7_75t_L g2669 ( 
.A(n_2552),
.B(n_2530),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2578),
.B(n_2533),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2603),
.B(n_2431),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2567),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2603),
.B(n_2432),
.Y(n_2673)
);

NOR2x1_ASAP7_75t_L g2674 ( 
.A(n_2609),
.B(n_2485),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2612),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2584),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2612),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2621),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2559),
.B(n_2590),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2569),
.B(n_2482),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2581),
.B(n_2432),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2609),
.B(n_2541),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2563),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2652),
.B(n_2571),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2667),
.B(n_2575),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2623),
.B(n_2583),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2629),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2646),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2625),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2625),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_L g2691 ( 
.A(n_2674),
.B(n_2583),
.C(n_2590),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_R g2692 ( 
.A(n_2622),
.B(n_2562),
.Y(n_2692)
);

HB1xp67_ASAP7_75t_L g2693 ( 
.A(n_2629),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2631),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2631),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2667),
.B(n_2571),
.Y(n_2696)
);

AOI21xp33_ASAP7_75t_L g2697 ( 
.A1(n_2635),
.A2(n_2608),
.B(n_2615),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2637),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2641),
.B(n_2613),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2628),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2637),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_SL g2702 ( 
.A1(n_2645),
.A2(n_2464),
.B1(n_2608),
.B2(n_2554),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2679),
.B(n_2554),
.Y(n_2703)
);

INVx1_ASAP7_75t_SL g2704 ( 
.A(n_2637),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2665),
.B(n_2576),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2682),
.A2(n_2620),
.B(n_2464),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2679),
.B(n_2566),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2642),
.B(n_2570),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2683),
.Y(n_2709)
);

AOI22x1_ASAP7_75t_L g2710 ( 
.A1(n_2663),
.A2(n_2593),
.B1(n_2586),
.B2(n_2587),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2644),
.B(n_2598),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2665),
.B(n_2618),
.Y(n_2712)
);

INVxp67_ASAP7_75t_L g2713 ( 
.A(n_2644),
.Y(n_2713)
);

AOI211xp5_ASAP7_75t_L g2714 ( 
.A1(n_2655),
.A2(n_2611),
.B(n_2593),
.C(n_2586),
.Y(n_2714)
);

CKINVDCx16_ASAP7_75t_R g2715 ( 
.A(n_2639),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2668),
.B(n_2595),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2683),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_R g2718 ( 
.A(n_2633),
.B(n_2585),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2624),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2632),
.Y(n_2720)
);

NAND3xp33_ASAP7_75t_SL g2721 ( 
.A(n_2630),
.B(n_2610),
.C(n_2556),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2668),
.B(n_2597),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2634),
.Y(n_2723)
);

OR2x6_ASAP7_75t_L g2724 ( 
.A(n_2624),
.B(n_2587),
.Y(n_2724)
);

NAND4xp25_ASAP7_75t_L g2725 ( 
.A(n_2680),
.B(n_2556),
.C(n_2601),
.D(n_2589),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2649),
.B(n_2599),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2627),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2656),
.B(n_2591),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2656),
.B(n_2602),
.Y(n_2729)
);

INVxp67_ASAP7_75t_L g2730 ( 
.A(n_2626),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2704),
.B(n_2658),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2705),
.B(n_2626),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2687),
.Y(n_2733)
);

INVx2_ASAP7_75t_SL g2734 ( 
.A(n_2684),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2687),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2713),
.B(n_2636),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2715),
.B(n_2638),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2696),
.B(n_2654),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2693),
.Y(n_2739)
);

BUFx12f_ASAP7_75t_L g2740 ( 
.A(n_2719),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2693),
.Y(n_2741)
);

NAND2x1p5_ASAP7_75t_L g2742 ( 
.A(n_2688),
.B(n_2636),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2684),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_2691),
.B(n_2640),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2698),
.Y(n_2745)
);

INVxp67_ASAP7_75t_L g2746 ( 
.A(n_2727),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2713),
.Y(n_2747)
);

INVxp33_ASAP7_75t_L g2748 ( 
.A(n_2692),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2722),
.B(n_2716),
.Y(n_2749)
);

HB1xp67_ASAP7_75t_L g2750 ( 
.A(n_2727),
.Y(n_2750)
);

OR2x2_ASAP7_75t_L g2751 ( 
.A(n_2701),
.B(n_2653),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2689),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2724),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2685),
.B(n_2654),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2690),
.B(n_2630),
.Y(n_2755)
);

INVxp67_ASAP7_75t_L g2756 ( 
.A(n_2724),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2711),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2724),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2694),
.Y(n_2759)
);

NAND3xp33_ASAP7_75t_L g2760 ( 
.A(n_2686),
.B(n_2659),
.C(n_2663),
.Y(n_2760)
);

OR2x4_ASAP7_75t_L g2761 ( 
.A(n_2723),
.B(n_2648),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2712),
.B(n_2678),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2695),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2709),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2730),
.B(n_2699),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2710),
.Y(n_2766)
);

OR2x6_ASAP7_75t_L g2767 ( 
.A(n_2730),
.B(n_2643),
.Y(n_2767)
);

OR2x6_ASAP7_75t_L g2768 ( 
.A(n_2686),
.B(n_2699),
.Y(n_2768)
);

NOR2x1_ASAP7_75t_L g2769 ( 
.A(n_2768),
.B(n_2767),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2760),
.A2(n_2702),
.B1(n_2706),
.B2(n_2714),
.Y(n_2770)
);

AOI222xp33_ASAP7_75t_L g2771 ( 
.A1(n_2760),
.A2(n_2706),
.B1(n_2721),
.B2(n_2744),
.C1(n_2737),
.C2(n_2755),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2740),
.A2(n_2721),
.B1(n_2728),
.B2(n_2697),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2734),
.B(n_2729),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2750),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2743),
.A2(n_2697),
.B1(n_2669),
.B2(n_2670),
.Y(n_2775)
);

OAI221xp5_ASAP7_75t_SL g2776 ( 
.A1(n_2768),
.A2(n_2703),
.B1(n_2726),
.B2(n_2707),
.C(n_2725),
.Y(n_2776)
);

INVxp67_ASAP7_75t_SL g2777 ( 
.A(n_2742),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2733),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2735),
.Y(n_2779)
);

NOR3xp33_ASAP7_75t_L g2780 ( 
.A(n_2766),
.B(n_2700),
.C(n_2720),
.Y(n_2780)
);

OAI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2768),
.A2(n_2676),
.B1(n_2708),
.B2(n_2653),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2739),
.Y(n_2782)
);

OAI21xp33_ASAP7_75t_L g2783 ( 
.A1(n_2748),
.A2(n_2718),
.B(n_2670),
.Y(n_2783)
);

AOI322xp5_ASAP7_75t_L g2784 ( 
.A1(n_2755),
.A2(n_2647),
.A3(n_2650),
.B1(n_2661),
.B2(n_2666),
.C1(n_2664),
.C2(n_2660),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2741),
.Y(n_2785)
);

OA21x2_ASAP7_75t_L g2786 ( 
.A1(n_2746),
.A2(n_2717),
.B(n_2676),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2742),
.Y(n_2787)
);

AOI21xp33_ASAP7_75t_SL g2788 ( 
.A1(n_2757),
.A2(n_2731),
.B(n_2751),
.Y(n_2788)
);

AND2x4_ASAP7_75t_L g2789 ( 
.A(n_2756),
.B(n_2738),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2736),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2749),
.B(n_2669),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2736),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2767),
.Y(n_2793)
);

OAI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2756),
.A2(n_2669),
.B1(n_2681),
.B2(n_2614),
.Y(n_2794)
);

AOI211xp5_ASAP7_75t_L g2795 ( 
.A1(n_2732),
.A2(n_2672),
.B(n_2651),
.C(n_2675),
.Y(n_2795)
);

OAI21xp33_ASAP7_75t_L g2796 ( 
.A1(n_2754),
.A2(n_2681),
.B(n_2657),
.Y(n_2796)
);

INVx2_ASAP7_75t_SL g2797 ( 
.A(n_2767),
.Y(n_2797)
);

AND3x1_ASAP7_75t_L g2798 ( 
.A(n_2753),
.B(n_2677),
.C(n_2671),
.Y(n_2798)
);

HB1xp67_ASAP7_75t_L g2799 ( 
.A(n_2746),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2762),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2772),
.B(n_2765),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_2777),
.B(n_2765),
.Y(n_2802)
);

NAND4xp25_ASAP7_75t_L g2803 ( 
.A(n_2771),
.B(n_2758),
.C(n_2745),
.D(n_2747),
.Y(n_2803)
);

INVxp67_ASAP7_75t_SL g2804 ( 
.A(n_2769),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2786),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2789),
.B(n_2764),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2783),
.B(n_2761),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2786),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2789),
.B(n_2764),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2787),
.B(n_2752),
.Y(n_2810)
);

OAI21xp5_ASAP7_75t_SL g2811 ( 
.A1(n_2770),
.A2(n_2763),
.B(n_2759),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2799),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2797),
.B(n_2761),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2800),
.B(n_2657),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2775),
.B(n_2671),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2773),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2774),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2781),
.B(n_2673),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2776),
.A2(n_2662),
.B(n_2616),
.Y(n_2819)
);

INVx1_ASAP7_75t_SL g2820 ( 
.A(n_2791),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2793),
.Y(n_2821)
);

INVxp33_ASAP7_75t_L g2822 ( 
.A(n_2788),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2794),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2796),
.B(n_2673),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2778),
.Y(n_2825)
);

HB1xp67_ASAP7_75t_L g2826 ( 
.A(n_2808),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2802),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2805),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2806),
.B(n_2790),
.Y(n_2829)
);

XOR2x2_ASAP7_75t_L g2830 ( 
.A(n_2818),
.B(n_2798),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2809),
.Y(n_2831)
);

NAND2xp33_ASAP7_75t_L g2832 ( 
.A(n_2823),
.B(n_2780),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2814),
.B(n_2792),
.Y(n_2833)
);

OAI21xp33_ASAP7_75t_L g2834 ( 
.A1(n_2822),
.A2(n_2784),
.B(n_2782),
.Y(n_2834)
);

HB1xp67_ASAP7_75t_L g2835 ( 
.A(n_2804),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_SL g2836 ( 
.A(n_2803),
.B(n_2785),
.C(n_2779),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2813),
.Y(n_2837)
);

INVx1_ASAP7_75t_SL g2838 ( 
.A(n_2820),
.Y(n_2838)
);

NOR2x1_ASAP7_75t_L g2839 ( 
.A(n_2813),
.B(n_2662),
.Y(n_2839)
);

AOI221xp5_ASAP7_75t_SL g2840 ( 
.A1(n_2819),
.A2(n_2795),
.B1(n_2605),
.B2(n_2516),
.C(n_2513),
.Y(n_2840)
);

INVx1_ASAP7_75t_SL g2841 ( 
.A(n_2810),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2824),
.B(n_2437),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2812),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2821),
.B(n_2437),
.Y(n_2844)
);

OAI211xp5_ASAP7_75t_L g2845 ( 
.A1(n_2834),
.A2(n_2811),
.B(n_2801),
.C(n_2815),
.Y(n_2845)
);

NAND2xp33_ASAP7_75t_L g2846 ( 
.A(n_2835),
.B(n_2815),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2838),
.A2(n_2807),
.B1(n_2816),
.B2(n_2817),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2827),
.B(n_2825),
.Y(n_2848)
);

INVx2_ASAP7_75t_SL g2849 ( 
.A(n_2841),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2826),
.Y(n_2850)
);

AOI21xp33_ASAP7_75t_L g2851 ( 
.A1(n_2837),
.A2(n_56),
.B(n_58),
.Y(n_2851)
);

NOR3xp33_ASAP7_75t_L g2852 ( 
.A(n_2832),
.B(n_2447),
.C(n_2444),
.Y(n_2852)
);

NAND3xp33_ASAP7_75t_L g2853 ( 
.A(n_2836),
.B(n_2447),
.C(n_2444),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2843),
.B(n_59),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2829),
.B(n_65),
.Y(n_2855)
);

NAND3xp33_ASAP7_75t_L g2856 ( 
.A(n_2839),
.B(n_620),
.C(n_619),
.Y(n_2856)
);

NOR3xp33_ASAP7_75t_L g2857 ( 
.A(n_2831),
.B(n_628),
.C(n_627),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2849),
.B(n_2833),
.Y(n_2858)
);

NAND4xp25_ASAP7_75t_L g2859 ( 
.A(n_2847),
.B(n_2842),
.C(n_2844),
.D(n_2828),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2850),
.B(n_2840),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_SL g2861 ( 
.A(n_2848),
.B(n_2830),
.Y(n_2861)
);

NAND2xp33_ASAP7_75t_L g2862 ( 
.A(n_2852),
.B(n_2853),
.Y(n_2862)
);

NOR2x1_ASAP7_75t_L g2863 ( 
.A(n_2845),
.B(n_2840),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2846),
.Y(n_2864)
);

NOR3xp33_ASAP7_75t_L g2865 ( 
.A(n_2855),
.B(n_639),
.C(n_635),
.Y(n_2865)
);

NOR2xp67_ASAP7_75t_L g2866 ( 
.A(n_2856),
.B(n_65),
.Y(n_2866)
);

NOR2x1_ASAP7_75t_L g2867 ( 
.A(n_2854),
.B(n_2851),
.Y(n_2867)
);

AOI311xp33_ASAP7_75t_L g2868 ( 
.A1(n_2857),
.A2(n_2188),
.A3(n_67),
.B(n_68),
.C(n_69),
.Y(n_2868)
);

NAND4xp25_ASAP7_75t_SL g2869 ( 
.A(n_2845),
.B(n_2273),
.C(n_2297),
.D(n_2261),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2846),
.Y(n_2870)
);

AOI221x1_ASAP7_75t_L g2871 ( 
.A1(n_2859),
.A2(n_2870),
.B1(n_2864),
.B2(n_2865),
.C(n_2863),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2867),
.B(n_2866),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2858),
.B(n_2299),
.Y(n_2873)
);

AOI222xp33_ASAP7_75t_L g2874 ( 
.A1(n_2860),
.A2(n_2092),
.B1(n_2134),
.B2(n_2188),
.C1(n_2325),
.C2(n_71),
.Y(n_2874)
);

NOR2x1_ASAP7_75t_L g2875 ( 
.A(n_2862),
.B(n_66),
.Y(n_2875)
);

AOI22xp33_ASAP7_75t_L g2876 ( 
.A1(n_2861),
.A2(n_2203),
.B1(n_2213),
.B2(n_2210),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2868),
.B(n_2325),
.Y(n_2877)
);

NAND5xp2_ASAP7_75t_L g2878 ( 
.A(n_2869),
.B(n_66),
.C(n_68),
.D(n_69),
.E(n_70),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2864),
.B(n_2188),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2870),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2864),
.B(n_2188),
.Y(n_2881)
);

NOR2x1_ASAP7_75t_L g2882 ( 
.A(n_2859),
.B(n_73),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2870),
.Y(n_2883)
);

INVx1_ASAP7_75t_SL g2884 ( 
.A(n_2870),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2864),
.B(n_2144),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2864),
.B(n_74),
.Y(n_2886)
);

NAND4xp75_ASAP7_75t_L g2887 ( 
.A(n_2863),
.B(n_78),
.C(n_75),
.D(n_76),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2884),
.B(n_75),
.Y(n_2888)
);

A2O1A1Ixp33_ASAP7_75t_L g2889 ( 
.A1(n_2880),
.A2(n_82),
.B(n_76),
.C(n_81),
.Y(n_2889)
);

AO22x2_ASAP7_75t_SL g2890 ( 
.A1(n_2883),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2890)
);

NOR2x1_ASAP7_75t_L g2891 ( 
.A(n_2887),
.B(n_85),
.Y(n_2891)
);

AOI31xp33_ASAP7_75t_L g2892 ( 
.A1(n_2875),
.A2(n_643),
.A3(n_648),
.B(n_641),
.Y(n_2892)
);

NOR3xp33_ASAP7_75t_L g2893 ( 
.A(n_2886),
.B(n_657),
.C(n_653),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2882),
.Y(n_2894)
);

NOR3xp33_ASAP7_75t_L g2895 ( 
.A(n_2872),
.B(n_668),
.C(n_661),
.Y(n_2895)
);

INVx1_ASAP7_75t_SL g2896 ( 
.A(n_2873),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2879),
.B(n_2877),
.Y(n_2897)
);

NOR3xp33_ASAP7_75t_L g2898 ( 
.A(n_2878),
.B(n_671),
.C(n_669),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2871),
.B(n_85),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2881),
.B(n_2180),
.Y(n_2900)
);

NAND4xp75_ASAP7_75t_L g2901 ( 
.A(n_2874),
.B(n_92),
.C(n_87),
.D(n_88),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2876),
.A2(n_2885),
.B1(n_2168),
.B2(n_2174),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2896),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2890),
.B(n_2885),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2894),
.B(n_679),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2888),
.Y(n_2906)
);

NAND4xp25_ASAP7_75t_L g2907 ( 
.A(n_2891),
.B(n_96),
.C(n_88),
.D(n_93),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2901),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2899),
.Y(n_2909)
);

OAI211xp5_ASAP7_75t_SL g2910 ( 
.A1(n_2897),
.A2(n_97),
.B(n_93),
.C(n_96),
.Y(n_2910)
);

NAND2x1p5_ASAP7_75t_L g2911 ( 
.A(n_2900),
.B(n_97),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2892),
.Y(n_2912)
);

OR3x1_ASAP7_75t_L g2913 ( 
.A(n_2898),
.B(n_99),
.C(n_100),
.Y(n_2913)
);

NOR3xp33_ASAP7_75t_L g2914 ( 
.A(n_2893),
.B(n_2895),
.C(n_2889),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2911),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2913),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2904),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2903),
.Y(n_2918)
);

NOR2x1_ASAP7_75t_L g2919 ( 
.A(n_2907),
.B(n_101),
.Y(n_2919)
);

NAND2x1_ASAP7_75t_L g2920 ( 
.A(n_2908),
.B(n_2902),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2910),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2909),
.Y(n_2922)
);

INVxp67_ASAP7_75t_L g2923 ( 
.A(n_2906),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2912),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2905),
.Y(n_2925)
);

XNOR2xp5_ASAP7_75t_L g2926 ( 
.A(n_2918),
.B(n_2914),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2915),
.Y(n_2927)
);

XNOR2x1_ASAP7_75t_L g2928 ( 
.A(n_2919),
.B(n_102),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2917),
.B(n_102),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2916),
.Y(n_2930)
);

NOR2x1_ASAP7_75t_L g2931 ( 
.A(n_2920),
.B(n_103),
.Y(n_2931)
);

OAI22x1_ASAP7_75t_L g2932 ( 
.A1(n_2921),
.A2(n_681),
.B1(n_682),
.B2(n_691),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2922),
.Y(n_2933)
);

HB1xp67_ASAP7_75t_L g2934 ( 
.A(n_2924),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2923),
.Y(n_2935)
);

AOI211xp5_ASAP7_75t_L g2936 ( 
.A1(n_2925),
.A2(n_103),
.B(n_104),
.C(n_105),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2919),
.Y(n_2937)
);

OAI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_2917),
.A2(n_2168),
.B1(n_2157),
.B2(n_2174),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2917),
.A2(n_696),
.B1(n_699),
.B2(n_700),
.Y(n_2939)
);

NAND4xp25_ASAP7_75t_L g2940 ( 
.A(n_2917),
.B(n_104),
.C(n_106),
.D(n_107),
.Y(n_2940)
);

NOR2x1_ASAP7_75t_L g2941 ( 
.A(n_2931),
.B(n_106),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_SL g2942 ( 
.A1(n_2937),
.A2(n_704),
.B1(n_709),
.B2(n_109),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2927),
.B(n_107),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2934),
.A2(n_2182),
.B1(n_2203),
.B2(n_2210),
.Y(n_2944)
);

AOI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2935),
.A2(n_2182),
.B1(n_110),
.B2(n_111),
.Y(n_2945)
);

OAI211xp5_ASAP7_75t_SL g2946 ( 
.A1(n_2933),
.A2(n_108),
.B(n_111),
.C(n_112),
.Y(n_2946)
);

NAND4xp25_ASAP7_75t_L g2947 ( 
.A(n_2930),
.B(n_108),
.C(n_112),
.D(n_113),
.Y(n_2947)
);

OA21x2_ASAP7_75t_L g2948 ( 
.A1(n_2926),
.A2(n_113),
.B(n_114),
.Y(n_2948)
);

AOI221x1_ASAP7_75t_L g2949 ( 
.A1(n_2932),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_2949)
);

OAI211xp5_ASAP7_75t_L g2950 ( 
.A1(n_2941),
.A2(n_2939),
.B(n_2940),
.C(n_2936),
.Y(n_2950)
);

INVxp67_ASAP7_75t_SL g2951 ( 
.A(n_2948),
.Y(n_2951)
);

AOI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2946),
.A2(n_2928),
.B1(n_2929),
.B2(n_2938),
.Y(n_2952)
);

NOR3xp33_ASAP7_75t_L g2953 ( 
.A(n_2943),
.B(n_116),
.C(n_118),
.Y(n_2953)
);

NAND4xp25_ASAP7_75t_L g2954 ( 
.A(n_2949),
.B(n_119),
.C(n_121),
.D(n_122),
.Y(n_2954)
);

NOR2x1_ASAP7_75t_L g2955 ( 
.A(n_2948),
.B(n_2947),
.Y(n_2955)
);

NAND4xp25_ASAP7_75t_L g2956 ( 
.A(n_2945),
.B(n_119),
.C(n_122),
.D(n_123),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2942),
.B(n_123),
.Y(n_2957)
);

INVx1_ASAP7_75t_SL g2958 ( 
.A(n_2944),
.Y(n_2958)
);

AND3x1_ASAP7_75t_L g2959 ( 
.A(n_2941),
.B(n_124),
.C(n_125),
.Y(n_2959)
);

AOI211xp5_ASAP7_75t_L g2960 ( 
.A1(n_2946),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_2960)
);

NOR4xp25_ASAP7_75t_L g2961 ( 
.A(n_2943),
.B(n_130),
.C(n_131),
.D(n_132),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2941),
.Y(n_2962)
);

NAND5xp2_ASAP7_75t_L g2963 ( 
.A(n_2945),
.B(n_133),
.C(n_134),
.D(n_135),
.E(n_141),
.Y(n_2963)
);

OAI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2945),
.A2(n_133),
.B1(n_134),
.B2(n_1959),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2941),
.B(n_2144),
.Y(n_2965)
);

XNOR2xp5_ASAP7_75t_L g2966 ( 
.A(n_2941),
.B(n_147),
.Y(n_2966)
);

OAI211xp5_ASAP7_75t_SL g2967 ( 
.A1(n_2941),
.A2(n_870),
.B(n_861),
.C(n_166),
.Y(n_2967)
);

XNOR2x1_ASAP7_75t_L g2968 ( 
.A(n_2941),
.B(n_152),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2941),
.B(n_2144),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2941),
.B(n_2144),
.Y(n_2970)
);

AOI321xp33_ASAP7_75t_L g2971 ( 
.A1(n_2941),
.A2(n_163),
.A3(n_170),
.B1(n_173),
.B2(n_174),
.C(n_179),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2959),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2951),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2968),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2966),
.Y(n_2975)
);

AOI22x1_ASAP7_75t_L g2976 ( 
.A1(n_2962),
.A2(n_918),
.B1(n_908),
.B2(n_897),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2954),
.Y(n_2977)
);

AOI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2953),
.A2(n_918),
.B1(n_908),
.B2(n_2021),
.Y(n_2978)
);

INVxp67_ASAP7_75t_SL g2979 ( 
.A(n_2955),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2960),
.B(n_180),
.Y(n_2980)
);

OAI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2952),
.A2(n_2029),
.B1(n_918),
.B2(n_908),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2965),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_R g2983 ( 
.A(n_2958),
.B(n_185),
.Y(n_2983)
);

XOR2xp5_ASAP7_75t_L g2984 ( 
.A(n_2956),
.B(n_187),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2969),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2970),
.A2(n_918),
.B1(n_908),
.B2(n_861),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2957),
.A2(n_918),
.B(n_908),
.Y(n_2987)
);

OR3x1_ASAP7_75t_L g2988 ( 
.A(n_2963),
.B(n_195),
.C(n_198),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2961),
.B(n_1305),
.Y(n_2989)
);

OAI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2964),
.A2(n_1307),
.B1(n_1305),
.B2(n_870),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2950),
.B(n_199),
.Y(n_2991)
);

OAI21x1_ASAP7_75t_L g2992 ( 
.A1(n_2971),
.A2(n_2967),
.B(n_2051),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2959),
.Y(n_2993)
);

INVx4_ASAP7_75t_L g2994 ( 
.A(n_2962),
.Y(n_2994)
);

AOI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2951),
.A2(n_888),
.B(n_1122),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2959),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2968),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2959),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2951),
.B(n_204),
.Y(n_2999)
);

CKINVDCx20_ASAP7_75t_R g3000 ( 
.A(n_2952),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_SL g3001 ( 
.A1(n_2952),
.A2(n_208),
.B(n_210),
.Y(n_3001)
);

OAI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2955),
.A2(n_2051),
.B(n_1998),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2979),
.B(n_211),
.Y(n_3003)
);

OR2x2_ASAP7_75t_L g3004 ( 
.A(n_2999),
.B(n_2991),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2973),
.Y(n_3005)
);

INVxp67_ASAP7_75t_L g3006 ( 
.A(n_2984),
.Y(n_3006)
);

AOI22xp5_ASAP7_75t_SL g3007 ( 
.A1(n_3000),
.A2(n_212),
.B1(n_216),
.B2(n_218),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2994),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2988),
.Y(n_3009)
);

OAI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2972),
.A2(n_1307),
.B1(n_1305),
.B2(n_888),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2993),
.Y(n_3011)
);

AND2x2_ASAP7_75t_SL g3012 ( 
.A(n_2996),
.B(n_219),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2998),
.Y(n_3013)
);

INVx1_ASAP7_75t_SL g3014 ( 
.A(n_2983),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2977),
.A2(n_1307),
.B1(n_1423),
.B2(n_1072),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2980),
.Y(n_3016)
);

NAND5xp2_ASAP7_75t_L g3017 ( 
.A(n_2982),
.B(n_221),
.C(n_223),
.D(n_224),
.E(n_229),
.Y(n_3017)
);

OAI222xp33_ASAP7_75t_L g3018 ( 
.A1(n_2994),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.C1(n_236),
.C2(n_244),
.Y(n_3018)
);

HB1xp67_ASAP7_75t_L g3019 ( 
.A(n_2985),
.Y(n_3019)
);

XOR2xp5_ASAP7_75t_L g3020 ( 
.A(n_2975),
.B(n_253),
.Y(n_3020)
);

OAI221xp5_ASAP7_75t_R g3021 ( 
.A1(n_2978),
.A2(n_254),
.B1(n_255),
.B2(n_262),
.C(n_264),
.Y(n_3021)
);

OAI322xp33_ASAP7_75t_L g3022 ( 
.A1(n_2989),
.A2(n_265),
.A3(n_267),
.B1(n_269),
.B2(n_270),
.C1(n_272),
.C2(n_274),
.Y(n_3022)
);

AOI221xp5_ASAP7_75t_L g3023 ( 
.A1(n_2990),
.A2(n_1122),
.B1(n_1072),
.B2(n_1092),
.C(n_987),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2974),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2997),
.A2(n_1122),
.B1(n_1092),
.B2(n_1072),
.Y(n_3025)
);

NAND5xp2_ASAP7_75t_L g3026 ( 
.A(n_3001),
.B(n_276),
.C(n_277),
.D(n_278),
.E(n_281),
.Y(n_3026)
);

XNOR2xp5_ASAP7_75t_L g3027 ( 
.A(n_2986),
.B(n_282),
.Y(n_3027)
);

NAND3xp33_ASAP7_75t_L g3028 ( 
.A(n_2987),
.B(n_987),
.C(n_1023),
.Y(n_3028)
);

NAND3xp33_ASAP7_75t_L g3029 ( 
.A(n_2976),
.B(n_987),
.C(n_1023),
.Y(n_3029)
);

OAI211xp5_ASAP7_75t_L g3030 ( 
.A1(n_2995),
.A2(n_287),
.B(n_293),
.C(n_307),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2992),
.B(n_308),
.Y(n_3031)
);

BUFx3_ASAP7_75t_L g3032 ( 
.A(n_2981),
.Y(n_3032)
);

INVxp33_ASAP7_75t_L g3033 ( 
.A(n_3002),
.Y(n_3033)
);

NAND4xp25_ASAP7_75t_SL g3034 ( 
.A(n_2991),
.B(n_309),
.C(n_315),
.D(n_321),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_3008),
.Y(n_3035)
);

HB1xp67_ASAP7_75t_L g3036 ( 
.A(n_3008),
.Y(n_3036)
);

OAI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_3005),
.A2(n_327),
.B(n_329),
.Y(n_3037)
);

AOI22xp33_ASAP7_75t_SL g3038 ( 
.A1(n_3019),
.A2(n_3013),
.B1(n_3011),
.B2(n_3024),
.Y(n_3038)
);

XNOR2xp5_ASAP7_75t_L g3039 ( 
.A(n_3014),
.B(n_330),
.Y(n_3039)
);

INVx8_ASAP7_75t_L g3040 ( 
.A(n_3006),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_3012),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_3003),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_3031),
.Y(n_3043)
);

INVxp67_ASAP7_75t_L g3044 ( 
.A(n_3020),
.Y(n_3044)
);

OAI22xp5_ASAP7_75t_SL g3045 ( 
.A1(n_3009),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_3045)
);

AOI221xp5_ASAP7_75t_SL g3046 ( 
.A1(n_3010),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.C(n_343),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_3004),
.Y(n_3047)
);

OAI21x1_ASAP7_75t_L g3048 ( 
.A1(n_3027),
.A2(n_1998),
.B(n_1949),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_SL g3049 ( 
.A1(n_3016),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_3032),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_3036),
.A2(n_3033),
.B(n_3026),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_3035),
.A2(n_3034),
.B(n_3025),
.Y(n_3052)
);

OAI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_3038),
.A2(n_3044),
.B(n_3050),
.Y(n_3053)
);

OA21x2_ASAP7_75t_L g3054 ( 
.A1(n_3041),
.A2(n_3023),
.B(n_3028),
.Y(n_3054)
);

AOI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_3047),
.A2(n_3030),
.B1(n_3015),
.B2(n_3029),
.Y(n_3055)
);

CKINVDCx20_ASAP7_75t_R g3056 ( 
.A(n_3040),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_3040),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_3042),
.A2(n_3017),
.B(n_3007),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_SL g3059 ( 
.A1(n_3043),
.A2(n_3021),
.B1(n_3022),
.B2(n_3018),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_3045),
.A2(n_1023),
.B1(n_1078),
.B2(n_1037),
.Y(n_3060)
);

OAI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_3046),
.A2(n_350),
.B(n_352),
.Y(n_3061)
);

AOI222xp33_ASAP7_75t_L g3062 ( 
.A1(n_3049),
.A2(n_355),
.B1(n_358),
.B2(n_361),
.C1(n_362),
.C2(n_367),
.Y(n_3062)
);

AOI21x1_ASAP7_75t_L g3063 ( 
.A1(n_3051),
.A2(n_3053),
.B(n_3052),
.Y(n_3063)
);

AOI31xp67_ASAP7_75t_L g3064 ( 
.A1(n_3055),
.A2(n_3039),
.A3(n_3037),
.B(n_3048),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_SL g3065 ( 
.A1(n_3056),
.A2(n_374),
.B1(n_376),
.B2(n_379),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_3058),
.A2(n_380),
.B(n_382),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_3057),
.B(n_2072),
.Y(n_3067)
);

AOI221xp5_ASAP7_75t_L g3068 ( 
.A1(n_3060),
.A2(n_1092),
.B1(n_1023),
.B2(n_1078),
.C(n_1106),
.Y(n_3068)
);

A2O1A1Ixp33_ASAP7_75t_L g3069 ( 
.A1(n_3061),
.A2(n_383),
.B(n_384),
.C(n_385),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3059),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_3054),
.B(n_3062),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_3051),
.A2(n_386),
.B(n_387),
.Y(n_3072)
);

INVx1_ASAP7_75t_SL g3073 ( 
.A(n_3070),
.Y(n_3073)
);

INVxp67_ASAP7_75t_L g3074 ( 
.A(n_3071),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_3064),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3063),
.Y(n_3076)
);

INVxp67_ASAP7_75t_L g3077 ( 
.A(n_3072),
.Y(n_3077)
);

OR2x2_ASAP7_75t_L g3078 ( 
.A(n_3073),
.B(n_3069),
.Y(n_3078)
);

OAI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_3074),
.A2(n_3068),
.B(n_3067),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_3075),
.B(n_3066),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_3080),
.A2(n_3076),
.B(n_3077),
.Y(n_3081)
);

AOI211xp5_ASAP7_75t_L g3082 ( 
.A1(n_3081),
.A2(n_3078),
.B(n_3079),
.C(n_3065),
.Y(n_3082)
);


endmodule