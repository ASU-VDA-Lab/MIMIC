module fake_aes_9100_n_870 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_870);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_870;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g109 ( .A(n_68), .Y(n_109) );
BUFx5_ASAP7_75t_L g110 ( .A(n_95), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_89), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_97), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_40), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_21), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_74), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_47), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_88), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_67), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_60), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_51), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_6), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_32), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_44), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_1), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_59), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_6), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_12), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_49), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_69), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_9), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_80), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_65), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_78), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
BUFx2_ASAP7_75t_SL g140 ( .A(n_79), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_16), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_50), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_53), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_31), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_26), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_24), .Y(n_147) );
CKINVDCx14_ASAP7_75t_R g148 ( .A(n_29), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_142), .B(n_0), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_118), .B(n_18), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_110), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_137), .B(n_0), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_134), .B(n_1), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_139), .B(n_2), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_137), .B(n_2), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
BUFx12f_ASAP7_75t_L g163 ( .A(n_111), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_129), .B(n_3), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_129), .B(n_3), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_123), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
BUFx8_ASAP7_75t_SL g172 ( .A(n_125), .Y(n_172) );
BUFx8_ASAP7_75t_SL g173 ( .A(n_127), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_141), .B(n_4), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_120), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_167), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_173), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_169), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_172), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_163), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_163), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_163), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_158), .A2(n_140), .B1(n_122), .B2(n_131), .Y(n_186) );
NOR2xp33_ASAP7_75t_R g187 ( .A(n_164), .B(n_114), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_164), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_165), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_165), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_150), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_150), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_154), .B(n_157), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_150), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_154), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_157), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_170), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_170), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_159), .Y(n_202) );
NOR2xp67_ASAP7_75t_L g203 ( .A(n_171), .B(n_121), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_171), .Y(n_204) );
NAND2xp33_ASAP7_75t_R g205 ( .A(n_161), .B(n_112), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_161), .Y(n_206) );
AOI21x1_ASAP7_75t_L g207 ( .A1(n_152), .A2(n_149), .B(n_131), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_161), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_174), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_160), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_175), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_175), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
INVxp67_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_167), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_151), .Y(n_218) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_152), .A2(n_133), .B(n_109), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_153), .B(n_114), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_151), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_176), .B(n_133), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_151), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_153), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_151), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_151), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_156), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_156), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_151), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_151), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_151), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_210), .B(n_148), .Y(n_235) );
NOR2xp33_ASAP7_75t_R g236 ( .A(n_183), .B(n_148), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_234), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_190), .B(n_126), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_182), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_197), .B(n_113), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_198), .B(n_115), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_196), .Y(n_244) );
BUFx5_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_218), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_211), .B(n_132), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_200), .B(n_116), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g249 ( .A(n_233), .B(n_110), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_201), .B(n_117), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_232), .Y(n_251) );
BUFx5_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_168), .B1(n_128), .B2(n_162), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_204), .B(n_119), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_189), .B(n_126), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_191), .B(n_126), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_214), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_195), .B(n_124), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_193), .B(n_136), .Y(n_260) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_178), .B(n_176), .C(n_168), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_180), .B(n_176), .C(n_168), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_188), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_203), .B(n_138), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_213), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_181), .B(n_128), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_186), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_186), .A2(n_128), .B1(n_167), .B2(n_176), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_206), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_208), .Y(n_273) );
AND2x4_ASAP7_75t_SL g274 ( .A(n_213), .B(n_162), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_194), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_219), .A2(n_166), .B1(n_162), .B2(n_176), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_216), .B(n_143), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_220), .B(n_145), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_222), .Y(n_279) );
INVx6_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_179), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_221), .B(n_176), .C(n_166), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_219), .B(n_153), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_229), .A2(n_155), .B(n_162), .C(n_166), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_187), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
BUFx6f_ASAP7_75t_SL g287 ( .A(n_179), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_212), .B(n_153), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_224), .B(n_153), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_184), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_202), .B(n_153), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_212), .B(n_162), .Y(n_296) );
AO221x1_ASAP7_75t_L g297 ( .A1(n_185), .A2(n_166), .B1(n_155), .B2(n_7), .C(n_8), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_215), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_253), .B(n_223), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_268), .A2(n_166), .B1(n_228), .B2(n_225), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_245), .Y(n_302) );
AO22x1_ASAP7_75t_L g303 ( .A1(n_265), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_265), .Y(n_304) );
BUFx4f_ASAP7_75t_L g305 ( .A(n_237), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_287), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_245), .B(n_226), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_287), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_281), .Y(n_309) );
AO21x1_ASAP7_75t_L g310 ( .A1(n_269), .A2(n_227), .B(n_217), .Y(n_310) );
NOR2x1p5_ASAP7_75t_L g311 ( .A(n_241), .B(n_166), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_269), .A2(n_155), .B1(n_217), .B2(n_215), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_238), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_274), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
BUFx10_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_244), .B(n_155), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_236), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_245), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_270), .B(n_5), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_275), .B(n_273), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_279), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_235), .A2(n_110), .B1(n_227), .B2(n_226), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_252), .B(n_226), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_256), .B(n_8), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_252), .B(n_110), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_291), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_252), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
AOI22xp33_ASAP7_75t_SL g337 ( .A1(n_297), .A2(n_110), .B1(n_10), .B2(n_11), .Y(n_337) );
OAI22xp5_ASAP7_75t_SL g338 ( .A1(n_267), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_338) );
INVx5_ASAP7_75t_L g339 ( .A(n_238), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_247), .B(n_13), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_243), .B(n_13), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_248), .B(n_14), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_239), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_271), .Y(n_344) );
INVx5_ASAP7_75t_L g345 ( .A(n_238), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_254), .B(n_107), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_283), .B(n_249), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_336), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_321), .B(n_285), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_SL g350 ( .A1(n_329), .A2(n_296), .B(n_288), .C(n_260), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_323), .B(n_257), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_322), .B(n_250), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_321), .B(n_255), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_307), .A2(n_278), .B(n_259), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_340), .A2(n_266), .B(n_293), .C(n_242), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_321), .A2(n_277), .B1(n_261), .B2(n_262), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_SL g357 ( .A1(n_333), .A2(n_284), .B(n_290), .C(n_282), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_305), .B(n_264), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_302), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_SL g360 ( .A1(n_333), .A2(n_282), .B(n_262), .C(n_261), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_276), .B(n_294), .C(n_295), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_337), .A2(n_251), .B1(n_246), .B2(n_280), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_325), .B(n_246), .Y(n_365) );
AO32x2_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .Y(n_366) );
OR2x6_ASAP7_75t_L g367 ( .A(n_331), .B(n_251), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_251), .B(n_246), .C(n_298), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_305), .B(n_15), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_327), .A2(n_280), .B(n_19), .Y(n_370) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_302), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_305), .B(n_17), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_304), .A2(n_20), .B(n_22), .C(n_23), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_334), .B(n_25), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_27), .B(n_28), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_370), .A2(n_310), .B(n_346), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_346), .B(n_320), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_354), .A2(n_326), .B(n_300), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_374), .A2(n_320), .B(n_330), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_352), .B(n_315), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_348), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_372), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_344), .B(n_343), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
BUFx12f_ASAP7_75t_SL g390 ( .A(n_349), .Y(n_390) );
BUFx2_ASAP7_75t_SL g391 ( .A(n_376), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_362), .A2(n_344), .B(n_328), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_364), .B(n_315), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_351), .B(n_309), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
AOI22x1_ASAP7_75t_L g396 ( .A1(n_377), .A2(n_311), .B1(n_313), .B2(n_320), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_349), .A2(n_338), .B1(n_314), .B2(n_332), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_361), .A2(n_301), .B(n_335), .Y(n_400) );
INVx6_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_353), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_369), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_301), .B(n_335), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_365), .B(n_319), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_400), .A2(n_356), .B(n_330), .Y(n_414) );
BUFx10_ASAP7_75t_L g415 ( .A(n_409), .Y(n_415) );
AOI21x1_ASAP7_75t_L g416 ( .A1(n_383), .A2(n_303), .B(n_358), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_357), .B(n_350), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_393), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_397), .A2(n_375), .B1(n_309), .B2(n_308), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_397), .A2(n_306), .B1(n_308), .B2(n_316), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
CKINVDCx6p67_ASAP7_75t_R g422 ( .A(n_402), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_385), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_404), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_299), .B(n_360), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_386), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_408), .A2(n_316), .B1(n_318), .B2(n_319), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g429 ( .A1(n_402), .A2(n_316), .B1(n_318), .B2(n_339), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_402), .A2(n_345), .B1(n_339), .B2(n_313), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_404), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_398), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
AOI21x1_ASAP7_75t_L g439 ( .A1(n_383), .A2(n_355), .B(n_313), .Y(n_439) );
CKINVDCx11_ASAP7_75t_R g440 ( .A(n_405), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_378), .A2(n_317), .B(n_313), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_388), .A2(n_317), .B(n_345), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_393), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_403), .B(n_345), .Y(n_444) );
CKINVDCx11_ASAP7_75t_R g445 ( .A(n_405), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_403), .B(n_345), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
INVx4_ASAP7_75t_SL g451 ( .A(n_401), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_345), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_392), .A2(n_339), .B(n_33), .Y(n_453) );
OAI21x1_ASAP7_75t_L g454 ( .A1(n_378), .A2(n_339), .B(n_34), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
AOI21x1_ASAP7_75t_L g456 ( .A1(n_383), .A2(n_339), .B(n_35), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_391), .A2(n_30), .B1(n_36), .B2(n_37), .Y(n_457) );
OAI21x1_ASAP7_75t_L g458 ( .A1(n_378), .A2(n_38), .B(n_39), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
OAI21x1_ASAP7_75t_L g460 ( .A1(n_379), .A2(n_41), .B(n_42), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_407), .Y(n_461) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_392), .A2(n_43), .B(n_45), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_381), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_391), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_393), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_413), .B(n_405), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_451), .B(n_389), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_423), .B(n_389), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_435), .A2(n_408), .B1(n_406), .B2(n_390), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_415), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_440), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_453), .B(n_390), .C(n_384), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_444), .B(n_409), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_445), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_446), .B(n_409), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_446), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_415), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_451), .B(n_389), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_452), .B(n_409), .Y(n_483) );
NOR2xp33_ASAP7_75t_R g484 ( .A(n_422), .B(n_410), .Y(n_484) );
NOR3xp33_ASAP7_75t_SL g485 ( .A(n_453), .B(n_384), .C(n_410), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_409), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_424), .B(n_406), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_422), .Y(n_488) );
NOR2xp33_ASAP7_75t_R g489 ( .A(n_465), .B(n_410), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_412), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_437), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_451), .B(n_389), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_447), .Y(n_494) );
NOR2xp33_ASAP7_75t_R g495 ( .A(n_465), .B(n_410), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_425), .A2(n_406), .B1(n_401), .B2(n_380), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_464), .A2(n_393), .B1(n_401), .B2(n_396), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_427), .B(n_382), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
NAND2xp33_ASAP7_75t_R g500 ( .A(n_465), .B(n_382), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
NOR2xp33_ASAP7_75t_R g502 ( .A(n_465), .B(n_401), .Y(n_502) );
NAND2xp33_ASAP7_75t_R g503 ( .A(n_464), .B(n_382), .Y(n_503) );
OAI21x1_ASAP7_75t_SL g504 ( .A1(n_418), .A2(n_396), .B(n_407), .Y(n_504) );
AO31x2_ASAP7_75t_L g505 ( .A1(n_432), .A2(n_379), .A3(n_380), .B(n_382), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_415), .B(n_401), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_427), .B(n_449), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_412), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_448), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_449), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_434), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_421), .B(n_381), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_455), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_421), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_421), .A2(n_381), .B1(n_379), .B2(n_52), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_430), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_419), .A2(n_46), .B1(n_48), .B2(n_54), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_455), .B(n_106), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_418), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_420), .B(n_56), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_430), .B(n_57), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_433), .B(n_58), .Y(n_522) );
NAND3xp33_ASAP7_75t_SL g523 ( .A(n_428), .B(n_61), .C(n_62), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_451), .B(n_63), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_443), .A2(n_64), .B(n_66), .C(n_70), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_451), .B(n_71), .Y(n_527) );
CKINVDCx11_ASAP7_75t_R g528 ( .A(n_463), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_433), .B(n_72), .Y(n_529) );
NAND3xp33_ASAP7_75t_SL g530 ( .A(n_429), .B(n_73), .C(n_75), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_443), .B(n_76), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_431), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_436), .B(n_77), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_438), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_438), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_450), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_457), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_537) );
NOR3xp33_ASAP7_75t_SL g538 ( .A(n_462), .B(n_85), .C(n_86), .Y(n_538) );
NOR3xp33_ASAP7_75t_SL g539 ( .A(n_462), .B(n_87), .C(n_90), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_463), .B(n_105), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_92), .Y(n_541) );
AO32x2_ASAP7_75t_L g542 ( .A1(n_417), .A2(n_94), .A3(n_96), .B1(n_99), .B2(n_100), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_463), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_442), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_450), .Y(n_545) );
AO32x2_ASAP7_75t_L g546 ( .A1(n_417), .A2(n_101), .A3(n_102), .B1(n_104), .B2(n_450), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_442), .A2(n_417), .B1(n_462), .B2(n_461), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_454), .A2(n_460), .B(n_458), .C(n_441), .Y(n_548) );
AO31x2_ASAP7_75t_L g549 ( .A1(n_432), .A2(n_461), .A3(n_459), .B(n_416), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_432), .Y(n_550) );
NOR3xp33_ASAP7_75t_SL g551 ( .A(n_456), .B(n_416), .C(n_458), .Y(n_551) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_456), .A2(n_454), .B(n_441), .Y(n_552) );
OR2x6_ASAP7_75t_L g553 ( .A(n_460), .B(n_459), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_511), .Y(n_554) );
NOR2x1_ASAP7_75t_SL g555 ( .A(n_499), .B(n_442), .Y(n_555) );
OR2x2_ASAP7_75t_SL g556 ( .A(n_509), .B(n_414), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_473), .B(n_459), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_461), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_543), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_494), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_476), .B(n_414), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_501), .B(n_414), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_475), .A2(n_486), .B1(n_483), .B2(n_478), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_510), .B(n_414), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_532), .A2(n_426), .B1(n_439), .B2(n_470), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_482), .B(n_426), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_553), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_513), .B(n_439), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_426), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_466), .B(n_487), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_487), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_496), .A2(n_520), .B1(n_469), .B2(n_506), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_535), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_477), .B(n_471), .Y(n_576) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_468), .B(n_530), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_536), .B(n_545), .Y(n_578) );
INVx4_ASAP7_75t_L g579 ( .A(n_480), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_512), .B(n_508), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_498), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_474), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_489), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_498), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_490), .B(n_514), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_549), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_549), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_521), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_549), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_505), .B(n_544), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_505), .B(n_553), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
AOI31xp33_ASAP7_75t_L g595 ( .A1(n_488), .A2(n_503), .A3(n_484), .B(n_500), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_495), .B(n_485), .Y(n_596) );
BUFx3_ASAP7_75t_L g597 ( .A(n_528), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_553), .B(n_547), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_467), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_531), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_472), .B(n_502), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_522), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_467), .B(n_481), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_525), .B(n_533), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_525), .B(n_492), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_492), .B(n_541), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_531), .A2(n_523), .B1(n_524), .B2(n_527), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_497), .B(n_546), .Y(n_611) );
NOR2x1_ASAP7_75t_SL g612 ( .A(n_497), .B(n_540), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_546), .B(n_551), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_504), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_515), .B(n_548), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_552), .B(n_515), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_526), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_538), .A2(n_539), .B(n_517), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_542), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_537), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_542), .B(n_491), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_491), .B(n_493), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_511), .B(n_435), .Y(n_624) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_470), .B(n_480), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_491), .B(n_493), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_511), .Y(n_627) );
INVx3_ASAP7_75t_SL g628 ( .A(n_488), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_534), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_511), .B(n_507), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_476), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_534), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_534), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_534), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_491), .B(n_493), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_511), .B(n_507), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_491), .B(n_493), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_491), .B(n_493), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
AO21x2_ASAP7_75t_L g642 ( .A1(n_551), .A2(n_504), .B(n_548), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_491), .B(n_493), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_491), .B(n_493), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_534), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_528), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_534), .Y(n_647) );
INVx3_ASAP7_75t_SL g648 ( .A(n_488), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_491), .B(n_493), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_511), .Y(n_650) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_519), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_491), .B(n_493), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_491), .B(n_493), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_511), .B(n_435), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_569), .B(n_631), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_637), .B(n_554), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_627), .B(n_639), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_624), .A2(n_654), .B(n_565), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_650), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_560), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_572), .B(n_578), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_609), .B(n_563), .Y(n_663) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_587), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_578), .B(n_557), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_581), .B(n_651), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_606), .B(n_566), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_606), .B(n_599), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_582), .B(n_585), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_623), .B(n_626), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_636), .B(n_638), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_640), .B(n_643), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_575), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_625), .B(n_595), .Y(n_675) );
NAND2x1_ASAP7_75t_SL g676 ( .A(n_628), .B(n_648), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_614), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_629), .Y(n_678) );
OA21x2_ASAP7_75t_L g679 ( .A1(n_593), .A2(n_590), .B(n_588), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_644), .B(n_649), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_644), .B(n_649), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_652), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_652), .B(n_653), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_653), .B(n_559), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_629), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_630), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_555), .B(n_568), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_568), .B(n_598), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_573), .B(n_632), .Y(n_689) );
AND2x4_ASAP7_75t_SL g690 ( .A(n_579), .B(n_600), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_562), .B(n_564), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_625), .A2(n_579), .B1(n_584), .B2(n_612), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_605), .B(n_603), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_579), .B(n_597), .Y(n_694) );
BUFx3_ASAP7_75t_L g695 ( .A(n_597), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_646), .B(n_654), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_630), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_646), .B(n_624), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_577), .B(n_610), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_586), .B(n_558), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_633), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_586), .B(n_558), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_633), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_589), .B(n_604), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_628), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_594), .B(n_602), .Y(n_707) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_611), .B(n_615), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_607), .B(n_641), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_635), .Y(n_710) );
INVx4_ASAP7_75t_L g711 ( .A(n_648), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_641), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_596), .B(n_613), .Y(n_713) );
AOI221x1_ASAP7_75t_L g714 ( .A1(n_619), .A2(n_613), .B1(n_620), .B2(n_616), .C(n_601), .Y(n_714) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_574), .A2(n_615), .B1(n_611), .B2(n_598), .C(n_621), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_645), .B(n_647), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_583), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_580), .Y(n_718) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_618), .B(n_621), .C(n_622), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_564), .B(n_622), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_568), .B(n_620), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_576), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_571), .B(n_561), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_571), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_587), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_567), .Y(n_726) );
INVx4_ASAP7_75t_L g727 ( .A(n_608), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_556), .B(n_592), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_591), .B(n_592), .Y(n_729) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_588), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_608), .B(n_617), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_709), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_705), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_691), .B(n_570), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_708), .A2(n_642), .B1(n_570), .B2(n_593), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_691), .B(n_642), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_667), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_695), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_720), .B(n_642), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_700), .B(n_702), .Y(n_740) );
BUFx2_ASAP7_75t_L g741 ( .A(n_676), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_711), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_657), .B(n_655), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_672), .B(n_680), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_731), .B(n_708), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_711), .B(n_695), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_724), .B(n_661), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_665), .B(n_729), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_692), .B(n_687), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_682), .B(n_693), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_694), .Y(n_751) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_711), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_687), .B(n_688), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_660), .B(n_671), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_684), .B(n_673), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_696), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_681), .B(n_683), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_662), .B(n_723), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_688), .B(n_668), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_722), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_659), .B(n_726), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_713), .B(n_712), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_713), .B(n_712), .Y(n_763) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_698), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_663), .B(n_670), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_658), .B(n_666), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_728), .B(n_667), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_689), .Y(n_768) );
AND2x4_ASAP7_75t_L g769 ( .A(n_687), .B(n_656), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_704), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_728), .B(n_669), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_707), .Y(n_772) );
BUFx3_ASAP7_75t_L g773 ( .A(n_690), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_719), .B(n_716), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_719), .B(n_690), .Y(n_775) );
AND4x1_ASAP7_75t_L g776 ( .A(n_714), .B(n_675), .C(n_692), .D(n_699), .Y(n_776) );
INVxp67_ASAP7_75t_L g777 ( .A(n_675), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_703), .B(n_706), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_748), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_737), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_771), .B(n_656), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_748), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_778), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_777), .A2(n_699), .B1(n_656), .B2(n_677), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_771), .B(n_677), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_734), .B(n_677), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_761), .B(n_710), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_735), .A2(n_721), .B1(n_727), .B2(n_725), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_758), .B(n_715), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_773), .B(n_727), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_732), .B(n_717), .Y(n_791) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_764), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_749), .A2(n_721), .B1(n_727), .B2(n_718), .Y(n_793) );
XNOR2x2_ASAP7_75t_L g794 ( .A(n_749), .B(n_715), .Y(n_794) );
INVxp67_ASAP7_75t_L g795 ( .A(n_760), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_736), .A2(n_664), .B1(n_730), .B2(n_725), .C(n_701), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g797 ( .A(n_776), .B(n_679), .C(n_730), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_773), .A2(n_686), .B1(n_674), .B2(n_678), .Y(n_798) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_752), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_733), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_758), .B(n_686), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_733), .B(n_685), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_747), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_747), .Y(n_804) );
OAI32xp33_ASAP7_75t_L g805 ( .A1(n_775), .A2(n_742), .A3(n_774), .B1(n_746), .B2(n_738), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_743), .B(n_697), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_750), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_770), .B(n_697), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_752), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_808), .Y(n_810) );
OAI21xp33_ASAP7_75t_L g811 ( .A1(n_789), .A2(n_736), .B(n_767), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_808), .Y(n_812) );
OAI221xp5_ASAP7_75t_SL g813 ( .A1(n_792), .A2(n_741), .B1(n_742), .B2(n_774), .C(n_756), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_791), .Y(n_814) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_780), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_801), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_784), .A2(n_751), .B(n_762), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_791), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_787), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_795), .A2(n_767), .B1(n_739), .B2(n_745), .Y(n_820) );
INVx1_ASAP7_75t_SL g821 ( .A(n_800), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_787), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_783), .Y(n_823) );
OAI21xp33_ASAP7_75t_L g824 ( .A1(n_805), .A2(n_739), .B(n_745), .Y(n_824) );
AOI21xp33_ASAP7_75t_SL g825 ( .A1(n_790), .A2(n_751), .B(n_769), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_797), .A2(n_752), .B(n_769), .Y(n_826) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_794), .B(n_766), .Y(n_827) );
OAI31xp33_ASAP7_75t_L g828 ( .A1(n_790), .A2(n_762), .A3(n_763), .B(n_769), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_798), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_779), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_782), .A2(n_763), .B1(n_752), .B2(n_753), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_816), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g833 ( .A1(n_826), .A2(n_793), .B(n_788), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_815), .Y(n_834) );
OAI22xp33_ASAP7_75t_SL g835 ( .A1(n_813), .A2(n_799), .B1(n_798), .B2(n_766), .Y(n_835) );
AOI32xp33_ASAP7_75t_L g836 ( .A1(n_824), .A2(n_796), .A3(n_802), .B1(n_785), .B2(n_781), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_814), .B(n_807), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_815), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_817), .B(n_786), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_828), .B(n_734), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_819), .B(n_806), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_827), .A2(n_797), .B1(n_753), .B2(n_772), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_813), .A2(n_753), .B1(n_765), .B2(n_757), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_834), .B(n_822), .Y(n_844) );
INVx2_ASAP7_75t_SL g845 ( .A(n_832), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_835), .A2(n_836), .B1(n_833), .B2(n_843), .C(n_829), .Y(n_846) );
NOR3x1_ASAP7_75t_L g847 ( .A(n_838), .B(n_809), .C(n_823), .Y(n_847) );
NOR2x1_ASAP7_75t_L g848 ( .A(n_840), .B(n_826), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_837), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_844), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_849), .B(n_842), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_847), .B(n_839), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g853 ( .A(n_846), .B(n_836), .C(n_811), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_852), .B(n_821), .Y(n_854) );
A2O1A1Ixp33_ASAP7_75t_L g855 ( .A1(n_853), .A2(n_848), .B(n_845), .C(n_825), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_850), .B(n_831), .Y(n_856) );
INVxp67_ASAP7_75t_L g857 ( .A(n_854), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_856), .Y(n_858) );
AOI31xp33_ASAP7_75t_L g859 ( .A1(n_857), .A2(n_855), .A3(n_851), .B(n_820), .Y(n_859) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_858), .B(n_841), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_860), .Y(n_861) );
INVx1_ASAP7_75t_SL g862 ( .A(n_859), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_861), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_863), .Y(n_864) );
AO22x2_ASAP7_75t_L g865 ( .A1(n_864), .A2(n_862), .B1(n_830), .B2(n_818), .Y(n_865) );
OAI22xp5_ASAP7_75t_SL g866 ( .A1(n_865), .A2(n_812), .B1(n_810), .B2(n_768), .Y(n_866) );
AOI21xp33_ASAP7_75t_SL g867 ( .A1(n_866), .A2(n_754), .B(n_803), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_867), .A2(n_804), .B1(n_755), .B2(n_759), .Y(n_868) );
XNOR2xp5_ASAP7_75t_L g869 ( .A(n_868), .B(n_755), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_869), .A2(n_759), .B1(n_740), .B2(n_744), .Y(n_870) );
endmodule