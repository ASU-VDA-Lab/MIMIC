module fake_jpeg_29101_n_373 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_373);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_63),
.Y(n_87)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_33),
.A2(n_10),
.B1(n_17),
.B2(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx2_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_84),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_79),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_41),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_109),
.Y(n_142)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_51),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_127),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_43),
.B(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_60),
.B(n_43),
.C(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_34),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_128),
.B(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_42),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_145),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_28),
.B1(n_55),
.B2(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_144),
.B1(n_149),
.B2(n_160),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_152),
.B1(n_159),
.B2(n_94),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_31),
.B1(n_35),
.B2(n_42),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_151),
.Y(n_166)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_75),
.B1(n_80),
.B2(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_25),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_95),
.A2(n_25),
.B1(n_39),
.B2(n_27),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_23),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_39),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_83),
.B1(n_72),
.B2(n_78),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_57),
.B1(n_56),
.B2(n_46),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_176),
.B1(n_178),
.B2(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_104),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_49),
.B1(n_52),
.B2(n_47),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_108),
.B1(n_99),
.B2(n_115),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_184),
.B1(n_168),
.B2(n_121),
.Y(n_201)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_195),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_152),
.C(n_128),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_123),
.B(n_151),
.C(n_146),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_158),
.B1(n_133),
.B2(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_196),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_154),
.B(n_142),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_157),
.B(n_150),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_161),
.B(n_90),
.Y(n_215)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_196),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_141),
.B1(n_125),
.B2(n_121),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_162),
.B1(n_164),
.B2(n_167),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_215),
.B(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_177),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_182),
.B1(n_184),
.B2(n_198),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_230),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_215),
.B1(n_210),
.B2(n_214),
.Y(n_234)
);

NAND2x1_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_190),
.C(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_207),
.C(n_212),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_189),
.B(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_171),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_170),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_202),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_171),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_187),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_211),
.B1(n_216),
.B2(n_210),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_249),
.B1(n_223),
.B2(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.C(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_207),
.C(n_215),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_206),
.B(n_201),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_205),
.B(n_183),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_206),
.C(n_203),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_221),
.B1(n_194),
.B2(n_230),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_220),
.A2(n_224),
.B1(n_202),
.B2(n_217),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_139),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_226),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_254),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_243),
.B1(n_240),
.B2(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_228),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_222),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_267),
.Y(n_289)
);

AND2x4_ASAP7_75t_SL g287 ( 
.A(n_257),
.B(n_148),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_172),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_163),
.C(n_173),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_164),
.B1(n_125),
.B2(n_130),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_163),
.C(n_177),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_205),
.Y(n_265)
);

XOR2x1_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_159),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_179),
.C(n_188),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_90),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_179),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_242),
.B1(n_245),
.B2(n_238),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_162),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_121),
.Y(n_302)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_279),
.B(n_289),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_238),
.B(n_183),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_172),
.C(n_131),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_265),
.C(n_251),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_136),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_288),
.Y(n_304)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_290),
.B1(n_155),
.B2(n_82),
.C(n_124),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_15),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_259),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_296),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_298),
.C(n_305),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_303),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_283),
.C(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_308),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_309),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_15),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_112),
.C(n_143),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_307),
.Y(n_321)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_156),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_297),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_314),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_289),
.B(n_156),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_313),
.A2(n_102),
.B(n_88),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_140),
.B(n_132),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_18),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_325),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_18),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_319),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_295),
.B(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_113),
.C(n_98),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_105),
.C(n_103),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_308),
.B1(n_296),
.B2(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_330),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_321),
.B(n_322),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_329),
.B(n_337),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_108),
.B(n_99),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_41),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_336),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_41),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_320),
.B(n_41),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_75),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_324),
.C(n_312),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_332),
.B(n_312),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_13),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_346),
.A2(n_347),
.B1(n_11),
.B2(n_15),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_37),
.B1(n_101),
.B2(n_97),
.Y(n_347)
);

OAI321xp33_ASAP7_75t_L g348 ( 
.A1(n_331),
.A2(n_12),
.A3(n_16),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_348),
.A2(n_37),
.B1(n_53),
.B2(n_50),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_350),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_37),
.C(n_53),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_353),
.B(n_355),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_37),
.C(n_50),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_11),
.C(n_16),
.Y(n_355)
);

AOI31xp67_ASAP7_75t_SL g356 ( 
.A1(n_344),
.A2(n_342),
.A3(n_338),
.B(n_3),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_356),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_350),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_9),
.C(n_14),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_359),
.B(n_5),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_363),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_9),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_366),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_5),
.Y(n_366)
);

AOI322xp5_ASAP7_75t_L g367 ( 
.A1(n_360),
.A2(n_358),
.A3(n_8),
.B1(n_13),
.B2(n_14),
.C1(n_17),
.C2(n_1),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_369),
.C(n_365),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_8),
.C(n_13),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_372),
.B(n_14),
.Y(n_373)
);


endmodule