module fake_jpeg_28719_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_10),
.B(n_5),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_50),
.Y(n_54)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_2),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_37),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_31),
.C(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_11),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_39),
.B1(n_32),
.B2(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_75),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_33),
.B1(n_36),
.B2(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_4),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_81),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_8),
.B(n_9),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_73),
.B1(n_70),
.B2(n_14),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_12),
.C(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_77),
.C(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_98),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_21),
.B(n_22),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_99),
.C(n_102),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_105),
.B(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_100),
.Y(n_111)
);


endmodule