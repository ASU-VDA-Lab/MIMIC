module fake_netlist_6_1379_n_2405 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2405);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2405;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_437;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2357;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_177),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_133),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_128),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_52),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_73),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_70),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_52),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_62),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_17),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_115),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_112),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_68),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_161),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_23),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_74),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_178),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_211),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_82),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_60),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_61),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_101),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_28),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_222),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_33),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_59),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_203),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_191),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_129),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_120),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_126),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_201),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_154),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_131),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_66),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_142),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_140),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_42),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_213),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_199),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_9),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_181),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_65),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_94),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_169),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_114),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_33),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_107),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_55),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_155),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_72),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_48),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_14),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_30),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_78),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_183),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_59),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_87),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_21),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_102),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_10),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_30),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_176),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_35),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_83),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_91),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_151),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_44),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_18),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_125),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_25),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_117),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_75),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_20),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_67),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_97),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_60),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_89),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_50),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_159),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_205),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_162),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_164),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_97),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_228),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_14),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_216),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_11),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_28),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_56),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_224),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_7),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_186),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_101),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_166),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_23),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_168),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_89),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_62),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_27),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_63),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_138),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_20),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_121),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_212),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_136),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_208),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_150),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_98),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_75),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_91),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_13),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_1),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_69),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_22),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_9),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_50),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_58),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_46),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_221),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_167),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_111),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_173),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_196),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_80),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_157),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_122),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_19),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_104),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_134),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_206),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_0),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_226),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_124),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_102),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_36),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_19),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_24),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_193),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_209),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_83),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_96),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_27),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_72),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_108),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_172),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_144),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_67),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_88),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_81),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_197),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_43),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_35),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_106),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_25),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_76),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_13),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_103),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_194),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_184),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_1),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_210),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_158),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_71),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_160),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_36),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_11),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_99),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_104),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_84),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_43),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_188),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_15),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_71),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_46),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_190),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_137),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_220),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_54),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_171),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_182),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_255),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_263),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_243),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_295),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_229),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_233),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_236),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_240),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_263),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_248),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_251),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_278),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_254),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_260),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_287),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_333),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_295),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_349),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_371),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_265),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_371),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_292),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_257),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_272),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_292),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_241),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_279),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_396),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_323),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_282),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_323),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_263),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_391),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_292),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_318),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_318),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_318),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_410),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_415),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_284),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_286),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_435),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_396),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_289),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_305),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_294),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_383),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_305),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_300),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_395),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_2),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_423),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_428),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_291),
.B(n_2),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_395),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_307),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_336),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_338),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_346),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_347),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_348),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_330),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_351),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_354),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_275),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_275),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_275),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_412),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_3),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_235),
.B(n_4),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_330),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_360),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_361),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_301),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_235),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_329),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_363),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_365),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_372),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_252),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_374),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_375),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_376),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_390),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_393),
.B(n_109),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_252),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_4),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_304),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_269),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_269),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_281),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_281),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_293),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_273),
.B(n_5),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_293),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_298),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_304),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_399),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_257),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_298),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_400),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_230),
.B(n_8),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_402),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_409),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_299),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_329),
.B(n_10),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_416),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_434),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_513),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_452),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_481),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

CKINVDCx8_ASAP7_75t_R g579 ( 
.A(n_554),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_463),
.B(n_421),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_453),
.A2(n_370),
.B(n_230),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_481),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_481),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_458),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_546),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_459),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_463),
.B(n_329),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_466),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_552),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_463),
.B(n_429),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_532),
.B(n_450),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_568),
.B(n_450),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_481),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

BUFx8_ASAP7_75t_L g601 ( 
.A(n_532),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_451),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_460),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_446),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_505),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_469),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_454),
.B(n_450),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_574),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_470),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_556),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_556),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_557),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_464),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_447),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_465),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_565),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_565),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_565),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_467),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_565),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_453),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_529),
.B(n_230),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_454),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

OA21x2_ASAP7_75t_L g629 ( 
.A1(n_457),
.A2(n_404),
.B(n_370),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_468),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_561),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_558),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_489),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_490),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_477),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_559),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_482),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_530),
.B(n_448),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_461),
.B(n_257),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_471),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_553),
.B(n_242),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_471),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_559),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_485),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_475),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_488),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_R g652 ( 
.A(n_520),
.B(n_244),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_490),
.B(n_475),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_499),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_509),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_486),
.B(n_231),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_283),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_566),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_462),
.B(n_434),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_571),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_476),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_476),
.B(n_370),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_500),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_504),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_506),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_474),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_531),
.B(n_404),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_478),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_656),
.B(n_510),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_604),
.B(n_519),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_625),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_640),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_646),
.Y(n_677)
);

INVx6_ASAP7_75t_L g678 ( 
.A(n_653),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_634),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_580),
.B(n_523),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_580),
.B(n_527),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_589),
.B(n_531),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_596),
.B(n_533),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_661),
.B(n_512),
.C(n_502),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_596),
.B(n_533),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_586),
.B(n_528),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_633),
.B(n_456),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_627),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_628),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_628),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_600),
.A2(n_537),
.B1(n_536),
.B2(n_433),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_652),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_628),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_639),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_588),
.B(n_543),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_627),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_639),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_639),
.Y(n_701)
);

AO21x1_ASAP7_75t_L g702 ( 
.A1(n_604),
.A2(n_560),
.B(n_572),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_603),
.B(n_544),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_616),
.B(n_547),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_641),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_617),
.A2(n_484),
.B1(n_487),
.B2(n_472),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_634),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_641),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_643),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_643),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_576),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_577),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_592),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_577),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_596),
.B(n_534),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_645),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_645),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_617),
.A2(n_526),
.B1(n_443),
.B2(n_536),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_645),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_649),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_661),
.A2(n_524),
.B1(n_525),
.B2(n_521),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_600),
.A2(n_443),
.B1(n_386),
.B2(n_407),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_626),
.B(n_534),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_649),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_640),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_602),
.B(n_548),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_577),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_594),
.B(n_564),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_619),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_670),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_670),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_627),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_653),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_653),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_602),
.B(n_567),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_480),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_623),
.B(n_570),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_646),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_626),
.B(n_480),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_653),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_664),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_594),
.B(n_573),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_646),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_607),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_646),
.Y(n_750)
);

CKINVDCx16_ASAP7_75t_R g751 ( 
.A(n_609),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_630),
.B(n_538),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_664),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_664),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_635),
.B(n_539),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_663),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_637),
.B(n_545),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_577),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_663),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_589),
.A2(n_312),
.B1(n_314),
.B2(n_299),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_607),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_664),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_631),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_648),
.B(n_549),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_606),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_663),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_589),
.B(n_478),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_607),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_663),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_640),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_582),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_582),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_638),
.B(n_455),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_585),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_607),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_601),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_638),
.B(n_479),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_585),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_611),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_611),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_575),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_597),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_631),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_611),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_587),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_597),
.B(n_404),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_611),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_587),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_590),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_590),
.Y(n_793)
);

BUFx4f_ASAP7_75t_L g794 ( 
.A(n_581),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_575),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_610),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_597),
.B(n_483),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_657),
.B(n_516),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_593),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_593),
.Y(n_800)
);

BUFx4f_ASAP7_75t_L g801 ( 
.A(n_581),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_657),
.B(n_340),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_595),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_651),
.B(n_569),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_597),
.B(n_483),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_601),
.B(n_479),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_626),
.B(n_492),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_595),
.B(n_492),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_583),
.B(n_433),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_609),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_640),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_605),
.B(n_271),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_621),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_601),
.B(n_540),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_598),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_621),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_598),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_605),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_621),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_668),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_655),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_621),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_608),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_640),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_621),
.Y(n_828)
);

AO21x2_ASAP7_75t_L g829 ( 
.A1(n_669),
.A2(n_237),
.B(n_232),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_612),
.B(n_493),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_601),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_654),
.B(n_665),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_702),
.A2(n_642),
.B1(n_550),
.B2(n_666),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_786),
.A2(n_667),
.B1(n_491),
.B2(n_498),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_729),
.B(n_669),
.Y(n_835)
);

INVx6_ASAP7_75t_L g836 ( 
.A(n_797),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_581),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_780),
.B(n_581),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_681),
.B(n_511),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_678),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_798),
.B(n_655),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_737),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_737),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_702),
.A2(n_581),
.B1(n_629),
.B2(n_433),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_685),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_785),
.B(n_257),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_672),
.B(n_744),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_811),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_518),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_785),
.B(n_257),
.Y(n_850)
);

BUFx4f_ASAP7_75t_L g851 ( 
.A(n_789),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_731),
.B(n_497),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_740),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_744),
.A2(n_501),
.B1(n_389),
.B2(n_237),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_684),
.B(n_629),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_684),
.B(n_629),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_745),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_749),
.A2(n_239),
.B1(n_246),
.B2(n_232),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_794),
.B(n_801),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_794),
.A2(n_584),
.B(n_583),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_738),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_747),
.B(n_579),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_684),
.B(n_629),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_794),
.B(n_257),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_764),
.B(n_671),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_745),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_749),
.B(n_629),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_778),
.B(n_599),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_753),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_685),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_801),
.B(n_579),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_753),
.Y(n_872)
);

XNOR2xp5_ASAP7_75t_L g873 ( 
.A(n_714),
.B(n_579),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_801),
.B(n_238),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_754),
.A2(n_640),
.B1(n_246),
.B2(n_250),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_789),
.B(n_238),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_778),
.B(n_238),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_764),
.B(n_707),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_707),
.B(n_802),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_768),
.B(n_238),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_738),
.B(n_238),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_798),
.B(n_239),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_754),
.B(n_238),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_699),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_763),
.B(n_238),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_740),
.B(n_797),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_789),
.B(n_238),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_802),
.B(n_612),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_687),
.B(n_613),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_740),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_733),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_797),
.B(n_599),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_805),
.B(n_599),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_763),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_784),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_805),
.B(n_599),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_695),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_812),
.B(n_238),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_805),
.B(n_640),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_807),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_679),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_687),
.B(n_640),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_789),
.B(n_310),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_784),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_717),
.Y(n_905)
);

BUFx5_ASAP7_75t_L g906 ( 
.A(n_789),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_807),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_762),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_807),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_812),
.B(n_310),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_762),
.B(n_613),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_686),
.B(n_245),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_812),
.B(n_310),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_798),
.B(n_247),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_717),
.B(n_583),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_827),
.B(n_310),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_798),
.A2(n_250),
.B1(n_258),
.B2(n_253),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_699),
.A2(n_314),
.B1(n_315),
.B2(n_312),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_811),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_725),
.B(n_584),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_725),
.B(n_584),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_743),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_733),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_770),
.B(n_253),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_691),
.A2(n_620),
.B(n_591),
.Y(n_926)
);

AND2x6_ASAP7_75t_SL g927 ( 
.A(n_752),
.B(n_315),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_773),
.B(n_591),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_679),
.B(n_614),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_773),
.B(n_591),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_774),
.B(n_620),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_770),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_827),
.B(n_310),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_774),
.B(n_620),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_827),
.B(n_310),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_806),
.B(n_310),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_777),
.Y(n_937)
);

INVx8_ASAP7_75t_L g938 ( 
.A(n_789),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_789),
.A2(n_264),
.B1(n_280),
.B2(n_258),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_795),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_829),
.A2(n_280),
.B1(n_290),
.B2(n_264),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_829),
.A2(n_296),
.B1(n_309),
.B2(n_290),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_690),
.B(n_614),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_678),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_777),
.B(n_622),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_678),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_689),
.B(n_249),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_814),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_781),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_829),
.A2(n_309),
.B1(n_313),
.B2(n_296),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_795),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_695),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_698),
.B(n_256),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_809),
.B(n_310),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_678),
.A2(n_321),
.B1(n_358),
.B2(n_313),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_781),
.B(n_622),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_788),
.B(n_622),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_736),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_788),
.B(n_624),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_675),
.B(n_310),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_L g961 ( 
.A(n_809),
.B(n_675),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_791),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_791),
.B(n_624),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_676),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_688),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_675),
.B(n_321),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_792),
.B(n_624),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_792),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_793),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_793),
.A2(n_373),
.B1(n_392),
.B2(n_358),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_703),
.B(n_259),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_690),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_704),
.B(n_261),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_799),
.B(n_578),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_799),
.B(n_578),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_373),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_800),
.B(n_392),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_803),
.A2(n_417),
.B1(n_424),
.B2(n_403),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_803),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_688),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_701),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_814),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_824),
.B(n_615),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_817),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_736),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_741),
.B(n_776),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_817),
.B(n_403),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_675),
.B(n_417),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_819),
.B(n_424),
.Y(n_989)
);

AND2x6_ASAP7_75t_L g990 ( 
.A(n_779),
.B(n_831),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_819),
.B(n_430),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_820),
.B(n_430),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_701),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_820),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_675),
.B(n_432),
.Y(n_995)
);

AO21x2_ASAP7_75t_L g996 ( 
.A1(n_767),
.A2(n_432),
.B(n_551),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_826),
.B(n_615),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_826),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_776),
.B(n_262),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_691),
.A2(n_662),
.B1(n_660),
.B2(n_659),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_767),
.B(n_618),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_769),
.B(n_618),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_706),
.B(n_266),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_769),
.B(n_632),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_771),
.B(n_632),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_771),
.B(n_636),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_808),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_742),
.B(n_636),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_832),
.B(n_319),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_865),
.B(n_720),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_835),
.B(n_694),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_855),
.A2(n_677),
.B(n_676),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_857),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_857),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_866),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_906),
.B(n_675),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_SL g1017 ( 
.A(n_854),
.B(n_723),
.C(n_821),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_845),
.B(n_694),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_866),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_938),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_869),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_884),
.B(n_808),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_869),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_845),
.B(n_694),
.Y(n_1024)
);

BUFx5_ASAP7_75t_L g1025 ( 
.A(n_842),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_878),
.B(n_733),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_872),
.Y(n_1027)
);

CKINVDCx11_ASAP7_75t_R g1028 ( 
.A(n_924),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_SL g1029 ( 
.A(n_859),
.B(n_870),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_870),
.B(n_694),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_872),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_894),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_905),
.B(n_830),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_SL g1034 ( 
.A(n_1003),
.B(n_724),
.C(n_824),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_901),
.B(n_751),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_894),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_905),
.B(n_830),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_884),
.B(n_779),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_900),
.A2(n_680),
.B1(n_692),
.B2(n_674),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_895),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_907),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_848),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_909),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_912),
.A2(n_680),
.B1(n_692),
.B2(n_674),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_911),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_911),
.Y(n_1047)
);

BUFx10_ASAP7_75t_L g1048 ( 
.A(n_891),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_944),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_911),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_895),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_889),
.B(n_742),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_834),
.B(n_751),
.C(n_714),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_958),
.B(n_831),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_937),
.B(n_746),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_958),
.B(n_853),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_904),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_904),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_920),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_924),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_860),
.A2(n_746),
.B(n_730),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_940),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_940),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_949),
.B(n_761),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_941),
.A2(n_696),
.B1(n_697),
.B2(n_693),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_847),
.A2(n_816),
.B1(n_757),
.B2(n_765),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_985),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_962),
.B(n_693),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_888),
.B(n_821),
.Y(n_1069)
);

OR2x6_ASAP7_75t_L g1070 ( 
.A(n_938),
.B(n_804),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_838),
.B(n_696),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_944),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_840),
.B(n_728),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_999),
.B(n_755),
.C(n_766),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_SL g1075 ( 
.A(n_833),
.B(n_796),
.C(n_766),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_972),
.B(n_712),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_948),
.B(n_823),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_861),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_951),
.Y(n_1079)
);

NOR2x2_ASAP7_75t_L g1080 ( 
.A(n_882),
.B(n_796),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_906),
.B(n_728),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_951),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_890),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_983),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_965),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_968),
.B(n_697),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_969),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_861),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_944),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_861),
.B(n_644),
.Y(n_1090)
);

INVx6_ASAP7_75t_L g1091 ( 
.A(n_861),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_982),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_879),
.B(n_644),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_979),
.B(n_700),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_836),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_946),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_984),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_891),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_994),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_998),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_897),
.B(n_268),
.C(n_267),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1008),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_943),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1007),
.B(n_700),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_886),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_916),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_897),
.B(n_274),
.C(n_270),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_965),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_908),
.B(n_647),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_923),
.B(n_705),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1001),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_837),
.B(n_705),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_908),
.B(n_932),
.Y(n_1113)
);

BUFx8_ASAP7_75t_L g1114 ( 
.A(n_891),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_986),
.A2(n_716),
.B1(n_719),
.B2(n_711),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1002),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_839),
.B(n_234),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1004),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_952),
.B(n_277),
.C(n_276),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_929),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_847),
.B(n_708),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_980),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_836),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_980),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_841),
.Y(n_1125)
);

BUFx8_ASAP7_75t_L g1126 ( 
.A(n_990),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_906),
.B(n_851),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_862),
.B(n_711),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_871),
.A2(n_719),
.B1(n_721),
.B2(n_716),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_836),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_932),
.B(n_721),
.Y(n_1132)
);

INVx3_ASAP7_75t_SL g1133 ( 
.A(n_952),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_849),
.B(n_647),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_852),
.B(n_350),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_938),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_841),
.B(n_650),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_908),
.B(n_650),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_871),
.B(n_357),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_908),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_990),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_938),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_946),
.B(n_658),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_914),
.B(n_418),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_990),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_851),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_946),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_925),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_840),
.B(n_658),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_981),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_981),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_873),
.Y(n_1153)
);

BUFx8_ASAP7_75t_L g1154 ( 
.A(n_990),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_997),
.B(n_722),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_947),
.B(n_953),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_915),
.B(n_722),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_928),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_867),
.B(n_727),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_840),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_927),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_L g1162 ( 
.A(n_841),
.B(n_420),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_841),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_906),
.B(n_728),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_906),
.B(n_728),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_993),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_930),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_931),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1009),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_882),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_934),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_942),
.A2(n_732),
.B1(n_734),
.B2(n_727),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_950),
.A2(n_734),
.B1(n_732),
.B2(n_709),
.Y(n_1173)
);

INVx3_ASAP7_75t_SL g1174 ( 
.A(n_1009),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_851),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_918),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1009),
.B(n_659),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_971),
.A2(n_322),
.B(n_324),
.C(n_319),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_993),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_SL g1180 ( 
.A(n_973),
.B(n_288),
.C(n_285),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_921),
.B(n_708),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_906),
.B(n_728),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_945),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_906),
.B(n_728),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_902),
.B(n_772),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_990),
.B(n_876),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_922),
.B(n_709),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_859),
.B(n_772),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1000),
.B(n_710),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_856),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_990),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1009),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_882),
.B(n_660),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_956),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_882),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_925),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_863),
.B(n_710),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_957),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_964),
.Y(n_1199)
);

INVx3_ASAP7_75t_SL g1200 ( 
.A(n_881),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_964),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_881),
.B(n_662),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_959),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_919),
.B(n_301),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_964),
.B(n_899),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1156),
.A2(n_936),
.B(n_864),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_1201),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1112),
.A2(n_864),
.B(n_874),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1061),
.A2(n_874),
.B(n_844),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1156),
.B(n_974),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1190),
.A2(n_877),
.B(n_936),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1015),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1190),
.A2(n_877),
.B(n_898),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1011),
.A2(n_939),
.B1(n_893),
.B2(n_896),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1134),
.B(n_975),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1111),
.B(n_976),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1061),
.A2(n_885),
.B(n_883),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1197),
.A2(n_910),
.B(n_898),
.Y(n_1218)
);

AND3x2_ASAP7_75t_L g1219 ( 
.A(n_1135),
.B(n_324),
.C(n_322),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1117),
.A2(n_885),
.B1(n_883),
.B2(n_892),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1160),
.A2(n_903),
.B(n_887),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1019),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1012),
.A2(n_967),
.B(n_963),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1188),
.A2(n_1205),
.B(n_1160),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1199),
.A2(n_903),
.B(n_961),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1069),
.B(n_996),
.Y(n_1226)
);

BUFx4_ASAP7_75t_SL g1227 ( 
.A(n_1043),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1116),
.A2(n_868),
.B1(n_858),
.B2(n_846),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1188),
.A2(n_926),
.B(n_880),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1069),
.B(n_996),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1127),
.A2(n_880),
.B(n_910),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1199),
.A2(n_961),
.B(n_677),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1178),
.A2(n_955),
.A3(n_987),
.B(n_977),
.Y(n_1233)
);

AO21x1_ASAP7_75t_L g1234 ( 
.A1(n_1029),
.A2(n_991),
.B(n_989),
.Y(n_1234)
);

NOR2xp67_ASAP7_75t_L g1235 ( 
.A(n_1074),
.B(n_992),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1178),
.A2(n_726),
.A3(n_735),
.B(n_718),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1059),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1127),
.A2(n_917),
.B(n_913),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1010),
.A2(n_1024),
.A3(n_1030),
.B(n_1018),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1025),
.B(n_913),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1121),
.A2(n_933),
.B(n_917),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1133),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1133),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1121),
.A2(n_935),
.B(n_933),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1199),
.A2(n_677),
.B(n_676),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1205),
.A2(n_935),
.B(n_850),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1118),
.A2(n_846),
.B1(n_850),
.B2(n_970),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1201),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1025),
.B(n_748),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1073),
.A2(n_1136),
.B(n_1020),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1185),
.A2(n_960),
.B(n_730),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1185),
.A2(n_1187),
.B(n_1181),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1117),
.A2(n_978),
.B(n_425),
.Y(n_1253)
);

AOI221xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1010),
.A2(n_352),
.B1(n_431),
.B2(n_394),
.C(n_387),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1139),
.A2(n_988),
.B1(n_995),
.B2(n_966),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1131),
.B(n_1145),
.Y(n_1256)
);

BUFx5_ASAP7_75t_L g1257 ( 
.A(n_1141),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1144),
.B(n_966),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1055),
.A2(n_730),
.B(n_713),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1093),
.B(n_718),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1028),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1088),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_758),
.B(n_713),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1019),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1029),
.A2(n_1128),
.B(n_1066),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1102),
.B(n_726),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1129),
.A2(n_960),
.B(n_758),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1105),
.A2(n_1200),
.B1(n_1175),
.B2(n_1147),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1033),
.B(n_1037),
.Y(n_1269)
);

NAND2x1_ASAP7_75t_L g1270 ( 
.A(n_1201),
.B(n_713),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1179),
.A2(n_782),
.B(n_758),
.Y(n_1271)
);

AOI31xp67_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_735),
.A3(n_988),
.B(n_995),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1046),
.B(n_782),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1021),
.A2(n_790),
.B(n_782),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1028),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1158),
.B(n_875),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1139),
.A2(n_368),
.B(n_449),
.C(n_431),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1021),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1023),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1167),
.B(n_1168),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1088),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1073),
.A2(n_750),
.B(n_748),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1201),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1060),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1092),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1171),
.B(n_790),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1020),
.A2(n_750),
.B(n_748),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1183),
.B(n_790),
.Y(n_1288)
);

AO22x2_ASAP7_75t_L g1289 ( 
.A1(n_1017),
.A2(n_1075),
.B1(n_1204),
.B2(n_1137),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1157),
.A2(n_327),
.A3(n_341),
.B(n_449),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1103),
.B(n_493),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1159),
.A2(n_954),
.B(n_756),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1179),
.A2(n_815),
.B(n_810),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1023),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1085),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1020),
.A2(n_756),
.B(n_750),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1020),
.A2(n_759),
.B(n_756),
.Y(n_1297)
);

OA22x2_ASAP7_75t_L g1298 ( 
.A1(n_1120),
.A2(n_327),
.B1(n_341),
.B2(n_343),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1013),
.A2(n_343),
.A3(n_352),
.B(n_394),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_1020),
.B(n_759),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1014),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1085),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1084),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1194),
.B(n_810),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1068),
.A2(n_815),
.B(n_810),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1025),
.B(n_759),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1088),
.Y(n_1307)
);

OAI22x1_ASAP7_75t_L g1308 ( 
.A1(n_1144),
.A2(n_306),
.B1(n_297),
.B2(n_303),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1136),
.B(n_760),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1060),
.B(n_359),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1049),
.A2(n_818),
.B(n_815),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1049),
.A2(n_1089),
.B(n_1072),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1159),
.A2(n_954),
.B(n_760),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1026),
.B(n_301),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1193),
.A2(n_809),
.B(n_302),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1035),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1176),
.A2(n_760),
.B1(n_825),
.B2(n_818),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1049),
.A2(n_825),
.B(n_818),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1203),
.B(n_825),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1041),
.B(n_311),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1027),
.A2(n_359),
.A3(n_367),
.B(n_368),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1149),
.A2(n_377),
.B(n_367),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1086),
.A2(n_495),
.B(n_494),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1198),
.B(n_320),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1094),
.A2(n_495),
.B(n_494),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1040),
.A2(n_503),
.B(n_496),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1040),
.A2(n_503),
.B(n_496),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1087),
.A2(n_387),
.B(n_377),
.C(n_381),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1159),
.A2(n_809),
.B(n_772),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_L g1330 ( 
.A(n_1186),
.B(n_772),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1198),
.B(n_325),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1058),
.A2(n_508),
.B(n_507),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1077),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1058),
.A2(n_508),
.B(n_507),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1177),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1114),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1136),
.A2(n_772),
.B(n_683),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_772),
.B(n_683),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1022),
.B(n_301),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_1076),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1100),
.B(n_326),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1136),
.A2(n_683),
.B(n_673),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1072),
.A2(n_515),
.B(n_514),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1108),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1067),
.Y(n_1346)
);

O2A1O1Ixp5_ASAP7_75t_L g1347 ( 
.A1(n_1155),
.A2(n_522),
.B(n_514),
.C(n_515),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1106),
.B(n_328),
.Y(n_1348)
);

O2A1O1Ixp5_ASAP7_75t_L g1349 ( 
.A1(n_1031),
.A2(n_517),
.B(n_522),
.C(n_381),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1072),
.A2(n_517),
.B(n_809),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_1048),
.Y(n_1351)
);

OA22x2_ASAP7_75t_L g1352 ( 
.A1(n_1169),
.A2(n_1192),
.B1(n_1174),
.B2(n_1195),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1022),
.B(n_331),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_SL g1354 ( 
.A1(n_1149),
.A2(n_809),
.B(n_113),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1176),
.A2(n_809),
.B1(n_302),
.B2(n_813),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1032),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1036),
.A2(n_12),
.A3(n_16),
.B(n_17),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1051),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1132),
.A2(n_683),
.B(n_673),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1079),
.A2(n_683),
.B(n_673),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1070),
.B(n_673),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1159),
.A2(n_1071),
.B(n_1052),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1079),
.A2(n_715),
.B(n_673),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1057),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1200),
.A2(n_828),
.B1(n_822),
.B2(n_813),
.Y(n_1365)
);

AOI211x1_ASAP7_75t_L g1366 ( 
.A1(n_1064),
.A2(n_384),
.B(n_308),
.C(n_316),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1108),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1025),
.B(n_828),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1089),
.A2(n_1148),
.B(n_1096),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1022),
.B(n_332),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1189),
.A2(n_12),
.A3(n_16),
.B(n_18),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1088),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1122),
.A2(n_828),
.B(n_822),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1076),
.B(n_334),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1360),
.A2(n_1045),
.B(n_1122),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1207),
.B(n_1142),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1212),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1362),
.A2(n_1104),
.B(n_1110),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1210),
.B(n_1196),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1239),
.B(n_1090),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1258),
.A2(n_1202),
.B(n_1143),
.Y(n_1382)
);

OAI221xp5_ASAP7_75t_L g1383 ( 
.A1(n_1253),
.A2(n_1034),
.B1(n_1162),
.B2(n_1180),
.C(n_1053),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1212),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1222),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1258),
.A2(n_1153),
.B1(n_1070),
.B2(n_1125),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1222),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1359),
.A2(n_1265),
.B(n_1234),
.Y(n_1388)
);

OAI222xp33_ASAP7_75t_L g1389 ( 
.A1(n_1256),
.A2(n_1070),
.B1(n_1042),
.B2(n_1044),
.C1(n_1083),
.C2(n_1170),
.Y(n_1389)
);

AOI31xp67_ASAP7_75t_L g1390 ( 
.A1(n_1220),
.A2(n_1152),
.A3(n_1124),
.B(n_1151),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1206),
.A2(n_1277),
.A3(n_1214),
.B(n_1247),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1323),
.A2(n_1172),
.B(n_1065),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1360),
.A2(n_1151),
.B(n_1124),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1207),
.B(n_1142),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1363),
.A2(n_1166),
.B(n_1152),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1242),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1289),
.A2(n_1153),
.B1(n_1070),
.B2(n_1163),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1275),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1264),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1363),
.A2(n_1166),
.B(n_1063),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1351),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1323),
.A2(n_1173),
.B(n_1082),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1305),
.A2(n_1186),
.B(n_1062),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1373),
.A2(n_1096),
.B(n_1089),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1373),
.A2(n_1148),
.B(n_1096),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1207),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1239),
.B(n_1090),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1215),
.B(n_1056),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1341),
.B(n_1056),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1305),
.A2(n_1274),
.B(n_1259),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1264),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1334),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1280),
.B(n_1056),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1216),
.A2(n_1147),
.B1(n_1175),
.B2(n_1050),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1207),
.Y(n_1416)
);

NAND2x1_ASAP7_75t_L g1417 ( 
.A(n_1361),
.B(n_1142),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_SL g1418 ( 
.A1(n_1277),
.A2(n_1047),
.B(n_1081),
.C(n_1016),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1278),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1237),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1269),
.B(n_1226),
.Y(n_1421)
);

INVx4_ASAP7_75t_SL g1422 ( 
.A(n_1361),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1274),
.A2(n_1148),
.B(n_1039),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1230),
.B(n_1090),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1228),
.A2(n_1071),
.A3(n_1159),
.B(n_1025),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1341),
.B(n_1174),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1224),
.A2(n_1223),
.B(n_1312),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1268),
.A2(n_1147),
.B1(n_1175),
.B2(n_1113),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1341),
.B(n_1067),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1325),
.A2(n_1202),
.B(n_1138),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1325),
.A2(n_1138),
.B(n_1109),
.Y(n_1431)
);

INVx8_ASAP7_75t_L g1432 ( 
.A(n_1361),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1278),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1295),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1295),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1316),
.B(n_1193),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1289),
.A2(n_1193),
.B1(n_1138),
.B2(n_1109),
.Y(n_1437)
);

INVx3_ASAP7_75t_SL g1438 ( 
.A(n_1243),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1235),
.A2(n_1202),
.B(n_1143),
.C(n_1109),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1276),
.A2(n_1175),
.B1(n_1147),
.B2(n_1113),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1369),
.A2(n_1081),
.B(n_1016),
.Y(n_1441)
);

AO31x2_ASAP7_75t_L g1442 ( 
.A1(n_1328),
.A2(n_1071),
.A3(n_1159),
.B(n_1025),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1324),
.B(n_1095),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1302),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1302),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_SL g1446 ( 
.A1(n_1354),
.A2(n_1130),
.B(n_1123),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1292),
.A2(n_1119),
.B(n_1107),
.C(n_1101),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1217),
.A2(n_1165),
.B(n_1164),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1241),
.A2(n_1143),
.B(n_1150),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1217),
.A2(n_1271),
.B(n_1263),
.Y(n_1450)
);

CKINVDCx8_ASAP7_75t_R g1451 ( 
.A(n_1243),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1345),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1285),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1345),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1331),
.B(n_1095),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1244),
.A2(n_1150),
.B(n_1071),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1293),
.A2(n_1165),
.B(n_1164),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1257),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1313),
.A2(n_1130),
.B(n_1123),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1367),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1219),
.B(n_1114),
.C(n_1054),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1209),
.A2(n_1184),
.B(n_1182),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1275),
.Y(n_1463)
);

BUFx8_ASAP7_75t_L g1464 ( 
.A(n_1351),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1337),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_R g1466 ( 
.A(n_1261),
.B(n_1161),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1367),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1336),
.B(n_1113),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1333),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1227),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1358),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1209),
.A2(n_1184),
.B(n_1182),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1311),
.A2(n_1071),
.B(n_1025),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1336),
.B(n_1078),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1364),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1318),
.A2(n_1071),
.B(n_1126),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1229),
.A2(n_1327),
.B(n_1326),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1289),
.A2(n_1038),
.B1(n_1054),
.B2(n_1078),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1374),
.A2(n_422),
.B1(n_364),
.B2(n_366),
.C(n_369),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1229),
.A2(n_1154),
.B(n_1126),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1330),
.A2(n_1150),
.B(n_1142),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1326),
.A2(n_1154),
.B(n_1126),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1255),
.A2(n_1146),
.B(n_1141),
.C(n_1038),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1262),
.Y(n_1484)
);

O2A1O1Ixp5_ASAP7_75t_L g1485 ( 
.A1(n_1208),
.A2(n_1054),
.B(n_1038),
.C(n_1080),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1227),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1327),
.A2(n_1191),
.B(n_1154),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1279),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1337),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1294),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1266),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1317),
.A2(n_1146),
.B1(n_1091),
.B2(n_1140),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1332),
.A2(n_1191),
.B(n_1140),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1257),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1257),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1352),
.B(n_1140),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1291),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1332),
.A2(n_1191),
.B(n_1140),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1346),
.B(n_1048),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1335),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1314),
.B(n_1161),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1301),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1251),
.A2(n_1091),
.B(n_1080),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1261),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1257),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1251),
.A2(n_1091),
.B(n_1048),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1356),
.A2(n_405),
.B1(n_339),
.B2(n_342),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1239),
.B(n_335),
.Y(n_1508)
);

AO32x2_ASAP7_75t_L g1509 ( 
.A1(n_1254),
.A2(n_1114),
.A3(n_384),
.B1(n_317),
.B2(n_316),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1213),
.A2(n_408),
.B(n_337),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1252),
.A2(n_379),
.B(n_378),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1315),
.A2(n_1098),
.B(n_822),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1308),
.A2(n_302),
.B1(n_1098),
.B2(n_308),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_SL g1514 ( 
.A(n_1284),
.B(n_1098),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1260),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1286),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1288),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1252),
.A2(n_414),
.B(n_344),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1344),
.A2(n_813),
.B(n_787),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1219),
.B(n_411),
.C(n_345),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1340),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1273),
.B(n_110),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1299),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1304),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1319),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1257),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1328),
.A2(n_1221),
.A3(n_1225),
.B(n_1365),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1352),
.A2(n_302),
.B1(n_308),
.B2(n_316),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1211),
.A2(n_419),
.B(n_353),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1273),
.B(n_116),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1239),
.B(n_308),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1353),
.A2(n_426),
.B1(n_355),
.B2(n_356),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1299),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1370),
.A2(n_316),
.B1(n_317),
.B2(n_384),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1273),
.A2(n_317),
.B1(n_384),
.B2(n_436),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1349),
.A2(n_438),
.B(n_380),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1262),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1298),
.A2(n_1348),
.B1(n_1320),
.B2(n_1342),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1246),
.A2(n_813),
.B(n_787),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_R g1540 ( 
.A(n_1284),
.B(n_362),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1299),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1299),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1246),
.A2(n_822),
.B(n_813),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1368),
.A2(n_822),
.B(n_787),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1368),
.A2(n_787),
.B(n_783),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1310),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1355),
.B(n_382),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1236),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1350),
.A2(n_1267),
.B(n_1231),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1267),
.A2(n_783),
.B(n_775),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1231),
.A2(n_783),
.B(n_775),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1233),
.B(n_317),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1349),
.A2(n_439),
.B(n_388),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1250),
.A2(n_787),
.B(n_783),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1236),
.Y(n_1555)
);

AOI22x1_ASAP7_75t_L g1556 ( 
.A1(n_1218),
.A2(n_437),
.B1(n_397),
.B2(n_398),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1238),
.A2(n_783),
.B(n_775),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1497),
.B(n_1290),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1384),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1398),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1479),
.A2(n_1534),
.B1(n_1383),
.B2(n_1513),
.C(n_1510),
.Y(n_1561)
);

NAND2xp33_ASAP7_75t_R g1562 ( 
.A(n_1426),
.B(n_1248),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1406),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_R g1564 ( 
.A(n_1381),
.B(n_1248),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1421),
.B(n_1290),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1384),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1413),
.B(n_1298),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1380),
.B(n_1366),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1436),
.B(n_1321),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1406),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1502),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1407),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1521),
.B(n_1321),
.Y(n_1573)
);

OR2x6_ASAP7_75t_SL g1574 ( 
.A(n_1504),
.B(n_385),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1381),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_R g1576 ( 
.A(n_1408),
.B(n_1283),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1386),
.A2(n_1240),
.B1(n_1283),
.B2(n_1310),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1407),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1409),
.A2(n_1310),
.B1(n_413),
.B2(n_427),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1408),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1508),
.B(n_1290),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1398),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1414),
.B(n_1290),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1529),
.A2(n_401),
.B1(n_440),
.B2(n_441),
.C(n_445),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1407),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1424),
.B(n_1240),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1502),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1474),
.B(n_1321),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1515),
.B(n_1307),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1501),
.A2(n_444),
.B1(n_1257),
.B2(n_1307),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1397),
.A2(n_1372),
.B1(n_1262),
.B2(n_1281),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1474),
.B(n_1321),
.Y(n_1592)
);

AO221x2_ASAP7_75t_L g1593 ( 
.A1(n_1389),
.A2(n_1371),
.B1(n_1357),
.B2(n_26),
.C(n_29),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1481),
.A2(n_1306),
.B(n_1249),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1382),
.B(n_1249),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1483),
.A2(n_1306),
.B(n_1232),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1471),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1531),
.A2(n_1322),
.B1(n_1238),
.B2(n_1372),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1385),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1538),
.A2(n_1372),
.B1(n_1281),
.B2(n_1262),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1385),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1474),
.B(n_1357),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1420),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1475),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1429),
.B(n_1281),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1420),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1508),
.B(n_1233),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1478),
.A2(n_1372),
.B1(n_1281),
.B2(n_1309),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1437),
.A2(n_1309),
.B1(n_1300),
.B2(n_1270),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1531),
.A2(n_1371),
.B1(n_1329),
.B2(n_1357),
.Y(n_1610)
);

BUFx8_ASAP7_75t_SL g1611 ( 
.A(n_1463),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1469),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1547),
.A2(n_1300),
.B1(n_1343),
.B2(n_1245),
.Y(n_1613)
);

NAND3x1_ASAP7_75t_L g1614 ( 
.A(n_1532),
.B(n_22),
.C(n_24),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_SL g1615 ( 
.A(n_1451),
.B(n_1338),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1535),
.A2(n_1347),
.B1(n_1282),
.B2(n_1287),
.C(n_1297),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1477),
.A2(n_1347),
.B(n_1272),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1443),
.A2(n_1296),
.B1(n_1339),
.B2(n_1233),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1455),
.A2(n_1233),
.B1(n_775),
.B2(n_715),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1439),
.A2(n_1236),
.B(n_1371),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1488),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1552),
.A2(n_1371),
.B1(n_1357),
.B2(n_31),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1453),
.A2(n_1468),
.B1(n_1515),
.B2(n_1451),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1432),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1522),
.B(n_1236),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1507),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.C(n_32),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1463),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1488),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1453),
.A2(n_775),
.B1(n_715),
.B2(n_37),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1552),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1432),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1490),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1465),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1490),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1377),
.B(n_118),
.Y(n_1635)
);

AOI21xp33_ASAP7_75t_L g1636 ( 
.A1(n_1556),
.A2(n_34),
.B(n_38),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1461),
.A2(n_1514),
.B1(n_1546),
.B2(n_1496),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1528),
.A2(n_1491),
.B1(n_1449),
.B2(n_1415),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1546),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1378),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1410),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1432),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1399),
.Y(n_1643)
);

AO31x2_ASAP7_75t_L g1644 ( 
.A1(n_1523),
.A2(n_41),
.A3(n_42),
.B(n_45),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1378),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1377),
.B(n_227),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1388),
.A2(n_225),
.B(n_219),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1387),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1396),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1556),
.A2(n_1491),
.B1(n_1520),
.B2(n_1516),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1484),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1522),
.B(n_47),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_R g1653 ( 
.A(n_1504),
.B(n_215),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1522),
.B(n_47),
.Y(n_1654)
);

OAI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1496),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1516),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1438),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1456),
.A2(n_55),
.B(n_57),
.C(n_58),
.Y(n_1658)
);

INVx3_ASAP7_75t_SL g1659 ( 
.A(n_1438),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1396),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1489),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1485),
.A2(n_1440),
.B(n_1517),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1422),
.B(n_214),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1388),
.A2(n_1459),
.B(n_1446),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1442),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1387),
.B(n_64),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1517),
.A2(n_66),
.B1(n_69),
.B2(n_74),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1524),
.B(n_77),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1524),
.B(n_77),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1477),
.A2(n_123),
.B(n_202),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1537),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1465),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1525),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1530),
.B(n_79),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_1470),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1530),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1496),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1399),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1525),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1412),
.B(n_90),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1496),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1530),
.A2(n_1447),
.B(n_1432),
.C(n_1503),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1484),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1428),
.A2(n_1492),
.B1(n_1499),
.B2(n_1416),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_R g1685 ( 
.A(n_1392),
.B(n_1458),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1486),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1489),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1509),
.B(n_99),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1379),
.A2(n_100),
.B1(n_103),
.B2(n_105),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1418),
.A2(n_100),
.B1(n_105),
.B2(n_119),
.C(n_127),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1484),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1433),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1533),
.B(n_130),
.C(n_132),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1541),
.B(n_135),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1379),
.A2(n_195),
.B1(n_146),
.B2(n_149),
.Y(n_1695)
);

OAI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1542),
.A2(n_139),
.B(n_153),
.C(n_156),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1417),
.A2(n_163),
.B1(n_170),
.B2(n_174),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1416),
.B(n_1417),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1484),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1379),
.A2(n_175),
.B1(n_192),
.B2(n_1433),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1503),
.A2(n_1434),
.B(n_1444),
.C(n_1454),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1537),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1412),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1434),
.B(n_1444),
.Y(n_1704)
);

AOI222xp33_ASAP7_75t_L g1705 ( 
.A1(n_1466),
.A2(n_1540),
.B1(n_1464),
.B2(n_1401),
.C1(n_1422),
.C2(n_1445),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1419),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1445),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1401),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1452),
.B(n_1454),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1484),
.Y(n_1710)
);

BUFx12f_ASAP7_75t_L g1711 ( 
.A(n_1401),
.Y(n_1711)
);

CKINVDCx11_ASAP7_75t_R g1712 ( 
.A(n_1464),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1419),
.B(n_1435),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1550),
.A2(n_1411),
.B(n_1539),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_SL g1715 ( 
.A(n_1464),
.B(n_1376),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1452),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1480),
.B(n_1459),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1435),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1376),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1720)
);

OAI222xp33_ASAP7_75t_L g1721 ( 
.A1(n_1460),
.A2(n_1467),
.B1(n_1376),
.B2(n_1394),
.C1(n_1555),
.C2(n_1548),
.Y(n_1721)
);

NAND2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1458),
.B(n_1526),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1509),
.B(n_1422),
.Y(n_1723)
);

CKINVDCx11_ASAP7_75t_R g1724 ( 
.A(n_1422),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1394),
.A2(n_1526),
.B1(n_1495),
.B2(n_1458),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1392),
.A2(n_1555),
.B1(n_1553),
.B2(n_1536),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1393),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1391),
.B(n_1425),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1509),
.B(n_1391),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1509),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1480),
.B(n_1482),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1509),
.B(n_1391),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1400),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1511),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1391),
.B(n_1442),
.Y(n_1735)
);

CKINVDCx16_ASAP7_75t_R g1736 ( 
.A(n_1431),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1392),
.A2(n_1494),
.B1(n_1505),
.B2(n_1495),
.Y(n_1737)
);

BUFx4f_ASAP7_75t_L g1738 ( 
.A(n_1394),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1494),
.A2(n_1495),
.B1(n_1526),
.B2(n_1505),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1391),
.B(n_1442),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1494),
.A2(n_1505),
.B1(n_1402),
.B2(n_1430),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1402),
.A2(n_1430),
.B1(n_1511),
.B2(n_1518),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1536),
.A2(n_1553),
.B1(n_1446),
.B2(n_1402),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1487),
.Y(n_1745)
);

NAND3x1_ASAP7_75t_L g1746 ( 
.A(n_1544),
.B(n_1442),
.C(n_1487),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_SL g1747 ( 
.A(n_1545),
.B(n_1431),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1493),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1400),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1393),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1425),
.B(n_1527),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1430),
.A2(n_1511),
.B1(n_1518),
.B2(n_1553),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1473),
.B(n_1506),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1425),
.B(n_1518),
.Y(n_1754)
);

BUFx4f_ASAP7_75t_SL g1755 ( 
.A(n_1711),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1724),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1561),
.B(n_1536),
.C(n_1500),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1590),
.A2(n_1425),
.B1(n_1527),
.B2(n_1390),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1575),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1579),
.A2(n_1431),
.B1(n_1512),
.B2(n_1498),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1575),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1694),
.A2(n_1403),
.B1(n_1512),
.B2(n_1545),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1579),
.B(n_1498),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1694),
.A2(n_1403),
.B1(n_1545),
.B2(n_1473),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1611),
.Y(n_1765)
);

CKINVDCx20_ASAP7_75t_R g1766 ( 
.A(n_1687),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1626),
.A2(n_1375),
.B1(n_1423),
.B2(n_1549),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1593),
.A2(n_1681),
.B1(n_1677),
.B2(n_1638),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1587),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1630),
.A2(n_1493),
.B1(n_1423),
.B2(n_1375),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1675),
.A2(n_1527),
.B1(n_1476),
.B2(n_1472),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1630),
.A2(n_1441),
.B1(n_1472),
.B2(n_1462),
.Y(n_1772)
);

OAI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1639),
.A2(n_1527),
.B1(n_1462),
.B2(n_1441),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1686),
.A2(n_1527),
.B1(n_1427),
.B2(n_1550),
.C(n_1448),
.Y(n_1774)
);

OR2x6_ASAP7_75t_L g1775 ( 
.A(n_1698),
.B(n_1427),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1661),
.A2(n_1448),
.B1(n_1395),
.B2(n_1551),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1593),
.A2(n_1551),
.B1(n_1557),
.B2(n_1543),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1675),
.A2(n_1457),
.B1(n_1404),
.B2(n_1405),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1569),
.B(n_1404),
.Y(n_1779)
);

BUFx10_ASAP7_75t_L g1780 ( 
.A(n_1633),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1570),
.B(n_1405),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1624),
.B(n_1557),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1586),
.B(n_1457),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1621),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1650),
.A2(n_1539),
.B(n_1543),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1623),
.A2(n_1554),
.B1(n_1519),
.B2(n_1450),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1686),
.A2(n_1395),
.B1(n_1450),
.B2(n_1519),
.C(n_1639),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1658),
.A2(n_1689),
.B(n_1584),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1593),
.A2(n_1688),
.B1(n_1653),
.B2(n_1577),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1658),
.A2(n_1676),
.B1(n_1689),
.B2(n_1667),
.C(n_1679),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1742),
.A2(n_1620),
.B(n_1753),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1636),
.A2(n_1655),
.B1(n_1690),
.B2(n_1656),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1586),
.B(n_1567),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1668),
.B(n_1669),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1650),
.A2(n_1660),
.B1(n_1637),
.B2(n_1606),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1655),
.A2(n_1673),
.B1(n_1679),
.B2(n_1667),
.Y(n_1796)
);

AOI222xp33_ASAP7_75t_L g1797 ( 
.A1(n_1656),
.A2(n_1673),
.B1(n_1695),
.B2(n_1652),
.C1(n_1654),
.C2(n_1674),
.Y(n_1797)
);

BUFx4f_ASAP7_75t_SL g1798 ( 
.A(n_1560),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1628),
.Y(n_1799)
);

OAI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1641),
.A2(n_1622),
.B(n_1695),
.C(n_1700),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1568),
.A2(n_1700),
.B1(n_1595),
.B2(n_1573),
.Y(n_1801)
);

INVx4_ASAP7_75t_L g1802 ( 
.A(n_1659),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1632),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1622),
.A2(n_1629),
.B1(n_1591),
.B2(n_1729),
.C(n_1732),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1581),
.A2(n_1565),
.B(n_1583),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1637),
.A2(n_1603),
.B1(n_1682),
.B2(n_1614),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1595),
.A2(n_1591),
.B1(n_1684),
.B2(n_1588),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1682),
.A2(n_1659),
.B1(n_1657),
.B2(n_1563),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1653),
.A2(n_1696),
.B1(n_1600),
.B2(n_1663),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1592),
.B(n_1602),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1612),
.A2(n_1649),
.B1(n_1558),
.B2(n_1738),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1671),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1705),
.A2(n_1604),
.B1(n_1597),
.B2(n_1666),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1589),
.B(n_1716),
.Y(n_1814)
);

BUFx8_ASAP7_75t_SL g1815 ( 
.A(n_1582),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1712),
.A2(n_1607),
.B1(n_1662),
.B2(n_1663),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1671),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1564),
.A2(n_1576),
.B1(n_1736),
.B2(n_1615),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1562),
.A2(n_1715),
.B1(n_1635),
.B2(n_1646),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_1672),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1738),
.A2(n_1693),
.B1(n_1598),
.B2(n_1605),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1580),
.B(n_1634),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1625),
.A2(n_1723),
.B1(n_1646),
.B2(n_1635),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1693),
.A2(n_1598),
.B1(n_1618),
.B2(n_1613),
.C(n_1616),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1619),
.A2(n_1610),
.B1(n_1697),
.B2(n_1730),
.C(n_1728),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1702),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1580),
.A2(n_1624),
.B1(n_1631),
.B2(n_1642),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1610),
.A2(n_1751),
.B1(n_1680),
.B2(n_1740),
.C(n_1735),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1627),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1731),
.B(n_1719),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1647),
.A2(n_1645),
.B1(n_1692),
.B2(n_1648),
.Y(n_1831)
);

BUFx4f_ASAP7_75t_SL g1832 ( 
.A(n_1651),
.Y(n_1832)
);

BUFx12f_ASAP7_75t_L g1833 ( 
.A(n_1708),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1651),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1564),
.A2(n_1576),
.B1(n_1647),
.B2(n_1608),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1574),
.A2(n_1631),
.B1(n_1642),
.B2(n_1698),
.Y(n_1836)
);

AO31x2_ASAP7_75t_L g1837 ( 
.A1(n_1747),
.A2(n_1701),
.A3(n_1741),
.B(n_1749),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1596),
.A2(n_1594),
.B(n_1734),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1640),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1609),
.A2(n_1754),
.B1(n_1665),
.B2(n_1698),
.Y(n_1840)
);

BUFx4f_ASAP7_75t_SL g1841 ( 
.A(n_1651),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1720),
.Y(n_1842)
);

BUFx4f_ASAP7_75t_SL g1843 ( 
.A(n_1651),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1562),
.A2(n_1685),
.B1(n_1737),
.B2(n_1707),
.Y(n_1844)
);

AND2x4_ASAP7_75t_SL g1845 ( 
.A(n_1719),
.B(n_1572),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1665),
.A2(n_1726),
.B1(n_1701),
.B2(n_1744),
.C(n_1704),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1664),
.A2(n_1585),
.B1(n_1743),
.B2(n_1719),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1585),
.B(n_1704),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1670),
.A2(n_1731),
.B(n_1744),
.C(n_1748),
.Y(n_1849)
);

AOI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1717),
.A2(n_1722),
.B(n_1725),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1726),
.A2(n_1721),
.B1(n_1718),
.B2(n_1733),
.C(n_1739),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1713),
.A2(n_1745),
.B1(n_1566),
.B2(n_1559),
.C(n_1599),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1699),
.Y(n_1853)
);

OAI222xp33_ASAP7_75t_L g1854 ( 
.A1(n_1717),
.A2(n_1703),
.B1(n_1599),
.B2(n_1601),
.C1(n_1706),
.C2(n_1643),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1710),
.B(n_1703),
.Y(n_1855)
);

O2A1O1Ixp5_ASAP7_75t_L g1856 ( 
.A1(n_1753),
.A2(n_1748),
.B(n_1750),
.C(n_1727),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1685),
.A2(n_1719),
.B1(n_1578),
.B2(n_1706),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1717),
.A2(n_1722),
.B1(n_1710),
.B2(n_1683),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1683),
.A2(n_1691),
.B1(n_1746),
.B2(n_1643),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1664),
.A2(n_1745),
.B1(n_1601),
.B2(n_1678),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1699),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1745),
.A2(n_1699),
.B(n_1644),
.C(n_1617),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1714),
.B(n_1569),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1714),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1714),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1558),
.B(n_1581),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1562),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1569),
.B(n_1588),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1870)
);

INVxp33_ASAP7_75t_L g1871 ( 
.A(n_1563),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1603),
.Y(n_1872)
);

OAI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.C(n_1135),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1594),
.A2(n_1156),
.B(n_1481),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1686),
.A2(n_1156),
.B1(n_560),
.B2(n_1117),
.C(n_1010),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1709),
.Y(n_1876)
);

OAI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.C(n_1135),
.Y(n_1877)
);

OAI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.C(n_1135),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1686),
.A2(n_1156),
.B1(n_560),
.B2(n_1117),
.C(n_1010),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1563),
.Y(n_1880)
);

OA21x2_ASAP7_75t_L g1881 ( 
.A1(n_1620),
.A2(n_1744),
.B(n_1734),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1571),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1724),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1639),
.A2(n_1135),
.B1(n_1676),
.B2(n_1655),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1888)
);

OAI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1639),
.A2(n_1135),
.B1(n_1676),
.B2(n_1655),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1586),
.B(n_1421),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1709),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1561),
.B(n_1156),
.C(n_1117),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1893)
);

OR2x6_ASAP7_75t_L g1894 ( 
.A(n_1698),
.B(n_1717),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1570),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1135),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1571),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1683),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1630),
.A2(n_1117),
.B(n_1156),
.C(n_1144),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1620),
.A2(n_1744),
.B(n_1734),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1571),
.Y(n_1901)
);

OAI33xp33_ASAP7_75t_L g1902 ( 
.A1(n_1686),
.A2(n_1639),
.A3(n_1655),
.B1(n_724),
.B2(n_720),
.B3(n_1568),
.Y(n_1902)
);

OA21x2_ASAP7_75t_L g1903 ( 
.A1(n_1620),
.A2(n_1744),
.B(n_1734),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1709),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1586),
.B(n_1421),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1135),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1561),
.A2(n_1156),
.B1(n_1117),
.B2(n_1144),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1675),
.B(n_712),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1586),
.B(n_1421),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1561),
.A2(n_1156),
.B(n_1117),
.Y(n_1910)
);

INVx11_ASAP7_75t_L g1911 ( 
.A(n_1711),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1570),
.Y(n_1912)
);

AOI221xp5_ASAP7_75t_L g1913 ( 
.A1(n_1686),
.A2(n_1156),
.B1(n_560),
.B2(n_1117),
.C(n_1010),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1561),
.A2(n_1156),
.B(n_1117),
.Y(n_1914)
);

AO31x2_ASAP7_75t_L g1915 ( 
.A1(n_1752),
.A2(n_1742),
.A3(n_1747),
.B(n_1730),
.Y(n_1915)
);

INVx4_ASAP7_75t_L g1916 ( 
.A(n_1659),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1686),
.A2(n_1156),
.B1(n_560),
.B2(n_1117),
.C(n_1010),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1863),
.B(n_1869),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1894),
.B(n_1775),
.Y(n_1919)
);

INVx4_ASAP7_75t_L g1920 ( 
.A(n_1894),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1779),
.B(n_1810),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1882),
.A2(n_1917),
.B1(n_1875),
.B2(n_1913),
.C(n_1879),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1908),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1890),
.B(n_1905),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1759),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1759),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1866),
.B(n_1761),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1769),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1775),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1783),
.B(n_1828),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1864),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1784),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1894),
.B(n_1775),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1799),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_SL g1935 ( 
.A(n_1821),
.B(n_1808),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1803),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1883),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1897),
.B(n_1901),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1761),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1839),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1805),
.B(n_1822),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1830),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1909),
.B(n_1842),
.Y(n_1943)
);

AO21x2_ASAP7_75t_L g1944 ( 
.A1(n_1785),
.A2(n_1757),
.B(n_1838),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1881),
.B(n_1900),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1880),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1830),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1862),
.Y(n_1948)
);

INVxp67_ASAP7_75t_SL g1949 ( 
.A(n_1781),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1793),
.B(n_1814),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1818),
.B(n_1848),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1818),
.B(n_1881),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1837),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1900),
.B(n_1903),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1856),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_SL g1956 ( 
.A(n_1791),
.B(n_1763),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1903),
.B(n_1840),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1856),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1791),
.B(n_1915),
.Y(n_1959)
);

NOR2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1892),
.B(n_1756),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1915),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1915),
.B(n_1758),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1868),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1855),
.B(n_1847),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_L g1965 ( 
.A(n_1914),
.B(n_1910),
.C(n_1870),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1915),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1868),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1846),
.B(n_1876),
.Y(n_1968)
);

AO31x2_ASAP7_75t_L g1969 ( 
.A1(n_1865),
.A2(n_1786),
.A3(n_1771),
.B(n_1849),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1871),
.B(n_1766),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1891),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_L g1972 ( 
.A(n_1867),
.B(n_1870),
.C(n_1893),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1904),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1778),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1811),
.Y(n_1975)
);

INVx5_ASAP7_75t_SL g1976 ( 
.A(n_1756),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1860),
.B(n_1801),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1895),
.B(n_1912),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1789),
.B(n_1825),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1844),
.B(n_1773),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1817),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1789),
.B(n_1804),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1844),
.B(n_1773),
.Y(n_1983)
);

NOR2xp67_ASAP7_75t_L g1984 ( 
.A(n_1850),
.B(n_1824),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1782),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1807),
.B(n_1857),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1782),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1794),
.B(n_1813),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1858),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1873),
.A2(n_1878),
.B1(n_1877),
.B2(n_1867),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1853),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1859),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1886),
.A2(n_1888),
.B1(n_1893),
.B2(n_1885),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1857),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1835),
.B(n_1851),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1813),
.B(n_1886),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1888),
.B(n_1907),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1760),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1831),
.B(n_1795),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1831),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1816),
.B(n_1806),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1777),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1835),
.B(n_1764),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1777),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1852),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1872),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1774),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1812),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1896),
.B(n_1906),
.Y(n_2009)
);

INVx4_ASAP7_75t_L g2010 ( 
.A(n_1756),
.Y(n_2010)
);

OA21x2_ASAP7_75t_L g2011 ( 
.A1(n_1961),
.A2(n_1874),
.B(n_1854),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1922),
.A2(n_1788),
.B1(n_1790),
.B2(n_1889),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1956),
.A2(n_1800),
.B(n_1887),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_L g2014 ( 
.A(n_1965),
.B(n_1899),
.C(n_1768),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1963),
.B(n_1816),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_2006),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1928),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_L g2018 ( 
.A(n_1990),
.B(n_1768),
.C(n_1796),
.D(n_1792),
.Y(n_2018)
);

BUFx2_ASAP7_75t_L g2019 ( 
.A(n_1929),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1972),
.A2(n_1889),
.B1(n_1887),
.B2(n_1902),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1918),
.B(n_1762),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1925),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1931),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1918),
.B(n_1772),
.Y(n_2024)
);

AOI33xp33_ASAP7_75t_L g2025 ( 
.A1(n_1979),
.A2(n_1826),
.A3(n_1809),
.B1(n_1827),
.B2(n_1823),
.B3(n_1902),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1993),
.A2(n_1809),
.B1(n_1819),
.B2(n_1836),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1979),
.A2(n_1797),
.B1(n_1916),
.B2(n_1802),
.Y(n_2027)
);

CKINVDCx16_ASAP7_75t_R g2028 ( 
.A(n_2010),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1923),
.B(n_1916),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1967),
.B(n_1802),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_2006),
.Y(n_2031)
);

OAI31xp33_ASAP7_75t_L g2032 ( 
.A1(n_1982),
.A2(n_1845),
.A3(n_1898),
.B(n_1770),
.Y(n_2032)
);

NAND3xp33_ASAP7_75t_L g2033 ( 
.A(n_2007),
.B(n_1787),
.C(n_1776),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_2006),
.Y(n_2034)
);

OR2x6_ASAP7_75t_L g2035 ( 
.A(n_1919),
.B(n_1756),
.Y(n_2035)
);

INVx5_ASAP7_75t_L g2036 ( 
.A(n_1947),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1982),
.A2(n_1755),
.B1(n_1798),
.B2(n_1884),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1927),
.B(n_1767),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1921),
.B(n_1767),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1927),
.B(n_1776),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1981),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1947),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1981),
.Y(n_2043)
);

AO21x1_ASAP7_75t_SL g2044 ( 
.A1(n_2002),
.A2(n_1843),
.B(n_1841),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1921),
.B(n_1834),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_2009),
.A2(n_1755),
.B1(n_1798),
.B2(n_1884),
.Y(n_2046)
);

OAI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1997),
.A2(n_1884),
.B1(n_1820),
.B2(n_1841),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1995),
.A2(n_1884),
.B1(n_1833),
.B2(n_1780),
.Y(n_2048)
);

OAI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1996),
.A2(n_1765),
.B1(n_1829),
.B2(n_1898),
.C(n_1861),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1934),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1971),
.B(n_1780),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1949),
.B(n_1832),
.Y(n_2052)
);

OAI332xp33_ASAP7_75t_L g2053 ( 
.A1(n_1988),
.A2(n_1815),
.A3(n_1832),
.B1(n_1843),
.B2(n_1911),
.B3(n_2007),
.C1(n_1999),
.C2(n_2001),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1936),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2001),
.A2(n_2010),
.B1(n_1999),
.B2(n_1980),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1952),
.B(n_1985),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1941),
.B(n_1974),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1930),
.B(n_1950),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1930),
.B(n_1943),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1952),
.B(n_1985),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1929),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1976),
.Y(n_2062)
);

AOI222xp33_ASAP7_75t_L g2063 ( 
.A1(n_1995),
.A2(n_1984),
.B1(n_2003),
.B2(n_1935),
.C1(n_1977),
.C2(n_1960),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1960),
.A2(n_1984),
.B1(n_1986),
.B2(n_1983),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1937),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_1929),
.Y(n_2066)
);

NAND3xp33_ASAP7_75t_L g2067 ( 
.A(n_1974),
.B(n_1998),
.C(n_2000),
.Y(n_2067)
);

CKINVDCx20_ASAP7_75t_R g2068 ( 
.A(n_1976),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1941),
.B(n_1939),
.Y(n_2069)
);

AOI221xp5_ASAP7_75t_L g2070 ( 
.A1(n_2000),
.A2(n_2003),
.B1(n_2004),
.B2(n_2002),
.C(n_1998),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2004),
.A2(n_1998),
.B1(n_1977),
.B2(n_2005),
.C(n_1957),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_2008),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1932),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1940),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1986),
.A2(n_1983),
.B1(n_1980),
.B2(n_1975),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1987),
.B(n_1957),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1939),
.B(n_1962),
.Y(n_2077)
);

AO21x2_ASAP7_75t_L g2078 ( 
.A1(n_1961),
.A2(n_1966),
.B(n_1953),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1989),
.A2(n_1968),
.B1(n_1994),
.B2(n_1951),
.Y(n_2079)
);

INVx5_ASAP7_75t_SL g2080 ( 
.A(n_1947),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1924),
.A2(n_1946),
.B1(n_1976),
.B2(n_1989),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_1947),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1987),
.B(n_1964),
.Y(n_2083)
);

AOI33xp33_ASAP7_75t_L g2084 ( 
.A1(n_1968),
.A2(n_1948),
.A3(n_1992),
.B1(n_1954),
.B2(n_2005),
.B3(n_1958),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_1991),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2057),
.B(n_1926),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2057),
.B(n_1962),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2056),
.B(n_1954),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2036),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2022),
.B(n_2069),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2069),
.B(n_2058),
.Y(n_2091)
);

INVx2_ASAP7_75t_SL g2092 ( 
.A(n_2036),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_2036),
.B(n_1919),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2056),
.B(n_1945),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2077),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_2023),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_1945),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2076),
.B(n_1955),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2059),
.B(n_1973),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_2036),
.B(n_1919),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2050),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2076),
.B(n_1955),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2036),
.B(n_1933),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2083),
.B(n_1958),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2054),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2054),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2065),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2083),
.B(n_1933),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_2077),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2024),
.B(n_1933),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2040),
.B(n_1969),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2019),
.B(n_1948),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2019),
.B(n_1920),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_2085),
.Y(n_2114)
);

NOR2x1_ASAP7_75t_L g2115 ( 
.A(n_2067),
.B(n_1920),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2074),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2040),
.B(n_1969),
.Y(n_2117)
);

HB1xp67_ASAP7_75t_L g2118 ( 
.A(n_2072),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2021),
.B(n_2039),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2035),
.B(n_1920),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2073),
.B(n_1938),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2021),
.B(n_2039),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2078),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2061),
.B(n_1969),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2017),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2061),
.B(n_1969),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2066),
.B(n_1969),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2035),
.B(n_1920),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_2078),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2066),
.B(n_1969),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2011),
.B(n_1944),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2038),
.B(n_1944),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2045),
.B(n_1964),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_2038),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2123),
.Y(n_2135)
);

INVxp67_ASAP7_75t_SL g2136 ( 
.A(n_2115),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2105),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2119),
.B(n_2071),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_2114),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2115),
.A2(n_2014),
.B(n_2063),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2088),
.B(n_2016),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2105),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2132),
.B(n_1944),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2120),
.A2(n_2013),
.B1(n_2033),
.B2(n_2018),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2112),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2119),
.B(n_2070),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2105),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2088),
.B(n_2034),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2087),
.B(n_2015),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2088),
.B(n_2045),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2119),
.B(n_2122),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2112),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2098),
.B(n_2031),
.Y(n_2153)
);

NAND2x2_ASAP7_75t_L g2154 ( 
.A(n_2089),
.B(n_2031),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2087),
.B(n_2030),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_2113),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2111),
.B(n_1959),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_2118),
.B(n_2051),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2098),
.B(n_2043),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2111),
.B(n_2117),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2098),
.B(n_2043),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2122),
.B(n_2084),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2102),
.B(n_2122),
.Y(n_2163)
);

INVxp67_ASAP7_75t_L g2164 ( 
.A(n_2125),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2123),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_2099),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2093),
.B(n_2042),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2117),
.B(n_1959),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2106),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2095),
.B(n_1992),
.Y(n_2170)
);

OAI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_2131),
.A2(n_2012),
.B(n_2020),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2102),
.B(n_2041),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2107),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2102),
.B(n_2042),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2123),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2094),
.B(n_2082),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2095),
.B(n_2011),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2107),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_2091),
.B(n_2029),
.Y(n_2179)
);

HB1xp67_ASAP7_75t_L g2180 ( 
.A(n_2104),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2094),
.B(n_2097),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2116),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2116),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2091),
.B(n_2013),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2094),
.B(n_2082),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2116),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2097),
.B(n_1942),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2101),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2188),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_2163),
.B(n_2093),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_SL g2191 ( 
.A1(n_2140),
.A2(n_2027),
.B(n_2026),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2171),
.B(n_2110),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2163),
.B(n_2110),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2151),
.B(n_2090),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2182),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2139),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2151),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2171),
.B(n_2110),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2182),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2160),
.B(n_2090),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2146),
.B(n_2104),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2160),
.B(n_2086),
.Y(n_2203)
);

INVx4_ASAP7_75t_L g2204 ( 
.A(n_2167),
.Y(n_2204)
);

OA21x2_ASAP7_75t_L g2205 ( 
.A1(n_2140),
.A2(n_2131),
.B(n_2096),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2134),
.B(n_2086),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2167),
.B(n_2108),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2186),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2146),
.B(n_2162),
.Y(n_2209)
);

AOI21xp33_ASAP7_75t_L g2210 ( 
.A1(n_2136),
.A2(n_2013),
.B(n_2064),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2186),
.Y(n_2211)
);

INVx1_ASAP7_75t_SL g2212 ( 
.A(n_2156),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2167),
.B(n_2108),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_2134),
.B(n_2109),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_2154),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2184),
.B(n_2109),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_2167),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2145),
.B(n_2108),
.Y(n_2218)
);

AND4x1_ASAP7_75t_L g2219 ( 
.A(n_2144),
.B(n_2037),
.C(n_2048),
.D(n_2046),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2188),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2164),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2164),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2162),
.B(n_2138),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2156),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2145),
.B(n_2097),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_R g2226 ( 
.A(n_2138),
.B(n_2062),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2184),
.B(n_2121),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2170),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2186),
.Y(n_2229)
);

INVx6_ASAP7_75t_L g2230 ( 
.A(n_2154),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2149),
.B(n_2121),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2179),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2166),
.B(n_2104),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2137),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2137),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2142),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2149),
.B(n_2133),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2158),
.B(n_2133),
.Y(n_2238)
);

NAND2x1_ASAP7_75t_L g2239 ( 
.A(n_2177),
.B(n_2089),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2150),
.B(n_2099),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2154),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2135),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2202),
.B(n_2143),
.Y(n_2243)
);

INVx1_ASAP7_75t_SL g2244 ( 
.A(n_2226),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2207),
.B(n_2152),
.Y(n_2245)
);

AOI322xp5_ASAP7_75t_L g2246 ( 
.A1(n_2223),
.A2(n_2079),
.A3(n_2131),
.B1(n_2152),
.B2(n_2075),
.C1(n_2124),
.C2(n_2126),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2196),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2189),
.Y(n_2248)
);

OAI31xp33_ASAP7_75t_L g2249 ( 
.A1(n_2191),
.A2(n_2047),
.A3(n_2049),
.B(n_2127),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2232),
.B(n_2155),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2239),
.Y(n_2251)
);

OAI21xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2219),
.A2(n_2209),
.B(n_2199),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2192),
.B(n_2150),
.Y(n_2253)
);

OAI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2210),
.A2(n_2143),
.B1(n_2177),
.B2(n_2032),
.C(n_2168),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2237),
.B(n_2157),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2238),
.B(n_2187),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2189),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2228),
.B(n_2187),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2212),
.B(n_2172),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2205),
.A2(n_2053),
.B(n_1935),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2207),
.B(n_2181),
.Y(n_2261)
);

INVx1_ASAP7_75t_SL g2262 ( 
.A(n_2230),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2221),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2230),
.A2(n_2055),
.B1(n_2100),
.B2(n_2093),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2224),
.B(n_2172),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2213),
.B(n_2181),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2222),
.B(n_2141),
.Y(n_2267)
);

OAI32xp33_ASAP7_75t_L g2268 ( 
.A1(n_2216),
.A2(n_2168),
.A3(n_2157),
.B1(n_2124),
.B2(n_2130),
.Y(n_2268)
);

OAI211xp5_ASAP7_75t_L g2269 ( 
.A1(n_2205),
.A2(n_2239),
.B(n_2197),
.C(n_2215),
.Y(n_2269)
);

AOI21xp33_ASAP7_75t_SL g2270 ( 
.A1(n_2205),
.A2(n_2081),
.B(n_2092),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2193),
.B(n_2141),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2193),
.B(n_2148),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2217),
.Y(n_2273)
);

AOI21xp33_ASAP7_75t_SL g2274 ( 
.A1(n_2215),
.A2(n_2092),
.B(n_2089),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2220),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2220),
.Y(n_2276)
);

OAI221xp5_ASAP7_75t_L g2277 ( 
.A1(n_2241),
.A2(n_2170),
.B1(n_2092),
.B2(n_2155),
.C(n_2126),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2234),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2195),
.Y(n_2279)
);

AO22x1_ASAP7_75t_L g2280 ( 
.A1(n_2241),
.A2(n_1978),
.B1(n_2093),
.B2(n_2100),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2194),
.B(n_2180),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2234),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2213),
.B(n_2204),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2230),
.A2(n_2093),
.B1(n_2100),
.B2(n_2103),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2235),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2283),
.B(n_2204),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2248),
.Y(n_2287)
);

AOI221xp5_ASAP7_75t_L g2288 ( 
.A1(n_2252),
.A2(n_2204),
.B1(n_2217),
.B2(n_2126),
.C(n_2124),
.Y(n_2288)
);

AOI211xp5_ASAP7_75t_L g2289 ( 
.A1(n_2249),
.A2(n_2214),
.B(n_2216),
.C(n_2206),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2248),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2260),
.B(n_2217),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2281),
.B(n_2194),
.Y(n_2292)
);

O2A1O1Ixp33_ASAP7_75t_SL g2293 ( 
.A1(n_2244),
.A2(n_2214),
.B(n_1970),
.C(n_2201),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_2247),
.B(n_2262),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2273),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2250),
.B(n_2218),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2275),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_SL g2298 ( 
.A1(n_2269),
.A2(n_2198),
.B(n_2195),
.C(n_2200),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2273),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2275),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2285),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2283),
.B(n_2190),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2285),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2264),
.A2(n_2206),
.B(n_2233),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_2245),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2257),
.Y(n_2306)
);

AOI211xp5_ASAP7_75t_L g2307 ( 
.A1(n_2270),
.A2(n_2130),
.B(n_2127),
.C(n_2190),
.Y(n_2307)
);

AOI21xp33_ASAP7_75t_L g2308 ( 
.A1(n_2263),
.A2(n_2227),
.B(n_2236),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2245),
.B(n_2190),
.Y(n_2309)
);

NOR2xp67_ASAP7_75t_L g2310 ( 
.A(n_2274),
.B(n_2201),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2284),
.A2(n_2230),
.B1(n_2100),
.B2(n_2103),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2246),
.B(n_2218),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2259),
.A2(n_2100),
.B1(n_2103),
.B2(n_2128),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2276),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2278),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_2281),
.B(n_2203),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2305),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2309),
.B(n_2261),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2301),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2294),
.B(n_2261),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2301),
.Y(n_2321)
);

NAND2xp33_ASAP7_75t_SL g2322 ( 
.A(n_2312),
.B(n_2251),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2296),
.B(n_2266),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2287),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2290),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_2292),
.Y(n_2326)
);

INVx1_ASAP7_75t_SL g2327 ( 
.A(n_2292),
.Y(n_2327)
);

XOR2xp5_ASAP7_75t_L g2328 ( 
.A(n_2299),
.B(n_2267),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2297),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2300),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_SL g2331 ( 
.A(n_2310),
.B(n_2254),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2295),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2289),
.B(n_2266),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2303),
.Y(n_2334)
);

NAND2xp33_ASAP7_75t_SL g2335 ( 
.A(n_2291),
.B(n_2251),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2306),
.Y(n_2336)
);

INVx3_ASAP7_75t_SL g2337 ( 
.A(n_2295),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2293),
.B(n_2265),
.Y(n_2338)
);

XOR2x2_ASAP7_75t_L g2339 ( 
.A(n_2288),
.B(n_2280),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2286),
.Y(n_2340)
);

NAND2xp33_ASAP7_75t_L g2341 ( 
.A(n_2326),
.B(n_2316),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2327),
.B(n_2314),
.Y(n_2342)
);

NOR3x1_ASAP7_75t_L g2343 ( 
.A(n_2333),
.B(n_2298),
.C(n_2291),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2331),
.B(n_2298),
.C(n_2293),
.Y(n_2344)
);

AND3x4_ASAP7_75t_L g2345 ( 
.A(n_2328),
.B(n_2103),
.C(n_2120),
.Y(n_2345)
);

NAND3x1_ASAP7_75t_L g2346 ( 
.A(n_2317),
.B(n_2315),
.C(n_2286),
.Y(n_2346)
);

INVxp67_ASAP7_75t_L g2347 ( 
.A(n_2335),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2318),
.B(n_2309),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2320),
.B(n_2316),
.Y(n_2349)
);

AOI21xp33_ASAP7_75t_L g2350 ( 
.A1(n_2338),
.A2(n_2307),
.B(n_2308),
.Y(n_2350)
);

XNOR2xp5_ASAP7_75t_L g2351 ( 
.A(n_2328),
.B(n_2311),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2332),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2319),
.Y(n_2353)
);

NAND4xp75_ASAP7_75t_L g2354 ( 
.A(n_2338),
.B(n_2302),
.C(n_2304),
.D(n_2313),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2321),
.Y(n_2355)
);

AOI222xp33_ASAP7_75t_L g2356 ( 
.A1(n_2344),
.A2(n_2322),
.B1(n_2335),
.B2(n_2339),
.C1(n_2337),
.C2(n_2336),
.Y(n_2356)
);

AOI321xp33_ASAP7_75t_L g2357 ( 
.A1(n_2350),
.A2(n_2323),
.A3(n_2318),
.B1(n_2322),
.B2(n_2339),
.C(n_2334),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2354),
.A2(n_2340),
.B1(n_2337),
.B2(n_2277),
.Y(n_2358)
);

OAI32xp33_ASAP7_75t_L g2359 ( 
.A1(n_2350),
.A2(n_2330),
.A3(n_2329),
.B1(n_2325),
.B2(n_2324),
.Y(n_2359)
);

AOI211xp5_ASAP7_75t_L g2360 ( 
.A1(n_2341),
.A2(n_2347),
.B(n_2351),
.C(n_2349),
.Y(n_2360)
);

AOI221x1_ASAP7_75t_L g2361 ( 
.A1(n_2352),
.A2(n_2282),
.B1(n_2302),
.B2(n_2279),
.C(n_2258),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2342),
.B(n_2253),
.Y(n_2362)
);

AOI222xp33_ASAP7_75t_L g2363 ( 
.A1(n_2342),
.A2(n_2268),
.B1(n_2280),
.B2(n_2279),
.C1(n_2256),
.C2(n_2272),
.Y(n_2363)
);

OAI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2343),
.A2(n_2348),
.B1(n_2271),
.B2(n_2355),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2346),
.A2(n_2255),
.B1(n_2203),
.B2(n_2243),
.Y(n_2365)
);

AOI222xp33_ASAP7_75t_L g2366 ( 
.A1(n_2353),
.A2(n_2268),
.B1(n_2127),
.B2(n_2130),
.C1(n_2225),
.C2(n_2229),
.Y(n_2366)
);

AOI21xp33_ASAP7_75t_SL g2367 ( 
.A1(n_2345),
.A2(n_2243),
.B(n_2255),
.Y(n_2367)
);

NAND4xp75_ASAP7_75t_L g2368 ( 
.A(n_2343),
.B(n_2225),
.C(n_2229),
.D(n_2236),
.Y(n_2368)
);

OAI221xp5_ASAP7_75t_L g2369 ( 
.A1(n_2357),
.A2(n_2356),
.B1(n_2360),
.B2(n_2358),
.C(n_2363),
.Y(n_2369)
);

OAI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2368),
.A2(n_2227),
.B1(n_2231),
.B2(n_1976),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_R g2371 ( 
.A(n_2362),
.B(n_2062),
.Y(n_2371)
);

AOI21xp33_ASAP7_75t_SL g2372 ( 
.A1(n_2364),
.A2(n_2231),
.B(n_2235),
.Y(n_2372)
);

INVxp67_ASAP7_75t_L g2373 ( 
.A(n_2361),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2365),
.Y(n_2374)
);

OAI21xp33_ASAP7_75t_SL g2375 ( 
.A1(n_2366),
.A2(n_2367),
.B(n_2359),
.Y(n_2375)
);

AOI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_2242),
.B1(n_2198),
.B2(n_2211),
.C(n_2208),
.Y(n_2376)
);

AOI222xp33_ASAP7_75t_L g2377 ( 
.A1(n_2375),
.A2(n_2242),
.B1(n_2200),
.B2(n_2211),
.C1(n_2208),
.C2(n_2175),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2374),
.Y(n_2378)
);

NOR3xp33_ASAP7_75t_L g2379 ( 
.A(n_2373),
.B(n_2025),
.C(n_2240),
.Y(n_2379)
);

OAI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2372),
.A2(n_2165),
.B(n_2135),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2370),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2371),
.B(n_2148),
.Y(n_2382)
);

NOR2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2374),
.B(n_2052),
.Y(n_2383)
);

OA22x2_ASAP7_75t_L g2384 ( 
.A1(n_2378),
.A2(n_2135),
.B1(n_2165),
.B2(n_2175),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2382),
.Y(n_2385)
);

AND4x1_ASAP7_75t_L g2386 ( 
.A(n_2379),
.B(n_1976),
.C(n_2153),
.D(n_2159),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2381),
.A2(n_2103),
.B1(n_2080),
.B2(n_2120),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2376),
.A2(n_2377),
.B(n_2380),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2383),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_L g2390 ( 
.A(n_2378),
.B(n_2165),
.C(n_2175),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_2385),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2389),
.Y(n_2392)
);

CKINVDCx16_ASAP7_75t_R g2393 ( 
.A(n_2386),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2387),
.B(n_2388),
.Y(n_2394)
);

OR5x1_ASAP7_75t_L g2395 ( 
.A(n_2393),
.B(n_2384),
.C(n_2390),
.D(n_2129),
.E(n_2185),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2395),
.A2(n_2394),
.B1(n_2391),
.B2(n_2392),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2396),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2396),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2397),
.B(n_2394),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2398),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2400),
.A2(n_2153),
.B1(n_2159),
.B2(n_2161),
.Y(n_2401)
);

OAI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2399),
.A2(n_2169),
.B1(n_2183),
.B2(n_2142),
.C(n_2178),
.Y(n_2402)
);

AOI322xp5_ASAP7_75t_L g2403 ( 
.A1(n_2401),
.A2(n_2174),
.A3(n_2161),
.B1(n_2176),
.B2(n_2185),
.C1(n_2113),
.C2(n_2173),
.Y(n_2403)
);

OAI221xp5_ASAP7_75t_R g2404 ( 
.A1(n_2403),
.A2(n_2402),
.B1(n_2068),
.B2(n_2028),
.C(n_2044),
.Y(n_2404)
);

AOI211xp5_ASAP7_75t_L g2405 ( 
.A1(n_2404),
.A2(n_2183),
.B(n_2178),
.C(n_2147),
.Y(n_2405)
);


endmodule