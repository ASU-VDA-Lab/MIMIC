module fake_jpeg_13162_n_458 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_458);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_458;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_49),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_50),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_55),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_24),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_75),
.Y(n_122)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_86),
.Y(n_135)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_15),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_15),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_25),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_97),
.B(n_1),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_23),
.B1(n_36),
.B2(n_21),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_109),
.B1(n_123),
.B2(n_130),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_23),
.B1(n_36),
.B2(n_21),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_36),
.B1(n_23),
.B2(n_46),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_138),
.B1(n_85),
.B2(n_60),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_18),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_133),
.B1(n_137),
.B2(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_18),
.B1(n_43),
.B2(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_32),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_32),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_28),
.B1(n_43),
.B2(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_48),
.A2(n_39),
.B1(n_31),
.B2(n_26),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_38),
.B1(n_39),
.B2(n_31),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_68),
.A2(n_46),
.B1(n_38),
.B2(n_26),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_74),
.A2(n_46),
.B1(n_25),
.B2(n_20),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_69),
.Y(n_155)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_160),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_159),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_86),
.B1(n_49),
.B2(n_51),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_105),
.B1(n_102),
.B2(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_69),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_146),
.B(n_96),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_82),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_187),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_91),
.B1(n_59),
.B2(n_56),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_164),
.A2(n_188),
.B1(n_130),
.B2(n_144),
.Y(n_223)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_100),
.A2(n_60),
.B(n_58),
.C(n_50),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_194),
.Y(n_204)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_171),
.Y(n_208)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_77),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_100),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_182),
.Y(n_233)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_79),
.B1(n_77),
.B2(n_58),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_186),
.B1(n_193),
.B2(n_131),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_118),
.A2(n_79),
.B1(n_50),
.B2(n_3),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_97),
.B(n_1),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_135),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_98),
.B(n_2),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_2),
.Y(n_237)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_107),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_196),
.A2(n_223),
.B(n_224),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_146),
.B(n_124),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_205),
.A2(n_121),
.B(n_185),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_207),
.A2(n_156),
.B(n_193),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_230),
.B1(n_156),
.B2(n_184),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_107),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_183),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_157),
.A2(n_127),
.B1(n_119),
.B2(n_144),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_168),
.A2(n_127),
.B1(n_119),
.B2(n_105),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_161),
.A2(n_99),
.B1(n_126),
.B2(n_102),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_186),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_99),
.B1(n_108),
.B2(n_131),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_152),
.A2(n_108),
.B1(n_121),
.B2(n_143),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_231),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_238),
.B(n_243),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_240),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_183),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_222),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_245),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_163),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_249),
.B(n_255),
.Y(n_306)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_204),
.A2(n_163),
.B(n_188),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_251),
.A2(n_197),
.B(n_220),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_160),
.C(n_147),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_259),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_207),
.B1(n_234),
.B2(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_168),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_264),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_201),
.B(n_165),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_205),
.A2(n_164),
.B(n_179),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_260),
.B(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_221),
.B(n_213),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_154),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_223),
.A2(n_164),
.B(n_158),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_222),
.B1(n_214),
.B2(n_197),
.Y(n_289)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_269),
.B1(n_216),
.B2(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_177),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_153),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_266),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_208),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_151),
.C(n_195),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_272),
.Y(n_298)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_270),
.A2(n_274),
.B(n_261),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_199),
.B(n_167),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_170),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_143),
.B(n_150),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_196),
.A2(n_192),
.B(n_175),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_200),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_227),
.Y(n_304)
);

BUFx4f_ASAP7_75t_SL g324 ( 
.A(n_276),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_277),
.A2(n_244),
.B1(n_261),
.B2(n_272),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_230),
.B1(n_212),
.B2(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_278),
.A2(n_283),
.B1(n_286),
.B2(n_288),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_249),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_281),
.B(n_290),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_206),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_257),
.B(n_247),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_224),
.B1(n_216),
.B2(n_215),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_231),
.B1(n_149),
.B2(n_206),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_289),
.A2(n_245),
.B1(n_250),
.B2(n_269),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_214),
.C(n_227),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_256),
.C(n_248),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_305),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_261),
.B(n_262),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_242),
.A2(n_220),
.B1(n_226),
.B2(n_198),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_198),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_310),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_267),
.B(n_273),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_240),
.B(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_270),
.B(n_274),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_335),
.B1(n_288),
.B2(n_331),
.Y(n_341)
);

XOR2x1_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_251),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_313),
.B(n_328),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_333),
.B(n_339),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_318),
.C(n_319),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_268),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_256),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_306),
.B(n_255),
.Y(n_329)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_280),
.B(n_284),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_292),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_282),
.B(n_294),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_332),
.A2(n_308),
.B1(n_282),
.B2(n_296),
.Y(n_346)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_336),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_305),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_250),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_291),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_294),
.A2(n_226),
.B(n_258),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_269),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_330),
.C(n_319),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_360),
.B1(n_299),
.B2(n_324),
.Y(n_376)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_328),
.A2(n_339),
.B(n_327),
.C(n_313),
.D(n_326),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_342),
.A2(n_345),
.B(n_301),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_343),
.B(n_318),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_286),
.B1(n_293),
.B2(n_281),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_344),
.A2(n_347),
.B1(n_353),
.B2(n_357),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_325),
.B1(n_322),
.B2(n_334),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_317),
.A2(n_286),
.B1(n_293),
.B2(n_278),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_356),
.C(n_314),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_277),
.B1(n_283),
.B2(n_279),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_292),
.C(n_307),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_338),
.A2(n_340),
.B1(n_332),
.B2(n_315),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_315),
.A2(n_323),
.B1(n_306),
.B2(n_298),
.Y(n_358)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_338),
.A2(n_298),
.B1(n_308),
.B2(n_303),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_362),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_337),
.A2(n_300),
.B1(n_301),
.B2(n_299),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_263),
.B1(n_241),
.B2(n_228),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_372),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_374),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_326),
.C(n_333),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_383),
.C(n_387),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_347),
.B1(n_341),
.B2(n_357),
.Y(n_390)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_365),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_343),
.B(n_363),
.Y(n_372)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_324),
.B(n_285),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_384),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_SL g378 ( 
.A1(n_361),
.A2(n_324),
.B(n_321),
.C(n_263),
.Y(n_378)
);

BUFx12f_ASAP7_75t_SL g401 ( 
.A(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_228),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_379),
.B(n_388),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_362),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_380),
.B(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_364),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_211),
.B(n_241),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_211),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_6),
.C(n_7),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_178),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_351),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_139),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_381),
.B1(n_378),
.B2(n_372),
.Y(n_413)
);

OAI321xp33_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_351),
.A3(n_354),
.B1(n_348),
.B2(n_353),
.C(n_342),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_396),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_352),
.C(n_344),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_370),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_398),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_385),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_369),
.B(n_375),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_SL g405 ( 
.A1(n_368),
.A2(n_366),
.A3(n_355),
.B1(n_365),
.B2(n_10),
.C1(n_7),
.C2(n_12),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_405),
.B(n_9),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_407),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_383),
.C(n_386),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_401),
.A2(n_377),
.B(n_378),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_411),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_375),
.C(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_395),
.B1(n_391),
.B2(n_402),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_378),
.C(n_8),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_417),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_7),
.B(n_8),
.Y(n_415)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_8),
.B(n_9),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_419),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_399),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_410),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_425),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_406),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_404),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_427),
.B(n_428),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_404),
.C(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_431),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_423),
.A2(n_416),
.B(n_409),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_435),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_392),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_416),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_439),
.B(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_438),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_420),
.A2(n_417),
.B(n_415),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_403),
.C(n_11),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_432),
.B(n_433),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_441),
.B(n_403),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_434),
.B(n_426),
.Y(n_444)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_425),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_447),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_430),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_429),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_10),
.B(n_11),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_451),
.A2(n_445),
.B(n_442),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g455 ( 
.A(n_453),
.B(n_454),
.C(n_449),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_452),
.C(n_10),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_10),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_12),
.Y(n_458)
);


endmodule