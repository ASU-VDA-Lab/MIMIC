module fake_jpeg_30865_n_44 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_9),
.B(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_26),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_31),
.B(n_32),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_13),
.B1(n_24),
.B2(n_25),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.C(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

AOI221xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.C(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_15),
.B1(n_23),
.B2(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_21),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_32),
.Y(n_43)
);

OAI321xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_21),
.A3(n_24),
.B1(n_28),
.B2(n_41),
.C(n_37),
.Y(n_44)
);


endmodule