module fake_jpeg_21155_n_355 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_46),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_8),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_14),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_51),
.Y(n_84)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_16),
.B1(n_24),
.B2(n_19),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_58),
.A2(n_63),
.B1(n_69),
.B2(n_85),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_16),
.B1(n_19),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_78),
.B1(n_82),
.B2(n_86),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_43),
.B1(n_54),
.B2(n_42),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_84),
.B1(n_56),
.B2(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_27),
.C(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_36),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_55),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_20),
.B1(n_30),
.B2(n_29),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_20),
.B1(n_30),
.B2(n_29),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_41),
.A2(n_26),
.B1(n_22),
.B2(n_35),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_81),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_13),
.B(n_12),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_98),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_105),
.B(n_44),
.Y(n_144)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_27),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_109),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_112),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_104),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_51),
.B(n_38),
.C(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_38),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_90),
.C(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_35),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_44),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_41),
.B1(n_44),
.B2(n_3),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_84),
.B1(n_64),
.B2(n_56),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_84),
.B1(n_67),
.B2(n_66),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_58),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_128),
.C(n_117),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_138),
.B1(n_140),
.B2(n_159),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_145),
.B1(n_91),
.B2(n_122),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_60),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_93),
.B(n_118),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_67),
.B1(n_76),
.B2(n_83),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_76),
.B1(n_57),
.B2(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_160),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_105),
.B(n_93),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_107),
.B1(n_125),
.B2(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_97),
.A2(n_12),
.B(n_11),
.C(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_1),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_96),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_57),
.B1(n_2),
.B2(n_4),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_165),
.Y(n_202)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_180),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_185),
.B(n_192),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_114),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_168),
.B(n_178),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_105),
.B1(n_127),
.B2(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_133),
.B1(n_141),
.B2(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_184),
.B1(n_159),
.B2(n_138),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_94),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_117),
.B1(n_122),
.B2(n_118),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_190),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_196),
.B1(n_135),
.B2(n_148),
.Y(n_211)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_183),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_134),
.B1(n_146),
.B2(n_131),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_94),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_121),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_143),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_10),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_136),
.C(n_141),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_208),
.C(n_167),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_226),
.B1(n_187),
.B2(n_175),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_164),
.C(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_217),
.B1(n_221),
.B2(n_224),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_156),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_153),
.B1(n_155),
.B2(n_160),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_121),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_110),
.B1(n_102),
.B2(n_100),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_197),
.B1(n_189),
.B2(n_193),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_129),
.B1(n_148),
.B2(n_158),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_96),
.A3(n_119),
.B1(n_92),
.B2(n_116),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_106),
.B1(n_10),
.B2(n_9),
.Y(n_224)
);

AO21x2_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_106),
.B(n_2),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_4),
.B(n_5),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_170),
.B(n_171),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_224),
.B1(n_201),
.B2(n_227),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_250),
.B1(n_252),
.B2(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_192),
.B(n_167),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_240),
.C(n_206),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_190),
.C(n_172),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_177),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_210),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_196),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_174),
.B1(n_185),
.B2(n_180),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_215),
.B1(n_225),
.B2(n_220),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_202),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_201),
.B(n_193),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_213),
.A2(n_5),
.B(n_6),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_263),
.C(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_254),
.C(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_208),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_225),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_240),
.B(n_218),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_211),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_209),
.C(n_217),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_199),
.C(n_215),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_256),
.B1(n_261),
.B2(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_225),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_284),
.B1(n_281),
.B2(n_278),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_232),
.B1(n_280),
.B2(n_225),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_232),
.B(n_256),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_301),
.B(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_246),
.B1(n_234),
.B2(n_252),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_297),
.B1(n_243),
.B2(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_296),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_237),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_242),
.C(n_230),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_274),
.C(n_263),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_261),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_315),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_265),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_308),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_6),
.Y(n_310)
);

BUFx12f_ASAP7_75t_SL g312 ( 
.A(n_294),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_6),
.B(n_7),
.C(n_285),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_287),
.B(n_291),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_293),
.B1(n_287),
.B2(n_295),
.Y(n_323)
);

BUFx12_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_296),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_309),
.B(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_288),
.B1(n_297),
.B2(n_283),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_326),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_292),
.C(n_299),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_327),
.C(n_320),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_310),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_293),
.C(n_300),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_334),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_319),
.A2(n_306),
.B1(n_289),
.B2(n_311),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_335),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_314),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_324),
.B(n_316),
.CI(n_313),
.CON(n_335),
.SN(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_316),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_335),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_329),
.C(n_331),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_319),
.B1(n_325),
.B2(n_322),
.Y(n_338)
);

NOR2x1_ASAP7_75t_SL g347 ( 
.A(n_338),
.B(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_337),
.B(n_327),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_340),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_344),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_348),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_347),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_349),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_346),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_350),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_349),
.Y(n_355)
);


endmodule