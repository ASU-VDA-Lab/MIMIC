module fake_netlist_6_1321_n_1568 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1568);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1568;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1558;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_49),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_169),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_360),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_1),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_217),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_17),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_216),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_78),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_95),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_57),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_196),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_78),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_96),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_356),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_14),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_55),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_40),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_322),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_274),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_179),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_210),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_272),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_97),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_63),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_16),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_231),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_133),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_237),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_240),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_138),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_98),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_193),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_290),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_119),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_206),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_282),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_223),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_211),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_79),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_265),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_139),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_239),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_336),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_57),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_153),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_82),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_369),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_262),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_203),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_354),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_174),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_16),
.Y(n_437)
);

INVx4_ASAP7_75t_R g438 ( 
.A(n_224),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_242),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_43),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_253),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_110),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_170),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_226),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_188),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_233),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_292),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_37),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_107),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_50),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_346),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_0),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_42),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_92),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_349),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_94),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_328),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_42),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_370),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_117),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_15),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_165),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_53),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_344),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_355),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_55),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_298),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_93),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_60),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_6),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_77),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_77),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_3),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_250),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_348),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_181),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_202),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_189),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_0),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_304),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_70),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_215),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_152),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_137),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_273),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_267),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_135),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_183),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_28),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_347),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_39),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_209),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_190),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_159),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_9),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_132),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_39),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_305),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_161),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_156),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_103),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_11),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_74),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_207),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_65),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_140),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_155),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_65),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_40),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_341),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_342),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_45),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_374),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_63),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_194),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_350),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_49),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_310),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_122),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_256),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_358),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_134),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_316),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_340),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_331),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_17),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_335),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_81),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_259),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_73),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_333),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_44),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_263),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_102),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_29),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_136),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_291),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_175),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_315),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_100),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_364),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_225),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_308),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_325),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_288),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_162),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_43),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_186),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_28),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_69),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_52),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_178),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_26),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_4),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_327),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_163),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_345),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_296),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_141),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_343),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_116),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_359),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_22),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_31),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_246),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_279),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_48),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_124),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_176),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_177),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_3),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_295),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_248),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_243),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_129),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_353),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_27),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_173),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_47),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_150),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_32),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_214),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_234),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_147),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_59),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_313),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_130),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_287),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_5),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_213),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_146),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_329),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_112),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_127),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_452),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_382),
.B(n_1),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_382),
.B(n_2),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_417),
.B(n_2),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_407),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_417),
.B(n_4),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_404),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_391),
.B(n_5),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_404),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_452),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_507),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_404),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_404),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_409),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_391),
.B(n_6),
.Y(n_611)
);

BUFx8_ASAP7_75t_L g612 ( 
.A(n_439),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

NOR2x1_ASAP7_75t_L g614 ( 
.A(n_399),
.B(n_7),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_407),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_409),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_465),
.B(n_7),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_409),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_587),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_587),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_409),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_436),
.B(n_8),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_380),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_436),
.B(n_8),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_443),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_397),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_407),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_532),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_443),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_443),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_447),
.B(n_9),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_483),
.Y(n_633)
);

BUFx8_ASAP7_75t_SL g634 ( 
.A(n_440),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_532),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_443),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_447),
.B(n_10),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_469),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_469),
.Y(n_639)
);

BUFx12f_ASAP7_75t_L g640 ( 
.A(n_532),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_469),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_385),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_491),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_559),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_388),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_559),
.B(n_10),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_376),
.B(n_11),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_442),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_442),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_442),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_465),
.B(n_12),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_399),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_458),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_475),
.Y(n_654)
);

BUFx12f_ASAP7_75t_L g655 ( 
.A(n_478),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_493),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

BUFx12f_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_478),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_556),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_458),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_466),
.B(n_12),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_466),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_543),
.B(n_13),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_13),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_544),
.B(n_547),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_544),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_389),
.B(n_14),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_547),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_375),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_377),
.Y(n_672)
);

BUFx12f_ASAP7_75t_L g673 ( 
.A(n_378),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_398),
.B(n_15),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_560),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_575),
.B(n_18),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_18),
.Y(n_677)
);

BUFx8_ASAP7_75t_SL g678 ( 
.A(n_472),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_567),
.B(n_19),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_514),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_528),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_379),
.B(n_19),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_468),
.B(n_20),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

CKINVDCx11_ASAP7_75t_R g687 ( 
.A(n_377),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_383),
.B(n_20),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_565),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_381),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_384),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_387),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_386),
.B(n_21),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_573),
.B(n_21),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_390),
.B(n_22),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_393),
.Y(n_697)
);

BUFx12f_ASAP7_75t_L g698 ( 
.A(n_392),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_488),
.B(n_23),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_403),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_395),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_414),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_579),
.B(n_23),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_418),
.B(n_24),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_438),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_396),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_394),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_420),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_406),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_495),
.B(n_24),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_400),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_424),
.B(n_25),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_425),
.B(n_25),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_426),
.B(n_430),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_435),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_422),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_572),
.B(n_26),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_448),
.B(n_27),
.Y(n_718)
);

BUFx12f_ASAP7_75t_L g719 ( 
.A(n_428),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_462),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_477),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_479),
.B(n_29),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_480),
.Y(n_723)
);

BUFx8_ASAP7_75t_SL g724 ( 
.A(n_530),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_437),
.B(n_450),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_486),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_487),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_489),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_705),
.B(n_401),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_603),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_603),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_674),
.A2(n_460),
.B1(n_463),
.B2(n_454),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_604),
.B(n_611),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_648),
.B(n_530),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_705),
.B(n_402),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_605),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_705),
.B(n_405),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_725),
.B(n_667),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_673),
.B(n_498),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_671),
.B(n_408),
.Y(n_742)
);

OA22x2_ASAP7_75t_L g743 ( 
.A1(n_654),
.A2(n_473),
.B1(n_474),
.B2(n_471),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_SL g744 ( 
.A1(n_672),
.A2(n_540),
.B1(n_548),
.B2(n_539),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_623),
.B(n_501),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_724),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_605),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_642),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_648),
.Y(n_749)
);

NAND3x1_ASAP7_75t_L g750 ( 
.A(n_614),
.B(n_512),
.C(n_509),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_699),
.B(n_539),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_691),
.B(n_410),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_699),
.A2(n_548),
.B1(n_550),
.B2(n_540),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_648),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_605),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_658),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_710),
.A2(n_561),
.B1(n_571),
.B2(n_550),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_672),
.A2(n_571),
.B1(n_561),
.B2(n_499),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_674),
.A2(n_504),
.B1(n_505),
.B2(n_481),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_676),
.A2(n_511),
.B1(n_516),
.B2(n_510),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_724),
.Y(n_761)
);

AO22x2_ASAP7_75t_L g762 ( 
.A1(n_679),
.A2(n_517),
.B1(n_518),
.B2(n_515),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_679),
.A2(n_521),
.B1(n_525),
.B2(n_520),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_676),
.A2(n_537),
.B1(n_549),
.B2(n_534),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_677),
.A2(n_553),
.B1(n_566),
.B2(n_551),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_608),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_677),
.A2(n_581),
.B1(n_583),
.B2(n_569),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_608),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_608),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_609),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_654),
.A2(n_591),
.B1(n_427),
.B2(n_431),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_647),
.A2(n_531),
.B1(n_541),
.B2(n_527),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_645),
.B(n_546),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_609),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_609),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_706),
.B(n_411),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_693),
.B(n_557),
.Y(n_777)
);

AO22x2_ASAP7_75t_L g778 ( 
.A1(n_617),
.A2(n_651),
.B1(n_664),
.B2(n_662),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_597),
.B(n_412),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_SL g780 ( 
.A1(n_647),
.A2(n_570),
.B1(n_584),
.B2(n_564),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_30),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_669),
.A2(n_444),
.B1(n_446),
.B2(n_416),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_669),
.A2(n_490),
.B1(n_494),
.B2(n_467),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_649),
.B(n_413),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_710),
.A2(n_526),
.B1(n_576),
.B2(n_496),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_598),
.A2(n_589),
.B1(n_592),
.B2(n_585),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_722),
.A2(n_593),
.B1(n_419),
.B2(n_421),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_631),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_707),
.B(n_415),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_722),
.A2(n_429),
.B1(n_432),
.B2(n_423),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_698),
.B(n_30),
.Y(n_792)
);

AO22x2_ASAP7_75t_L g793 ( 
.A1(n_689),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_649),
.B(n_650),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_598),
.A2(n_434),
.B1(n_441),
.B2(n_433),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_631),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_599),
.A2(n_449),
.B1(n_451),
.B2(n_445),
.Y(n_798)
);

OA22x2_ASAP7_75t_L g799 ( 
.A1(n_607),
.A2(n_456),
.B1(n_457),
.B2(n_453),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_689),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_717),
.A2(n_461),
.B1(n_464),
.B2(n_459),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_636),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_649),
.B(n_470),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_636),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_636),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_638),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_599),
.A2(n_482),
.B1(n_484),
.B2(n_476),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_650),
.B(n_485),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_638),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_701),
.B(n_34),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_717),
.A2(n_500),
.B1(n_502),
.B2(n_492),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_709),
.A2(n_506),
.B1(n_508),
.B2(n_503),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_650),
.Y(n_813)
);

OA22x2_ASAP7_75t_L g814 ( 
.A1(n_619),
.A2(n_522),
.B1(n_523),
.B2(n_513),
.Y(n_814)
);

OA22x2_ASAP7_75t_L g815 ( 
.A1(n_620),
.A2(n_529),
.B1(n_533),
.B2(n_524),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_638),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_711),
.B(n_535),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_718),
.A2(n_538),
.B1(n_542),
.B2(n_536),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_641),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_SL g820 ( 
.A1(n_600),
.A2(n_554),
.B1(n_558),
.B2(n_545),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_613),
.B(n_562),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_779),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_731),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_733),
.B(n_714),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_735),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_740),
.A2(n_602),
.B(n_600),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_735),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_733),
.B(n_714),
.Y(n_829)
);

XNOR2xp5_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_634),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_809),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_764),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

XOR2xp5_ASAP7_75t_L g834 ( 
.A(n_744),
.B(n_563),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_747),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_748),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_751),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_755),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_795),
.B(n_716),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_755),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_794),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_769),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_745),
.B(n_652),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_753),
.B(n_606),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_748),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_769),
.Y(n_846)
);

XNOR2x1_ASAP7_75t_L g847 ( 
.A(n_757),
.B(n_685),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_773),
.B(n_652),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_770),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_785),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_788),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_785),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_821),
.B(n_652),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_788),
.Y(n_855)
);

XOR2xp5_ASAP7_75t_L g856 ( 
.A(n_758),
.B(n_568),
.Y(n_856)
);

AND2x2_ASAP7_75t_SL g857 ( 
.A(n_781),
.B(n_694),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_809),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_789),
.B(n_659),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_778),
.B(n_708),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_818),
.B(n_791),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_801),
.B(n_716),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_730),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_811),
.B(n_716),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_742),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_782),
.B(n_703),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_818),
.B(n_653),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_738),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_766),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_768),
.Y(n_870)
);

XNOR2x2_ASAP7_75t_L g871 ( 
.A(n_793),
.B(n_614),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_793),
.B(n_719),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_804),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_746),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_775),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_790),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_797),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_802),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_778),
.B(n_720),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_805),
.B(n_723),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_756),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_806),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_816),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_761),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_752),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_819),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_776),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_804),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_817),
.B(n_666),
.Y(n_890)
);

XOR2xp5_ASAP7_75t_L g891 ( 
.A(n_812),
.B(n_574),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_666),
.Y(n_892)
);

INVx8_ASAP7_75t_L g893 ( 
.A(n_756),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_804),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_799),
.A2(n_622),
.B(n_602),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_814),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_815),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_784),
.B(n_601),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_803),
.B(n_615),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_762),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_762),
.Y(n_901)
);

XOR2xp5_ASAP7_75t_L g902 ( 
.A(n_743),
.B(n_577),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_763),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_808),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_729),
.B(n_728),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_736),
.Y(n_907)
);

OR2x2_ASAP7_75t_SL g908 ( 
.A(n_771),
.B(n_681),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_750),
.Y(n_909)
);

XOR2x2_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_678),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_739),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_754),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_786),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_772),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_907),
.B(n_694),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_823),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_825),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_896),
.B(n_696),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_796),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_827),
.B(n_800),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_881),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_873),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_841),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_881),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_827),
.B(n_800),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_826),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_828),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_854),
.B(n_798),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_843),
.B(n_787),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_833),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_888),
.B(n_734),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_844),
.B(n_783),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_874),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_861),
.B(n_732),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_897),
.B(n_696),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_836),
.B(n_741),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_835),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_861),
.B(n_807),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_843),
.B(n_780),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_841),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_874),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_857),
.B(n_820),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_857),
.B(n_704),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_886),
.B(n_813),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_906),
.B(n_704),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_895),
.A2(n_684),
.B(n_624),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_838),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_872),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_906),
.B(n_848),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_895),
.B(n_712),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_848),
.B(n_712),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_824),
.B(n_713),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_840),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_842),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_846),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_849),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_911),
.B(n_713),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_850),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_852),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_855),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_867),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_909),
.B(n_622),
.Y(n_962)
);

AND2x2_ASAP7_75t_SL g963 ( 
.A(n_862),
.B(n_624),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_901),
.B(n_633),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_824),
.B(n_697),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_887),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_822),
.B(n_737),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_863),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_829),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_860),
.A2(n_684),
.B(n_637),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_868),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_829),
.B(n_700),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_905),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_637),
.B(n_632),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_865),
.B(n_626),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_SL g976 ( 
.A(n_845),
.B(n_678),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_869),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_902),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_837),
.B(n_765),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_890),
.B(n_767),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_913),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_914),
.B(n_644),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_900),
.B(n_641),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_870),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_882),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_876),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_831),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_877),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_878),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_880),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_893),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_880),
.A2(n_646),
.B(n_632),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_866),
.B(n_644),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_837),
.B(n_687),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_903),
.B(n_630),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_839),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_904),
.B(n_760),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_864),
.B(n_656),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_832),
.B(n_578),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_879),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_883),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_884),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_889),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_873),
.B(n_682),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_859),
.B(n_741),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_893),
.Y(n_1006)
);

AND2x2_ASAP7_75t_SL g1007 ( 
.A(n_871),
.B(n_646),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_894),
.B(n_858),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_898),
.A2(n_718),
.B(n_695),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_899),
.B(n_644),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_873),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_912),
.B(n_847),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_892),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_908),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_891),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_923),
.B(n_687),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_940),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_969),
.B(n_999),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_991),
.Y(n_1019)
);

INVx6_ASAP7_75t_L g1020 ( 
.A(n_991),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_916),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_916),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_917),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_975),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_917),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_949),
.B(n_969),
.Y(n_1026)
);

AND2x6_ASAP7_75t_L g1027 ( 
.A(n_950),
.B(n_665),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_921),
.B(n_692),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_990),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_933),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_932),
.B(n_961),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_990),
.B(n_851),
.Y(n_1032)
);

BUFx4f_ASAP7_75t_L g1033 ( 
.A(n_990),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_985),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_973),
.B(n_777),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_931),
.B(n_777),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_965),
.B(n_853),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_965),
.B(n_834),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_985),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_933),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_926),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1014),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_990),
.Y(n_1044)
);

AND2x6_ASAP7_75t_L g1045 ( 
.A(n_950),
.B(n_665),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_934),
.B(n_830),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_981),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_975),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_933),
.B(n_641),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_1006),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_930),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_934),
.B(n_893),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_1003),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_973),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_964),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_924),
.B(n_972),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_999),
.B(n_856),
.Y(n_1057)
);

INVx6_ASAP7_75t_L g1058 ( 
.A(n_1006),
.Y(n_1058)
);

CKINVDCx11_ASAP7_75t_R g1059 ( 
.A(n_922),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_930),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_996),
.B(n_621),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_972),
.B(n_792),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_964),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_947),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1004),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_792),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_998),
.B(n_810),
.Y(n_1067)
);

BUFx4f_ASAP7_75t_L g1068 ( 
.A(n_962),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_964),
.B(n_643),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_947),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_953),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_998),
.B(n_810),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_962),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_974),
.B(n_692),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_996),
.B(n_657),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_1007),
.B(n_875),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_996),
.B(n_987),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_938),
.B(n_885),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_994),
.B(n_627),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_953),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1003),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_952),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_954),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1012),
.B(n_628),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_992),
.B(n_692),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_L g1086 ( 
.A(n_943),
.B(n_580),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_952),
.B(n_702),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_954),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_946),
.B(n_702),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_945),
.B(n_702),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_956),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_963),
.B(n_715),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_SL g1093 ( 
.A(n_920),
.B(n_910),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1032),
.A2(n_938),
.B1(n_963),
.B2(n_942),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_1044),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_1044),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1023),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_1059),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1043),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1033),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1016),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1025),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1030),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1044),
.Y(n_1104)
);

BUFx2_ASAP7_75t_SL g1105 ( 
.A(n_1019),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_1027),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1026),
.B(n_920),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1056),
.B(n_925),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_L g1109 ( 
.A(n_1027),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1056),
.B(n_925),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1030),
.Y(n_1111)
);

BUFx5_ASAP7_75t_L g1112 ( 
.A(n_1027),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1017),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1020),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1017),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1020),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1058),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1031),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1021),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1022),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_1082),
.B(n_995),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1026),
.B(n_1007),
.Y(n_1122)
);

INVxp67_ASAP7_75t_SL g1123 ( 
.A(n_1033),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1039),
.Y(n_1124)
);

BUFx2_ASAP7_75t_SL g1125 ( 
.A(n_1029),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1042),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1054),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1041),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1058),
.Y(n_1129)
);

INVx6_ASAP7_75t_L g1130 ( 
.A(n_1029),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1029),
.B(n_1012),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1041),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1081),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1060),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1034),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1081),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1081),
.B(n_1000),
.Y(n_1137)
);

BUFx24_ASAP7_75t_L g1138 ( 
.A(n_1035),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1040),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1051),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1054),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1050),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1075),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1053),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1065),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1080),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1082),
.B(n_995),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1018),
.B(n_951),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1037),
.Y(n_1149)
);

BUFx2_ASAP7_75t_SL g1150 ( 
.A(n_1035),
.Y(n_1150)
);

BUFx16f_ASAP7_75t_R g1151 ( 
.A(n_1069),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1088),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1068),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1077),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1038),
.B(n_970),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1064),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1053),
.B(n_1000),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1119),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1107),
.A2(n_1073),
.B1(n_1068),
.B2(n_1057),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1094),
.A2(n_1073),
.B1(n_929),
.B2(n_1047),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1149),
.B(n_1046),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_1114),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_1135),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1155),
.A2(n_1076),
.B1(n_1078),
.B2(n_1052),
.Y(n_1164)
);

BUFx8_ASAP7_75t_L g1165 ( 
.A(n_1098),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1097),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1155),
.A2(n_1015),
.B1(n_1076),
.B2(n_1084),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1098),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1120),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1149),
.A2(n_1052),
.B1(n_976),
.B2(n_1005),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1122),
.A2(n_1110),
.B1(n_1108),
.B2(n_1045),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1101),
.A2(n_1005),
.B1(n_1009),
.B2(n_936),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1097),
.Y(n_1173)
);

INVx6_ASAP7_75t_L g1174 ( 
.A(n_1114),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1124),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1127),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1122),
.A2(n_1027),
.B1(n_1045),
.B2(n_1062),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1154),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1102),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1108),
.A2(n_1110),
.B1(n_1148),
.B2(n_1147),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1126),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1116),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1121),
.B(n_1045),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1113),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1121),
.B(n_1045),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1121),
.A2(n_1047),
.B1(n_997),
.B2(n_928),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1147),
.A2(n_942),
.B1(n_979),
.B2(n_997),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1140),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1147),
.B(n_1024),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1143),
.A2(n_979),
.B1(n_1075),
.B2(n_1048),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1156),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1130),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1143),
.A2(n_919),
.B1(n_1077),
.B2(n_1092),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1102),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_1151),
.Y(n_1195)
);

OAI22x1_ASAP7_75t_L g1196 ( 
.A1(n_1131),
.A2(n_978),
.B1(n_1063),
.B2(n_1055),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1145),
.A2(n_1072),
.B1(n_1067),
.B2(n_1069),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1118),
.B(n_1145),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1113),
.A2(n_1036),
.B1(n_980),
.B2(n_1092),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1116),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1099),
.A2(n_1011),
.B1(n_1079),
.B2(n_939),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1134),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1117),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1134),
.Y(n_1204)
);

CKINVDCx11_ASAP7_75t_R g1205 ( 
.A(n_1139),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1115),
.A2(n_1004),
.B1(n_915),
.B2(n_1066),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1141),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1146),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1115),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1117),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1146),
.Y(n_1211)
);

BUFx4f_ASAP7_75t_SL g1212 ( 
.A(n_1129),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1130),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1153),
.A2(n_936),
.B1(n_612),
.B2(n_1011),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1129),
.B(n_1091),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1139),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1154),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1138),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1152),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1142),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1152),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1138),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1153),
.A2(n_1079),
.B1(n_1093),
.B2(n_635),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1164),
.A2(n_695),
.B1(n_1071),
.B2(n_1070),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1158),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1186),
.B(n_1150),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1160),
.A2(n_1083),
.B1(n_612),
.B2(n_1087),
.Y(n_1227)
);

OAI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1167),
.A2(n_1011),
.B1(n_1028),
.B2(n_1087),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1160),
.A2(n_1089),
.B1(n_1028),
.B2(n_1085),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1159),
.A2(n_1089),
.B1(n_1074),
.B2(n_1085),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1172),
.A2(n_1170),
.B1(n_1197),
.B2(n_1199),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1166),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1186),
.B(n_1142),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1214),
.A2(n_967),
.B(n_957),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1168),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1201),
.A2(n_915),
.B(n_918),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1165),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1161),
.A2(n_1123),
.B1(n_1100),
.B2(n_1109),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1173),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1159),
.A2(n_915),
.B1(n_1109),
.B2(n_1106),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1177),
.A2(n_1106),
.B1(n_1109),
.B2(n_1086),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1169),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1179),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1187),
.A2(n_1100),
.B1(n_1106),
.B2(n_1128),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1171),
.A2(n_927),
.B1(n_955),
.B2(n_937),
.Y(n_1245)
);

AOI211xp5_ASAP7_75t_L g1246 ( 
.A1(n_1223),
.A2(n_686),
.B(n_935),
.C(n_918),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1206),
.A2(n_1130),
.B1(n_1105),
.B2(n_1125),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1180),
.A2(n_958),
.B1(n_959),
.B2(n_956),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1192),
.B(n_1095),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1175),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1180),
.A2(n_960),
.B1(n_1079),
.B2(n_977),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1181),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1196),
.A2(n_1135),
.B1(n_640),
.B2(n_1013),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1183),
.A2(n_960),
.B1(n_984),
.B2(n_968),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1183),
.A2(n_989),
.B1(n_1001),
.B2(n_988),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1165),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1190),
.A2(n_1074),
.B1(n_661),
.B2(n_663),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1185),
.A2(n_986),
.B1(n_971),
.B2(n_1112),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1205),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1188),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1185),
.A2(n_986),
.B1(n_971),
.B2(n_1112),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1191),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1202),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1213),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1216),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1218),
.A2(n_1112),
.B1(n_1130),
.B2(n_1154),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1198),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1204),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1163),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1208),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1209),
.A2(n_1154),
.B1(n_1061),
.B2(n_983),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1193),
.A2(n_1112),
.B1(n_966),
.B2(n_1090),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1189),
.B(n_918),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1176),
.A2(n_1090),
.B(n_1013),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1218),
.A2(n_1112),
.B1(n_1154),
.B2(n_1111),
.Y(n_1275)
);

OAI222xp33_ASAP7_75t_L g1276 ( 
.A1(n_1222),
.A2(n_582),
.B1(n_586),
.B2(n_588),
.C1(n_590),
.C2(n_594),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1193),
.A2(n_1112),
.B1(n_987),
.B2(n_1002),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1207),
.A2(n_982),
.B(n_993),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1184),
.B(n_935),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1222),
.A2(n_1215),
.B1(n_1112),
.B2(n_1220),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1215),
.A2(n_987),
.B1(n_1002),
.B2(n_1000),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1219),
.A2(n_661),
.B1(n_663),
.B2(n_653),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1220),
.A2(n_1096),
.B1(n_1144),
.B2(n_1111),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1174),
.B(n_935),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1221),
.A2(n_661),
.B1(n_663),
.B2(n_653),
.Y(n_1285)
);

CKINVDCx8_ASAP7_75t_R g1286 ( 
.A(n_1162),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1194),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1211),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1178),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1231),
.A2(n_1195),
.B1(n_690),
.B2(n_688),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1227),
.A2(n_690),
.B1(n_683),
.B2(n_670),
.Y(n_1291)
);

OAI221xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1234),
.A2(n_1210),
.B1(n_1182),
.B2(n_1200),
.C(n_1010),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1267),
.B(n_1178),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1232),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1253),
.B(n_1217),
.Y(n_1295)
);

OAI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1227),
.A2(n_1061),
.B1(n_1008),
.B2(n_983),
.C(n_1203),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1224),
.A2(n_670),
.B1(n_660),
.B2(n_715),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1224),
.A2(n_670),
.B1(n_660),
.B2(n_715),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1233),
.B(n_1217),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1279),
.B(n_1213),
.Y(n_1300)
);

CKINVDCx11_ASAP7_75t_R g1301 ( 
.A(n_1265),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1228),
.A2(n_1002),
.B1(n_1003),
.B2(n_948),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1228),
.A2(n_727),
.B1(n_726),
.B2(n_721),
.C(n_596),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1251),
.A2(n_1003),
.B1(n_948),
.B2(n_1192),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1213),
.Y(n_1305)
);

AOI222xp33_ASAP7_75t_L g1306 ( 
.A1(n_1276),
.A2(n_595),
.B1(n_680),
.B2(n_675),
.C1(n_666),
.C2(n_668),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1226),
.A2(n_948),
.B1(n_1163),
.B2(n_1144),
.Y(n_1307)
);

OAI222xp33_ASAP7_75t_L g1308 ( 
.A1(n_1247),
.A2(n_1257),
.B1(n_1280),
.B2(n_1238),
.C1(n_1266),
.C2(n_1245),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1239),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1246),
.A2(n_1212),
.B1(n_1174),
.B2(n_1203),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1225),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1286),
.A2(n_1137),
.B1(n_1157),
.B2(n_1096),
.Y(n_1312)
);

INVxp67_ASAP7_75t_SL g1313 ( 
.A(n_1283),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1243),
.B(n_1104),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1240),
.A2(n_1137),
.B1(n_1157),
.B2(n_1096),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1287),
.B(n_1104),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1274),
.A2(n_1144),
.B1(n_1111),
.B2(n_1132),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1244),
.A2(n_1096),
.B1(n_1132),
.B2(n_1103),
.Y(n_1318)
);

OAI221xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1236),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.C(n_38),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1288),
.B(n_1104),
.Y(n_1320)
);

OAI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1255),
.A2(n_1137),
.B1(n_1157),
.B2(n_941),
.C(n_727),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1242),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1254),
.A2(n_1096),
.B1(n_1132),
.B2(n_1103),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1250),
.B(n_1104),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1248),
.A2(n_1103),
.B1(n_1104),
.B2(n_726),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1257),
.A2(n_727),
.B1(n_726),
.B2(n_721),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1252),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1260),
.B(n_1133),
.Y(n_1328)
);

OAI222xp33_ASAP7_75t_L g1329 ( 
.A1(n_1275),
.A2(n_668),
.B1(n_675),
.B2(n_680),
.C1(n_625),
.C2(n_621),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1229),
.A2(n_721),
.B1(n_675),
.B2(n_680),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1241),
.A2(n_1136),
.B1(n_1133),
.B2(n_1049),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1271),
.A2(n_1136),
.B1(n_1133),
.B2(n_668),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1229),
.A2(n_625),
.B(n_36),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1284),
.A2(n_1136),
.B1(n_1133),
.B2(n_644),
.Y(n_1334)
);

OAI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1278),
.A2(n_1136),
.B(n_1133),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1269),
.B(n_1259),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1262),
.B(n_1136),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1230),
.A2(n_38),
.B1(n_41),
.B2(n_44),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1263),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1230),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1237),
.A2(n_1049),
.B1(n_639),
.B2(n_629),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1272),
.A2(n_1277),
.B(n_1282),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1235),
.A2(n_629),
.B1(n_618),
.B2(n_616),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1268),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1270),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1258),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1256),
.A2(n_639),
.B1(n_629),
.B2(n_618),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1289),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1283),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1249),
.B(n_54),
.Y(n_1350)
);

NOR3xp33_ASAP7_75t_L g1351 ( 
.A(n_1249),
.B(n_1261),
.C(n_1282),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1281),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1264),
.A2(n_639),
.B1(n_618),
.B2(n_616),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1264),
.B(n_56),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1264),
.A2(n_616),
.B1(n_610),
.B2(n_61),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1293),
.B(n_1264),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1300),
.B(n_1285),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1306),
.B(n_1290),
.C(n_1338),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1290),
.A2(n_1285),
.B1(n_610),
.B2(n_61),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1319),
.A2(n_610),
.B1(n_60),
.B2(n_62),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_58),
.C(n_62),
.Y(n_1361)
);

NOR3xp33_ASAP7_75t_L g1362 ( 
.A(n_1292),
.B(n_64),
.C(n_66),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1305),
.B(n_1322),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1340),
.B(n_64),
.C(n_66),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1340),
.B(n_67),
.C(n_68),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1299),
.B(n_67),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1335),
.A2(n_68),
.B(n_69),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1327),
.B(n_70),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1311),
.B(n_71),
.Y(n_1369)
);

AOI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1344),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.C(n_74),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1339),
.B(n_72),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1348),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1295),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1294),
.B(n_75),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1308),
.B(n_76),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1309),
.B(n_80),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1324),
.B(n_83),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1337),
.B(n_1316),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1344),
.B(n_84),
.C(n_85),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1350),
.B(n_371),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1328),
.B(n_86),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1296),
.B(n_1313),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1297),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1349),
.B(n_1354),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1345),
.A2(n_90),
.B1(n_91),
.B2(n_99),
.C(n_101),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1320),
.B(n_104),
.Y(n_1386)
);

OAI21xp33_ASAP7_75t_L g1387 ( 
.A1(n_1345),
.A2(n_105),
.B(n_106),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1314),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1307),
.B(n_1291),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1303),
.B(n_108),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1297),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1291),
.B(n_114),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1342),
.A2(n_1302),
.B(n_1330),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1318),
.B(n_115),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1352),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1352),
.A2(n_123),
.B(n_125),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1346),
.A2(n_126),
.B1(n_128),
.B2(n_131),
.C(n_142),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1346),
.B(n_1351),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1333),
.B(n_143),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1298),
.B(n_144),
.Y(n_1400)
);

AOI211xp5_ASAP7_75t_L g1401 ( 
.A1(n_1310),
.A2(n_145),
.B(n_148),
.C(n_149),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1332),
.B(n_368),
.Y(n_1402)
);

OAI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1298),
.A2(n_151),
.B(n_154),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1312),
.B(n_1317),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1330),
.B(n_157),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1341),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1304),
.B(n_166),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1336),
.B(n_1315),
.Y(n_1408)
);

OAI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1355),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.C(n_172),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_L g1410 ( 
.A(n_1329),
.B(n_180),
.C(n_182),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1325),
.B(n_366),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1343),
.B(n_184),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1372),
.Y(n_1413)
);

NOR2x1_ASAP7_75t_L g1414 ( 
.A(n_1367),
.B(n_1321),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1378),
.B(n_1331),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1362),
.A2(n_1347),
.B1(n_1323),
.B2(n_1334),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1372),
.B(n_1363),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1356),
.B(n_1301),
.Y(n_1418)
);

NAND4xp75_ASAP7_75t_L g1419 ( 
.A(n_1375),
.B(n_1353),
.C(n_1326),
.D(n_191),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1388),
.B(n_1326),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1408),
.B(n_185),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1382),
.Y(n_1422)
);

OAI211xp5_ASAP7_75t_L g1423 ( 
.A1(n_1375),
.A2(n_187),
.B(n_192),
.C(n_195),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1384),
.B(n_197),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1362),
.B(n_198),
.C(n_199),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1404),
.B(n_1368),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_200),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1381),
.B(n_1380),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1357),
.B(n_201),
.Y(n_1429)
);

NAND4xp25_ASAP7_75t_L g1430 ( 
.A(n_1370),
.B(n_204),
.C(n_205),
.D(n_208),
.Y(n_1430)
);

NAND4xp75_ASAP7_75t_L g1431 ( 
.A(n_1398),
.B(n_212),
.C(n_218),
.D(n_219),
.Y(n_1431)
);

NOR3xp33_ASAP7_75t_L g1432 ( 
.A(n_1358),
.B(n_220),
.C(n_221),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1385),
.B(n_222),
.C(n_227),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1390),
.A2(n_363),
.B(n_229),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1367),
.Y(n_1435)
);

OAI211xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1373),
.A2(n_228),
.B(n_230),
.C(n_232),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1369),
.Y(n_1437)
);

NAND4xp75_ASAP7_75t_L g1438 ( 
.A(n_1390),
.B(n_236),
.C(n_238),
.D(n_241),
.Y(n_1438)
);

OAI211xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1387),
.A2(n_244),
.B(n_245),
.C(n_247),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1366),
.B(n_249),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1371),
.B(n_251),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_252),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_SL g1443 ( 
.A(n_1394),
.B(n_1402),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_R g1444 ( 
.A(n_1404),
.B(n_254),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1361),
.B(n_1365),
.C(n_1364),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1386),
.B(n_255),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1379),
.B(n_257),
.C(n_258),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1376),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1417),
.B(n_1393),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1413),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1435),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1437),
.Y(n_1454)
);

XNOR2xp5_ASAP7_75t_L g1455 ( 
.A(n_1418),
.B(n_1360),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1422),
.B(n_1393),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1449),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1426),
.B(n_1401),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1445),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1420),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1445),
.B(n_1428),
.Y(n_1462)
);

INVx5_ASAP7_75t_L g1463 ( 
.A(n_1421),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1429),
.B(n_1389),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1414),
.B(n_1399),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1420),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1432),
.A2(n_1397),
.B1(n_1410),
.B2(n_1395),
.Y(n_1467)
);

NAND4xp75_ASAP7_75t_L g1468 ( 
.A(n_1434),
.B(n_1411),
.C(n_1405),
.D(n_1392),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1440),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1427),
.B(n_1396),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1427),
.B(n_1440),
.Y(n_1471)
);

XOR2xp5_ASAP7_75t_L g1472 ( 
.A(n_1424),
.B(n_1406),
.Y(n_1472)
);

XOR2x2_ASAP7_75t_L g1473 ( 
.A(n_1455),
.B(n_1446),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1453),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1462),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_R g1476 ( 
.A(n_1463),
.B(n_1444),
.Y(n_1476)
);

XOR2x2_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1432),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1469),
.B(n_1443),
.Y(n_1478)
);

XOR2xp5_ASAP7_75t_L g1479 ( 
.A(n_1472),
.B(n_1419),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1460),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1451),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1460),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1451),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1454),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1471),
.B(n_1441),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1457),
.B(n_1416),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1454),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1475),
.Y(n_1488)
);

XOR2x2_ASAP7_75t_L g1489 ( 
.A(n_1473),
.B(n_1470),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1477),
.A2(n_1467),
.B1(n_1468),
.B2(n_1425),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1480),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1479),
.A2(n_1468),
.B1(n_1465),
.B2(n_1459),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1482),
.Y(n_1493)
);

XNOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1486),
.B(n_1462),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1478),
.A2(n_1459),
.B1(n_1452),
.B2(n_1456),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1481),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1484),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1483),
.Y(n_1498)
);

XNOR2xp5_ASAP7_75t_L g1499 ( 
.A(n_1476),
.B(n_1472),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1487),
.Y(n_1500)
);

AOI22x1_ASAP7_75t_L g1501 ( 
.A1(n_1474),
.A2(n_1453),
.B1(n_1452),
.B2(n_1466),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1474),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1478),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1498),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1498),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1497),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1500),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1492),
.A2(n_1430),
.B1(n_1433),
.B2(n_1457),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1488),
.Y(n_1509)
);

OAI322xp33_ASAP7_75t_L g1510 ( 
.A1(n_1490),
.A2(n_1466),
.A3(n_1461),
.B1(n_1485),
.B2(n_1458),
.C1(n_1450),
.C2(n_1460),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1490),
.Y(n_1511)
);

OAI322xp33_ASAP7_75t_L g1512 ( 
.A1(n_1499),
.A2(n_1485),
.A3(n_1458),
.B1(n_1450),
.B2(n_1359),
.C1(n_1464),
.C2(n_1442),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1489),
.A2(n_1503),
.B1(n_1494),
.B2(n_1495),
.Y(n_1513)
);

OAI322xp33_ASAP7_75t_L g1514 ( 
.A1(n_1511),
.A2(n_1513),
.A3(n_1504),
.B1(n_1505),
.B2(n_1507),
.C1(n_1506),
.C2(n_1509),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1511),
.A2(n_1491),
.B1(n_1493),
.B2(n_1496),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1512),
.A2(n_1502),
.B1(n_1423),
.B2(n_1436),
.C(n_1439),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1508),
.A2(n_1423),
.B1(n_1431),
.B2(n_1438),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1510),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1511),
.A2(n_1464),
.B1(n_1436),
.B2(n_1463),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1511),
.A2(n_1463),
.B1(n_1439),
.B2(n_1448),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1515),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1518),
.A2(n_1501),
.B1(n_1463),
.B2(n_1395),
.Y(n_1522)
);

OAI22x1_ASAP7_75t_L g1523 ( 
.A1(n_1517),
.A2(n_1520),
.B1(n_1519),
.B2(n_1501),
.Y(n_1523)
);

AO22x2_ASAP7_75t_L g1524 ( 
.A1(n_1514),
.A2(n_1410),
.B1(n_1447),
.B2(n_1383),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1516),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1515),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1521),
.B(n_1526),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1525),
.B(n_1463),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1523),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1522),
.B(n_1403),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1524),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1521),
.Y(n_1532)
);

AOI31xp33_ASAP7_75t_L g1533 ( 
.A1(n_1521),
.A2(n_1409),
.A3(n_1391),
.B(n_1407),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1528),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1529),
.A2(n_1400),
.B1(n_261),
.B2(n_264),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1531),
.A2(n_260),
.B1(n_266),
.B2(n_268),
.Y(n_1536)
);

NOR2x1_ASAP7_75t_L g1537 ( 
.A(n_1527),
.B(n_269),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1530),
.A2(n_270),
.B1(n_271),
.B2(n_276),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1532),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1535),
.A2(n_1530),
.B1(n_1533),
.B2(n_280),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1539),
.Y(n_1541)
);

AND5x1_ASAP7_75t_L g1542 ( 
.A(n_1536),
.B(n_361),
.C(n_278),
.D(n_281),
.E(n_283),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1538),
.B2(n_285),
.Y(n_1543)
);

NOR4xp75_ASAP7_75t_L g1544 ( 
.A(n_1534),
.B(n_277),
.C(n_284),
.D(n_286),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1541),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1544),
.Y(n_1546)
);

AND3x4_ASAP7_75t_L g1547 ( 
.A(n_1540),
.B(n_289),
.C(n_293),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1543),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1542),
.Y(n_1549)
);

OAI22x1_ASAP7_75t_L g1550 ( 
.A1(n_1547),
.A2(n_294),
.B1(n_297),
.B2(n_299),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1545),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1546),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1549),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_1553)
);

AO22x2_ASAP7_75t_L g1554 ( 
.A1(n_1548),
.A2(n_357),
.B1(n_307),
.B2(n_309),
.Y(n_1554)
);

NAND4xp75_ASAP7_75t_L g1555 ( 
.A(n_1545),
.B(n_306),
.C(n_311),
.D(n_312),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1551),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1552),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1553),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1554),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1557),
.A2(n_1558),
.B1(n_1559),
.B2(n_1550),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1558),
.A2(n_1555),
.B1(n_317),
.B2(n_318),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1560),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1561),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1562),
.A2(n_1556),
.B1(n_319),
.B2(n_323),
.Y(n_1564)
);

AOI211xp5_ASAP7_75t_L g1565 ( 
.A1(n_1563),
.A2(n_1556),
.B(n_326),
.C(n_330),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1565),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1566),
.A2(n_1564),
.B1(n_332),
.B2(n_334),
.C(n_337),
.Y(n_1567)
);

AOI211xp5_ASAP7_75t_L g1568 ( 
.A1(n_1567),
.A2(n_314),
.B(n_338),
.C(n_339),
.Y(n_1568)
);


endmodule