module fake_netlist_5_761_n_1505 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1505);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1505;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_1058;
wire n_586;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_259),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_60),
.Y(n_391)
);

CKINVDCx12_ASAP7_75t_R g392 ( 
.A(n_356),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_304),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_286),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_96),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_180),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_323),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_140),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_15),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_281),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_33),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_146),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_296),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_258),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_279),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_225),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_341),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_49),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_70),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_151),
.Y(n_414)
);

BUFx8_ASAP7_75t_SL g415 ( 
.A(n_334),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_175),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_126),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_347),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_357),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_178),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_60),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_270),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_69),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_23),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_128),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_384),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_166),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_333),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_65),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_43),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_2),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_121),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_163),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_202),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_37),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_231),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_63),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_236),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_179),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_50),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_112),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_212),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_309),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_111),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_16),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_348),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_331),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_294),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_311),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_199),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_90),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_120),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_78),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_282),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_379),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_251),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_361),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_69),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_226),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_328),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_161),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_297),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_210),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_154),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_265),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_368),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_147),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_81),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_93),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_268),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_66),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_233),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_176),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_170),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_256),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_84),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_321),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_81),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_300),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_247),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_274),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_222),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_12),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_293),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_167),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_86),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_374),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_92),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_208),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_192),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_153),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_125),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_239),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_327),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_19),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_337),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_380),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_322),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_22),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_143),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_291),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_349),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_302),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_365),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_189),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_16),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_55),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_359),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_12),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_6),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_346),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_336),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_377),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_173),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_370),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_201),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_98),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_24),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_73),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_340),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_307),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_35),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_366),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_254),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_353),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_39),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_14),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_95),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_40),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_264),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_227),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_195),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_299),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_160),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_41),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_7),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_308),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_40),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_271),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_375),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_267),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_385),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_102),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_188),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_118),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_276),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_358),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_109),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_27),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_64),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_53),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_250),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_193),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_75),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_292),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_87),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_78),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_10),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_132),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_103),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_30),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_138),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_262),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_76),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_316),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_85),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_242),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_382),
.Y(n_571)
);

CKINVDCx11_ASAP7_75t_R g572 ( 
.A(n_53),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_59),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_3),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_216),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_343),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_344),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_35),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_181),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_15),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_475),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_471),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_475),
.B(n_0),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_424),
.B(n_0),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_424),
.B(n_1),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_437),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_393),
.B(n_1),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_507),
.B(n_2),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_3),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_417),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_424),
.B(n_4),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_393),
.B(n_4),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

BUFx8_ASAP7_75t_L g598 ( 
.A(n_527),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_524),
.B(n_5),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_424),
.B(n_494),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_417),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_471),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_524),
.B(n_5),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_417),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_515),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_530),
.B(n_6),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_494),
.B(n_7),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_515),
.B(n_88),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_542),
.B(n_8),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_479),
.B(n_8),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_479),
.B(n_9),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_530),
.B(n_9),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_420),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_542),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_412),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_420),
.Y(n_622)
);

BUFx8_ASAP7_75t_SL g623 ( 
.A(n_510),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_479),
.B(n_10),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_404),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_391),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_421),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_398),
.B(n_89),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_559),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_432),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_510),
.Y(n_631)
);

BUFx8_ASAP7_75t_SL g632 ( 
.A(n_425),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_388),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_448),
.B(n_11),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_420),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_433),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_509),
.B(n_11),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_414),
.B(n_441),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_398),
.B(n_13),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_415),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_411),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_473),
.B(n_13),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_412),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_409),
.B(n_453),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_459),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_443),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_415),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_473),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_389),
.B(n_408),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_483),
.B(n_14),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_502),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_427),
.B(n_17),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_394),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_483),
.B(n_17),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_497),
.B(n_528),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_399),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_413),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_412),
.B(n_18),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_512),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_401),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_513),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_521),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_497),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_481),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_481),
.B(n_18),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_450),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_405),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_472),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_390),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_481),
.B(n_19),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_525),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_529),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_552),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_553),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_464),
.B(n_20),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_565),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_478),
.B(n_20),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_565),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_431),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_466),
.B(n_21),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_585),
.A2(n_574),
.B1(n_578),
.B2(n_573),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_508),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_638),
.A2(n_460),
.B1(n_493),
.B2(n_459),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_649),
.B(n_526),
.Y(n_685)
);

OA22x2_ASAP7_75t_L g686 ( 
.A1(n_584),
.A2(n_439),
.B1(n_461),
.B2(n_456),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_589),
.A2(n_493),
.B1(n_534),
.B2(n_460),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_596),
.A2(n_534),
.B1(n_400),
.B2(n_500),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_633),
.B(n_395),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_L g690 ( 
.A1(n_681),
.A2(n_564),
.B1(n_402),
.B2(n_486),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_681),
.A2(n_489),
.B1(n_498),
.B2(n_474),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_617),
.A2(n_580),
.B1(n_532),
.B2(n_538),
.Y(n_692)
);

AOI22x1_ASAP7_75t_SL g693 ( 
.A1(n_623),
.A2(n_522),
.B1(n_541),
.B2(n_539),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_581),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_652),
.A2(n_447),
.B1(n_568),
.B2(n_557),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_667),
.B(n_396),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_652),
.A2(n_560),
.B1(n_561),
.B2(n_554),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_625),
.B(n_540),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_SL g699 ( 
.A1(n_617),
.A2(n_569),
.B1(n_567),
.B2(n_397),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_617),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_676),
.A2(n_392),
.B1(n_407),
.B2(n_406),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_676),
.A2(n_410),
.B1(n_418),
.B2(n_416),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_641),
.Y(n_703)
);

OA22x2_ASAP7_75t_L g704 ( 
.A1(n_626),
.A2(n_423),
.B1(n_434),
.B2(n_403),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_R g706 ( 
.A1(n_678),
.A2(n_436),
.B1(n_445),
.B2(n_435),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_658),
.B(n_419),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_657),
.B(n_422),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_581),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_640),
.B(n_647),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_643),
.A2(n_457),
.B1(n_465),
.B2(n_455),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_SL g713 ( 
.A1(n_617),
.A2(n_480),
.B1(n_485),
.B2(n_470),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_601),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_622),
.A2(n_501),
.B1(n_504),
.B2(n_495),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_640),
.B(n_647),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_622),
.B(n_506),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_644),
.A2(n_428),
.B1(n_429),
.B2(n_426),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_632),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_648),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_SL g721 ( 
.A1(n_645),
.A2(n_517),
.B1(n_519),
.B2(n_514),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_430),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_665),
.B(n_523),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_678),
.A2(n_440),
.B1(n_442),
.B2(n_438),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_647),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_644),
.A2(n_446),
.B1(n_449),
.B2(n_444),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_601),
.Y(n_727)
);

AO22x2_ASAP7_75t_L g728 ( 
.A1(n_585),
.A2(n_535),
.B1(n_544),
.B2(n_533),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_643),
.A2(n_650),
.B1(n_642),
.B2(n_622),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_618),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_648),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_680),
.A2(n_452),
.B1(n_454),
.B2(n_451),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_SL g733 ( 
.A1(n_583),
.A2(n_570),
.B1(n_575),
.B2(n_555),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_653),
.B(n_656),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_590),
.A2(n_579),
.B1(n_23),
.B2(n_21),
.Y(n_735)
);

AO22x2_ASAP7_75t_L g736 ( 
.A1(n_590),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_SL g737 ( 
.A1(n_591),
.A2(n_462),
.B1(n_463),
.B2(n_458),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_670),
.A2(n_468),
.B1(n_469),
.B2(n_467),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_599),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_621),
.B(n_26),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_601),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_664),
.A2(n_477),
.B1(n_482),
.B2(n_476),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_647),
.B(n_484),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_648),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_601),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_599),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_609),
.A2(n_488),
.B1(n_490),
.B2(n_487),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_603),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_622),
.A2(n_492),
.B1(n_496),
.B2(n_491),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_635),
.A2(n_503),
.B1(n_505),
.B2(n_499),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_609),
.A2(n_516),
.B1(n_518),
.B2(n_511),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_602),
.B(n_31),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_SL g754 ( 
.A1(n_635),
.A2(n_531),
.B1(n_536),
.B2(n_520),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_582),
.B(n_537),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_SL g756 ( 
.A1(n_642),
.A2(n_650),
.B1(n_612),
.B2(n_624),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_648),
.Y(n_757)
);

AOI22x1_ASAP7_75t_L g758 ( 
.A1(n_655),
.A2(n_545),
.B1(n_546),
.B2(n_543),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_L g759 ( 
.A1(n_635),
.A2(n_548),
.B1(n_549),
.B2(n_547),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_604),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_635),
.A2(n_551),
.B1(n_556),
.B2(n_550),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_598),
.A2(n_562),
.B1(n_563),
.B2(n_558),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_592),
.B(n_566),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_593),
.A2(n_576),
.B1(n_577),
.B2(n_571),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_604),
.Y(n_765)
);

AO22x2_ASAP7_75t_L g766 ( 
.A1(n_603),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_593),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_720),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_731),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_744),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_757),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_730),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_709),
.Y(n_773)
);

XOR2xp5_ASAP7_75t_L g774 ( 
.A(n_719),
.B(n_632),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_755),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_756),
.B(n_605),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_763),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_709),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_710),
.Y(n_779)
);

BUFx5_ASAP7_75t_L g780 ( 
.A(n_711),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_710),
.Y(n_781)
);

BUFx6f_ASAP7_75t_SL g782 ( 
.A(n_740),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_727),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_727),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_694),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_700),
.B(n_594),
.Y(n_786)
);

XOR2xp5_ASAP7_75t_L g787 ( 
.A(n_684),
.B(n_626),
.Y(n_787)
);

XOR2xp5_ASAP7_75t_L g788 ( 
.A(n_688),
.B(n_636),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_705),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_714),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_741),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_683),
.B(n_619),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_745),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_748),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_760),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_765),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_753),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_704),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_717),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_682),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_653),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_708),
.B(n_611),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_698),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_689),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_696),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_728),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_767),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_728),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_703),
.B(n_619),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_723),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_697),
.B(n_656),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_686),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_729),
.B(n_614),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_758),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_718),
.B(n_660),
.Y(n_816)
);

XNOR2xp5_ASAP7_75t_L g817 ( 
.A(n_687),
.B(n_695),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_726),
.B(n_660),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_758),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_722),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_734),
.B(n_620),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_702),
.B(n_602),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_747),
.A2(n_615),
.B(n_612),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_743),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_766),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_766),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_716),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_736),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_736),
.Y(n_829)
);

XNOR2xp5_ASAP7_75t_L g830 ( 
.A(n_693),
.B(n_611),
.Y(n_830)
);

INVx4_ASAP7_75t_SL g831 ( 
.A(n_725),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_739),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_701),
.B(n_608),
.Y(n_833)
);

XNOR2x2_ASAP7_75t_L g834 ( 
.A(n_739),
.B(n_623),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_742),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_712),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_764),
.B(n_600),
.Y(n_837)
);

INVx4_ASAP7_75t_SL g838 ( 
.A(n_740),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_746),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_724),
.B(n_752),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_749),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_721),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_735),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_735),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_707),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_749),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_713),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_715),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_738),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_750),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_759),
.B(n_666),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_690),
.B(n_600),
.Y(n_853)
);

BUFx5_ASAP7_75t_L g854 ( 
.A(n_751),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_691),
.Y(n_855)
);

CKINVDCx14_ASAP7_75t_R g856 ( 
.A(n_737),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_733),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_732),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_754),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_796),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_805),
.B(n_666),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_792),
.B(n_634),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_785),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_819),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_804),
.B(n_762),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_806),
.B(n_637),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_803),
.B(n_588),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_803),
.B(n_588),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_790),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_821),
.B(n_666),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_824),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_791),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_793),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_797),
.B(n_811),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_794),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_801),
.B(n_597),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_818),
.B(n_761),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_823),
.B(n_597),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_669),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_821),
.B(n_666),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_841),
.B(n_692),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_810),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_856),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_831),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_799),
.B(n_668),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_768),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_798),
.B(n_669),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_769),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_835),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_822),
.B(n_776),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_831),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_770),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_772),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_815),
.B(n_668),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_771),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_616),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_773),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_837),
.B(n_668),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_827),
.B(n_837),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_775),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_778),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_779),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_781),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_813),
.A2(n_706),
.B1(n_624),
.B2(n_615),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_788),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_850),
.B(n_598),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_783),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_816),
.B(n_631),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_784),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_808),
.B(n_655),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_808),
.B(n_636),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_777),
.B(n_668),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_859),
.B(n_631),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_814),
.B(n_663),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_814),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_807),
.B(n_639),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_825),
.B(n_826),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_848),
.B(n_663),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_780),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_859),
.B(n_618),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_849),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_800),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_802),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_833),
.B(n_639),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_812),
.B(n_833),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_780),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_780),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_853),
.B(n_618),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_836),
.B(n_663),
.Y(n_933)
);

AND2x2_ASAP7_75t_SL g934 ( 
.A(n_851),
.B(n_654),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_780),
.B(n_852),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_809),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_844),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_780),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_855),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_853),
.B(n_654),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_854),
.B(n_663),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_786),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_854),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_860),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_854),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_854),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_860),
.B(n_651),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_851),
.B(n_618),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_845),
.B(n_627),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_858),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_828),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_829),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_832),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_857),
.B(n_629),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_839),
.B(n_630),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_840),
.B(n_646),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_842),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_847),
.B(n_628),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_846),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_890),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_879),
.B(n_817),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_892),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_887),
.B(n_843),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_894),
.B(n_929),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_919),
.B(n_787),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_871),
.B(n_838),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_887),
.B(n_830),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_890),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_919),
.B(n_677),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_882),
.B(n_677),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_899),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_899),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_871),
.B(n_874),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_887),
.Y(n_976)
);

NOR2x1_ASAP7_75t_L g977 ( 
.A(n_895),
.B(n_786),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_874),
.B(n_838),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_897),
.B(n_672),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_882),
.B(n_677),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_872),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_880),
.B(n_834),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_894),
.B(n_782),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_943),
.B(n_677),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_895),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_939),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_921),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_879),
.B(n_659),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_915),
.B(n_774),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_897),
.B(n_673),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_924),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_921),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_915),
.B(n_661),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_895),
.B(n_662),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_904),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_944),
.B(n_604),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_896),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_893),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_914),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_893),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_921),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_914),
.B(n_671),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_872),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_896),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_869),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_943),
.B(n_628),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_947),
.B(n_674),
.Y(n_1007)
);

BUFx4f_ASAP7_75t_L g1008 ( 
.A(n_921),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_904),
.Y(n_1009)
);

INVx5_ASAP7_75t_L g1010 ( 
.A(n_938),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_869),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_875),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_949),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_949),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_944),
.B(n_938),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_945),
.B(n_628),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_881),
.B(n_629),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_921),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_875),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_921),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_881),
.B(n_629),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_947),
.B(n_629),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_947),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_937),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_937),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_945),
.B(n_946),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_944),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_868),
.B(n_706),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_864),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_878),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_953),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_946),
.B(n_950),
.Y(n_1032)
);

NAND2x1_ASAP7_75t_L g1033 ( 
.A(n_938),
.B(n_610),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_951),
.B(n_91),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_886),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_951),
.B(n_94),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_923),
.B(n_606),
.Y(n_1037)
);

BUFx8_ASAP7_75t_L g1038 ( 
.A(n_1035),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_1026),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_998),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_1008),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_986),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_1008),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_962),
.A2(n_982),
.B1(n_966),
.B2(n_884),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1024),
.Y(n_1046)
);

CKINVDCx8_ASAP7_75t_R g1047 ( 
.A(n_1000),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_1005),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_991),
.B(n_863),
.Y(n_1049)
);

BUFx2_ASAP7_75t_SL g1050 ( 
.A(n_967),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_966),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_961),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_975),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_976),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_969),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1032),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_963),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_997),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_970),
.Y(n_1060)
);

BUFx8_ASAP7_75t_SL g1061 ( 
.A(n_964),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1004),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_976),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_991),
.B(n_863),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_985),
.B(n_1027),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1027),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1029),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_983),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_982),
.A2(n_903),
.B1(n_934),
.B2(n_912),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_967),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_983),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_985),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_989),
.Y(n_1073)
);

BUFx4_ASAP7_75t_SL g1074 ( 
.A(n_964),
.Y(n_1074)
);

BUFx2_ASAP7_75t_SL g1075 ( 
.A(n_978),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1013),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1014),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_1010),
.B(n_950),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_973),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_974),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1031),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_999),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_978),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1031),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_964),
.B(n_960),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_981),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_986),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1003),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_1023),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_965),
.A2(n_903),
.B1(n_935),
.B2(n_934),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_1005),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_995),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1007),
.B(n_928),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1025),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_995),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_994),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_999),
.B(n_900),
.Y(n_1097)
);

BUFx4f_ASAP7_75t_L g1098 ( 
.A(n_994),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1011),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1012),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1028),
.A2(n_934),
.B1(n_948),
.B2(n_928),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1019),
.Y(n_1102)
);

BUFx4_ASAP7_75t_SL g1103 ( 
.A(n_994),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1058),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1045),
.A2(n_917),
.B1(n_960),
.B2(n_910),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_1039),
.B(n_1010),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1040),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1042),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1058),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1097),
.B(n_1002),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_SL g1111 ( 
.A1(n_1051),
.A2(n_900),
.B1(n_693),
.B2(n_940),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1049),
.B(n_988),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1069),
.A2(n_993),
.B1(n_908),
.B2(n_925),
.Y(n_1113)
);

CKINVDCx11_ASAP7_75t_R g1114 ( 
.A(n_1047),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1052),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1048),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1064),
.B(n_940),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1055),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1060),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1059),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_1038),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1062),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_1038),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1040),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1067),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1101),
.A2(n_908),
.B1(n_932),
.B2(n_925),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1042),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1041),
.A2(n_1021),
.B1(n_1017),
.B2(n_992),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_1096),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1076),
.A2(n_587),
.B1(n_595),
.B2(n_586),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1077),
.A2(n_587),
.B1(n_595),
.B2(n_586),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1046),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1041),
.A2(n_1001),
.B1(n_1018),
.B2(n_987),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1090),
.A2(n_877),
.B1(n_1036),
.B2(n_1034),
.Y(n_1134)
);

INVx6_ASAP7_75t_L g1135 ( 
.A(n_1092),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_1073),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1039),
.B(n_1010),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1039),
.B(n_1010),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1071),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1087),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1060),
.Y(n_1141)
);

OAI22x1_ASAP7_75t_L g1142 ( 
.A1(n_1082),
.A2(n_1034),
.B1(n_1036),
.B2(n_886),
.Y(n_1142)
);

BUFx4f_ASAP7_75t_SL g1143 ( 
.A(n_1095),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1042),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1053),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1091),
.B(n_1011),
.Y(n_1146)
);

INVxp67_ASAP7_75t_SL g1147 ( 
.A(n_1056),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1061),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1056),
.A2(n_1020),
.B1(n_1009),
.B2(n_980),
.Y(n_1149)
);

CKINVDCx6p67_ASAP7_75t_R g1150 ( 
.A(n_1083),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1079),
.A2(n_877),
.B1(n_933),
.B2(n_922),
.Y(n_1151)
);

INVx8_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1100),
.A2(n_1030),
.B1(n_980),
.B2(n_972),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1043),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1080),
.A2(n_972),
.B1(n_918),
.B2(n_1022),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1080),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1073),
.A2(n_909),
.B1(n_968),
.B2(n_885),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1070),
.Y(n_1158)
);

INVx6_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

INVxp33_ASAP7_75t_L g1160 ( 
.A(n_1093),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1070),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1042),
.A2(n_1015),
.B(n_930),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_SL g1163 ( 
.A(n_1053),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1135),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1105),
.A2(n_902),
.B(n_883),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_SL g1166 ( 
.A1(n_1136),
.A2(n_1068),
.B1(n_1098),
.B2(n_782),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1111),
.A2(n_1085),
.B1(n_1068),
.B2(n_1022),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1152),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1126),
.A2(n_1085),
.B1(n_1082),
.B2(n_1061),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1126),
.A2(n_1085),
.B1(n_1096),
.B2(n_1088),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1115),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1118),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1111),
.A2(n_866),
.B(n_868),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1114),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1129),
.A2(n_1098),
.B1(n_1009),
.B2(n_1093),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1116),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1120),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1112),
.B(n_1099),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1139),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1147),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1122),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1157),
.A2(n_990),
.B1(n_979),
.B2(n_1007),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1113),
.A2(n_990),
.B1(n_979),
.B2(n_866),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1121),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1113),
.A2(n_1094),
.B1(n_1057),
.B2(n_870),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1117),
.A2(n_870),
.B(n_862),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1134),
.A2(n_1057),
.B1(n_1089),
.B2(n_1044),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1125),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1140),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1110),
.B(n_891),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1134),
.A2(n_1089),
.B1(n_1044),
.B2(n_1015),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1147),
.A2(n_1146),
.B1(n_1132),
.B2(n_1142),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1130),
.A2(n_1131),
.B1(n_1151),
.B2(n_1128),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1160),
.A2(n_907),
.B1(n_911),
.B2(n_878),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1154),
.B(n_891),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1156),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1145),
.B(n_956),
.Y(n_1197)
);

AOI222xp33_ASAP7_75t_L g1198 ( 
.A1(n_1130),
.A2(n_957),
.B1(n_956),
.B2(n_955),
.C1(n_920),
.C2(n_927),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1151),
.B(n_957),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1104),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1131),
.B(n_920),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1133),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1152),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1109),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_SL g1205 ( 
.A(n_1123),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1119),
.B(n_920),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1107),
.A2(n_1124),
.B1(n_1135),
.B2(n_1163),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1149),
.A2(n_1163),
.B1(n_1155),
.B2(n_911),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1153),
.A2(n_916),
.B(n_941),
.Y(n_1209)
);

OAI222xp33_ASAP7_75t_L g1210 ( 
.A1(n_1155),
.A2(n_1153),
.B1(n_1102),
.B2(n_1088),
.C1(n_1086),
.C2(n_1141),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1161),
.A2(n_1044),
.B1(n_1081),
.B2(n_1075),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_L g1212 ( 
.A1(n_1158),
.A2(n_867),
.B(n_864),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1145),
.A2(n_907),
.B1(n_905),
.B2(n_906),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1135),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1162),
.A2(n_873),
.B(n_971),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1145),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1108),
.A2(n_1074),
.B(n_1103),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1143),
.A2(n_1102),
.B1(n_1086),
.B2(n_971),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1143),
.A2(n_1044),
.B1(n_1074),
.B2(n_1050),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1127),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1106),
.A2(n_898),
.B(n_888),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1127),
.A2(n_905),
.B1(n_906),
.B2(n_901),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1144),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1148),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1144),
.A2(n_1081),
.B1(n_1084),
.B2(n_1072),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1159),
.B(n_958),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1159),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1106),
.A2(n_1103),
.B(n_954),
.Y(n_1229)
);

OAI21xp33_ASAP7_75t_L g1230 ( 
.A1(n_1137),
.A2(n_876),
.B(n_867),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1137),
.A2(n_954),
.B(n_952),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1150),
.A2(n_913),
.B1(n_901),
.B2(n_889),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1159),
.A2(n_913),
.B1(n_889),
.B2(n_876),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1152),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1138),
.B(n_958),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1138),
.A2(n_628),
.B1(n_861),
.B2(n_1084),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1170),
.A2(n_628),
.B1(n_610),
.B2(n_861),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1201),
.A2(n_1066),
.B1(n_1072),
.B2(n_1054),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1170),
.A2(n_610),
.B1(n_861),
.B2(n_1026),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1193),
.A2(n_1169),
.B1(n_1186),
.B2(n_1183),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1196),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1202),
.B(n_926),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1173),
.A2(n_1065),
.B1(n_1066),
.B2(n_1063),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1193),
.A2(n_610),
.B1(n_1026),
.B2(n_959),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1169),
.A2(n_610),
.B1(n_1026),
.B2(n_959),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1180),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1185),
.A2(n_959),
.B1(n_1054),
.B2(n_930),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1202),
.A2(n_959),
.B1(n_1054),
.B2(n_931),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1167),
.A2(n_931),
.B1(n_923),
.B2(n_921),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1182),
.A2(n_1065),
.B1(n_1063),
.B2(n_1078),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1178),
.A2(n_865),
.B1(n_927),
.B2(n_926),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1199),
.A2(n_865),
.B1(n_936),
.B2(n_953),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1180),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1192),
.A2(n_865),
.B1(n_936),
.B2(n_953),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1192),
.A2(n_1016),
.B1(n_1006),
.B2(n_952),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1212),
.A2(n_1006),
.B1(n_1016),
.B2(n_984),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1165),
.A2(n_984),
.B1(n_1078),
.B2(n_977),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1187),
.A2(n_996),
.B1(n_1033),
.B2(n_1037),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1232),
.A2(n_996),
.B1(n_942),
.B2(n_1037),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1176),
.A2(n_679),
.B1(n_675),
.B2(n_606),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1197),
.A2(n_679),
.B1(n_675),
.B2(n_606),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1175),
.A2(n_679),
.B1(n_675),
.B2(n_607),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1171),
.B(n_36),
.Y(n_1263)
);

AOI222xp33_ASAP7_75t_L g1264 ( 
.A1(n_1190),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.C1(n_41),
.C2(n_42),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1166),
.A2(n_1198),
.B1(n_1189),
.B2(n_1191),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1230),
.A2(n_679),
.B1(n_675),
.B2(n_606),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1205),
.A2(n_613),
.B1(n_43),
.B2(n_38),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1220),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1208),
.A2(n_607),
.B1(n_594),
.B2(n_613),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1205),
.A2(n_613),
.B1(n_46),
.B2(n_44),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1172),
.A2(n_613),
.B1(n_47),
.B2(n_45),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1229),
.A2(n_1207),
.B1(n_1218),
.B2(n_1179),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1209),
.A2(n_607),
.B1(n_594),
.B2(n_48),
.Y(n_1273)
);

OAI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1231),
.A2(n_1195),
.B1(n_1213),
.B2(n_1233),
.C(n_1194),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1181),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1164),
.A2(n_607),
.B1(n_594),
.B2(n_48),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1235),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1188),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1206),
.A2(n_1219),
.B1(n_1215),
.B2(n_1223),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1219),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1217),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1211),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1174),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1200),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1227),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1224),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1203),
.A2(n_99),
.B(n_97),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1184),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1234),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1228),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1214),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1221),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_1293)
);

AOI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1210),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.C(n_75),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1204),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1222),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1216),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1236),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1168),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1168),
.B(n_100),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1203),
.A2(n_1226),
.B1(n_1225),
.B2(n_105),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1203),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1203),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1276),
.B(n_113),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1297),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1285),
.B(n_119),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1285),
.B(n_122),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1279),
.B(n_123),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1279),
.B(n_124),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1241),
.B(n_127),
.Y(n_1310)
);

OAI221xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1289),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.C(n_133),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1242),
.B(n_134),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1264),
.A2(n_135),
.B(n_136),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1241),
.B(n_137),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1275),
.B(n_139),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1294),
.A2(n_141),
.B(n_142),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1275),
.B(n_144),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1242),
.B(n_145),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1240),
.B(n_148),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1246),
.B(n_149),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1263),
.B(n_387),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1296),
.B(n_150),
.C(n_152),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1246),
.B(n_155),
.Y(n_1323)
);

OAI221xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1265),
.A2(n_1282),
.B1(n_1290),
.B2(n_1291),
.C(n_1270),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1283),
.B(n_156),
.C(n_157),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1255),
.A2(n_158),
.B(n_159),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1253),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_L g1328 ( 
.A(n_1271),
.B(n_162),
.C(n_164),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1274),
.B(n_165),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1281),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1263),
.B(n_386),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1253),
.B(n_172),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1288),
.A2(n_1273),
.B(n_1272),
.Y(n_1333)
);

NOR3xp33_ASAP7_75t_L g1334 ( 
.A(n_1268),
.B(n_174),
.C(n_177),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1238),
.B(n_182),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1254),
.A2(n_183),
.B(n_184),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1267),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1300),
.B(n_190),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1280),
.B(n_191),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1278),
.B(n_194),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1286),
.B(n_196),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1295),
.B(n_197),
.C(n_198),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1292),
.B(n_200),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1257),
.A2(n_203),
.B(n_204),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1293),
.B(n_205),
.Y(n_1345)
);

NOR3xp33_ASAP7_75t_L g1346 ( 
.A(n_1303),
.B(n_206),
.C(n_207),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1287),
.B(n_209),
.C(n_211),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1247),
.B(n_213),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1300),
.B(n_214),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1301),
.B(n_383),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1248),
.B(n_215),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1299),
.B(n_1298),
.C(n_1288),
.Y(n_1352)
);

OAI221xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1277),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.C(n_220),
.Y(n_1353)
);

NAND4xp75_ASAP7_75t_L g1354 ( 
.A(n_1333),
.B(n_1302),
.C(n_1284),
.D(n_1243),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1329),
.B(n_1260),
.C(n_1261),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1327),
.B(n_1318),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1313),
.A2(n_1249),
.B1(n_1250),
.B2(n_1262),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_SL g1358 ( 
.A(n_1334),
.B(n_1284),
.C(n_1245),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_SL g1359 ( 
.A(n_1346),
.B(n_1239),
.C(n_1237),
.Y(n_1359)
);

NAND4xp75_ASAP7_75t_L g1360 ( 
.A(n_1329),
.B(n_1244),
.C(n_1269),
.D(n_224),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1327),
.B(n_1258),
.Y(n_1361)
);

NOR3xp33_ASAP7_75t_L g1362 ( 
.A(n_1311),
.B(n_1259),
.C(n_1251),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1332),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1352),
.A2(n_1252),
.B1(n_1266),
.B2(n_1256),
.Y(n_1364)
);

NAND4xp75_ASAP7_75t_L g1365 ( 
.A(n_1335),
.B(n_221),
.C(n_223),
.D(n_228),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1319),
.B(n_381),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1332),
.B(n_229),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1304),
.B(n_230),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1316),
.B(n_232),
.C(n_234),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1325),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1320),
.B(n_240),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1316),
.B(n_241),
.C(n_243),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1312),
.B(n_244),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1312),
.B(n_1323),
.Y(n_1374)
);

AND2x2_ASAP7_75t_SL g1375 ( 
.A(n_1326),
.B(n_245),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1305),
.B(n_246),
.C(n_248),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1317),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1353),
.B(n_249),
.C(n_252),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_253),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1335),
.A2(n_255),
.B(n_257),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1326),
.B(n_260),
.Y(n_1381)
);

OA211x2_ASAP7_75t_L g1382 ( 
.A1(n_1306),
.A2(n_1307),
.B(n_1308),
.C(n_1309),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1321),
.B(n_261),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1324),
.B(n_263),
.C(n_266),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1315),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1337),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.C(n_275),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1385),
.B(n_1344),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1363),
.B(n_1344),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1356),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1377),
.B(n_1344),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1361),
.B(n_1326),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1375),
.B(n_1336),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1384),
.A2(n_1328),
.B1(n_1322),
.B2(n_1342),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1369),
.B(n_1347),
.C(n_1339),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1381),
.Y(n_1395)
);

XOR2xp5_ASAP7_75t_L g1396 ( 
.A(n_1354),
.B(n_1331),
.Y(n_1396)
);

NAND4xp75_ASAP7_75t_SL g1397 ( 
.A(n_1366),
.B(n_1336),
.C(n_1350),
.D(n_1351),
.Y(n_1397)
);

XNOR2xp5_ASAP7_75t_L g1398 ( 
.A(n_1374),
.B(n_1338),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1372),
.B(n_1310),
.C(n_1314),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1381),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_L g1401 ( 
.A(n_1374),
.B(n_1336),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1367),
.B(n_1338),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1382),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1367),
.B(n_1349),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1379),
.B(n_1340),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1380),
.B(n_1348),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1379),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1380),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1400),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1395),
.Y(n_1410)
);

XOR2xp5_ASAP7_75t_L g1411 ( 
.A(n_1396),
.B(n_1355),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1395),
.Y(n_1412)
);

XOR2x2_ASAP7_75t_L g1413 ( 
.A(n_1398),
.B(n_1378),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1390),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1403),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1389),
.Y(n_1416)
);

XOR2x2_ASAP7_75t_L g1417 ( 
.A(n_1398),
.B(n_1365),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1407),
.Y(n_1418)
);

XNOR2xp5_ASAP7_75t_L g1419 ( 
.A(n_1397),
.B(n_1383),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1403),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1392),
.A2(n_1373),
.B1(n_1341),
.B2(n_1343),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1409),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1420),
.Y(n_1423)
);

AOI22x1_ASAP7_75t_L g1424 ( 
.A1(n_1411),
.A2(n_1392),
.B1(n_1406),
.B2(n_1408),
.Y(n_1424)
);

AOI22x1_ASAP7_75t_L g1425 ( 
.A1(n_1421),
.A2(n_1406),
.B1(n_1408),
.B2(n_1387),
.Y(n_1425)
);

AOI22x1_ASAP7_75t_L g1426 ( 
.A1(n_1419),
.A2(n_1387),
.B1(n_1405),
.B2(n_1391),
.Y(n_1426)
);

OAI22x1_ASAP7_75t_L g1427 ( 
.A1(n_1415),
.A2(n_1401),
.B1(n_1393),
.B2(n_1391),
.Y(n_1427)
);

OA22x2_ASAP7_75t_L g1428 ( 
.A1(n_1415),
.A2(n_1416),
.B1(n_1413),
.B2(n_1417),
.Y(n_1428)
);

AO22x2_ASAP7_75t_L g1429 ( 
.A1(n_1410),
.A2(n_1405),
.B1(n_1394),
.B2(n_1399),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1410),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1418),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1412),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1412),
.B(n_1388),
.Y(n_1433)
);

OA22x2_ASAP7_75t_SL g1434 ( 
.A1(n_1413),
.A2(n_1358),
.B1(n_1330),
.B2(n_1388),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_1414),
.Y(n_1435)
);

AOI22x1_ASAP7_75t_L g1436 ( 
.A1(n_1414),
.A2(n_1390),
.B1(n_1368),
.B2(n_1371),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1423),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1422),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1431),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1430),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1428),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1429),
.Y(n_1442)
);

INVx8_ASAP7_75t_L g1443 ( 
.A(n_1434),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1427),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1441),
.A2(n_1428),
.B1(n_1429),
.B2(n_1434),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1438),
.Y(n_1446)
);

AOI22x1_ASAP7_75t_L g1447 ( 
.A1(n_1442),
.A2(n_1429),
.B1(n_1432),
.B2(n_1424),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1443),
.A2(n_1426),
.B1(n_1425),
.B2(n_1436),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1441),
.A2(n_1443),
.B1(n_1444),
.B2(n_1437),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1439),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1446),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1450),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1449),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1445),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1448),
.A2(n_1443),
.B1(n_1440),
.B2(n_1435),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1447),
.A2(n_1435),
.B1(n_1433),
.B2(n_1402),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1454),
.A2(n_1433),
.B1(n_1362),
.B2(n_1386),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1453),
.A2(n_1376),
.B1(n_1360),
.B2(n_1359),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1451),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1452),
.B(n_1404),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1455),
.B(n_1456),
.C(n_1386),
.D(n_1357),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1454),
.A2(n_1370),
.B1(n_1364),
.B2(n_1345),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1451),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1454),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1461),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1457),
.A2(n_1458),
.B1(n_1462),
.B2(n_1464),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1460),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1459),
.A2(n_290),
.B1(n_295),
.B2(n_298),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1463),
.B(n_301),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1460),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1460),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1469),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1470),
.Y(n_1473)
);

AO22x2_ASAP7_75t_L g1474 ( 
.A1(n_1471),
.A2(n_303),
.B1(n_305),
.B2(n_310),
.Y(n_1474)
);

NOR4xp25_ASAP7_75t_L g1475 ( 
.A(n_1466),
.B(n_312),
.C(n_313),
.D(n_315),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1465),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1467),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1476),
.A2(n_1468),
.B1(n_319),
.B2(n_320),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1473),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1474),
.Y(n_1480)
);

INVxp33_ASAP7_75t_SL g1481 ( 
.A(n_1475),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1472),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1474),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1477),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1480),
.Y(n_1485)
);

OAI22x1_ASAP7_75t_L g1486 ( 
.A1(n_1483),
.A2(n_317),
.B1(n_324),
.B2(n_325),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1484),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1481),
.A2(n_326),
.B1(n_329),
.B2(n_330),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1479),
.Y(n_1489)
);

OAI211xp5_ASAP7_75t_L g1490 ( 
.A1(n_1482),
.A2(n_1478),
.B(n_335),
.C(n_338),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1485),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1487),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1489),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1486),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1488),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1491),
.A2(n_1478),
.B1(n_1490),
.B2(n_342),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1495),
.A2(n_332),
.B1(n_339),
.B2(n_345),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1494),
.A2(n_351),
.B1(n_352),
.B2(n_354),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1496),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1497),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1500),
.A2(n_1493),
.B1(n_1492),
.B2(n_1498),
.Y(n_1501)
);

AO22x2_ASAP7_75t_L g1502 ( 
.A1(n_1499),
.A2(n_355),
.B1(n_360),
.B2(n_362),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1501),
.Y(n_1503)
);

AO22x2_ASAP7_75t_L g1504 ( 
.A1(n_1503),
.A2(n_1502),
.B1(n_367),
.B2(n_371),
.Y(n_1504)
);

AOI211xp5_ASAP7_75t_L g1505 ( 
.A1(n_1504),
.A2(n_364),
.B(n_372),
.C(n_373),
.Y(n_1505)
);


endmodule