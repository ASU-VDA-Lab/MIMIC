module fake_jpeg_1390_n_688 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_688);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_688;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_70),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_71),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_83),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_80),
.Y(n_223)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_32),
.Y(n_82)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_82),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_18),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_84),
.B(n_94),
.Y(n_180)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_86),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_102),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_108),
.B(n_112),
.Y(n_213)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_31),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_114),
.B(n_35),
.Y(n_211)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_117),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx2_ASAP7_75t_R g120 ( 
.A(n_48),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_40),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_20),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_22),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_20),
.Y(n_128)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g129 ( 
.A(n_22),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g215 ( 
.A(n_129),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_20),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_22),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_25),
.Y(n_152)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_25),
.Y(n_132)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_59),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_149),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_152),
.B(n_170),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_25),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_153),
.B(n_156),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_57),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_158),
.B(n_178),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_71),
.A2(n_26),
.B(n_58),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_159),
.B(n_161),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_79),
.B(n_57),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_164),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_74),
.B(n_17),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_167),
.B(n_168),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_71),
.A2(n_26),
.B(n_58),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_57),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_111),
.B(n_17),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_82),
.B(n_39),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_181),
.B(n_182),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_39),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_38),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_185),
.B(n_192),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_61),
.A2(n_38),
.B1(n_35),
.B2(n_59),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_187),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_251)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_190),
.Y(n_286)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_38),
.Y(n_192)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_88),
.B(n_35),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_203),
.B(n_211),
.Y(n_297)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_88),
.B(n_21),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_219),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_110),
.A2(n_21),
.B1(n_58),
.B2(n_50),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_214),
.A2(n_49),
.B1(n_44),
.B2(n_36),
.Y(n_274)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_93),
.B(n_59),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_222),
.Y(n_262)
);

BUFx16f_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_229),
.Y(n_365)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_231),
.Y(n_318)
);

CKINVDCx9p33_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_232),
.Y(n_352)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_152),
.A2(n_123),
.B1(n_36),
.B2(n_37),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_237),
.A2(n_241),
.B1(n_246),
.B2(n_254),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_144),
.B(n_30),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_238),
.B(n_240),
.Y(n_324)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_239),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_144),
.B(n_30),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_170),
.A2(n_105),
.B1(n_103),
.B2(n_102),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_137),
.A2(n_72),
.B(n_27),
.C(n_50),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_242),
.A2(n_292),
.B(n_5),
.Y(n_319)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_244),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_245),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_153),
.A2(n_24),
.B1(n_21),
.B2(n_27),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_248),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_249),
.B(n_252),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_251),
.A2(n_218),
.B1(n_174),
.B2(n_136),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_147),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_137),
.B(n_27),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_259),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_181),
.A2(n_24),
.B1(n_30),
.B2(n_36),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_255),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_185),
.A2(n_95),
.B1(n_97),
.B2(n_24),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_256),
.A2(n_295),
.B1(n_299),
.B2(n_214),
.Y(n_308)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_147),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_135),
.Y(n_260)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_221),
.B(n_45),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_261),
.B(n_175),
.C(n_176),
.Y(n_354)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_192),
.A2(n_45),
.B1(n_37),
.B2(n_43),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_265),
.B(n_142),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_138),
.B(n_49),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

CKINVDCx12_ASAP7_75t_R g271 ( 
.A(n_215),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_271),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g272 ( 
.A1(n_189),
.A2(n_49),
.B1(n_43),
.B2(n_44),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_149),
.B(n_50),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_274),
.A2(n_175),
.B1(n_140),
.B2(n_203),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_158),
.B(n_44),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_275),
.B(n_278),
.Y(n_344)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_101),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_151),
.Y(n_279)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_282),
.B(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_226),
.B(n_92),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_96),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_291),
.Y(n_368)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_161),
.B(n_0),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_210),
.B(n_2),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_202),
.Y(n_298)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_183),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_163),
.Y(n_303)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_173),
.Y(n_304)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_177),
.Y(n_306)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_166),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_169),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_308),
.A2(n_321),
.B1(n_335),
.B2(n_243),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_313),
.B(n_354),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_319),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_280),
.A2(n_165),
.B1(n_157),
.B2(n_188),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_247),
.B(n_186),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_331),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_236),
.A2(n_174),
.B1(n_172),
.B2(n_171),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_327),
.A2(n_307),
.B1(n_303),
.B2(n_281),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_269),
.Y(n_331)
);

FAx1_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_205),
.CI(n_197),
.CON(n_334),
.SN(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_334),
.A2(n_261),
.B(n_295),
.C(n_274),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_237),
.A2(n_220),
.B1(n_224),
.B2(n_194),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_236),
.B(n_297),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_360),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_272),
.A2(n_140),
.B1(n_177),
.B2(n_225),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_351),
.B1(n_353),
.B2(n_359),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_272),
.A2(n_225),
.B1(n_193),
.B2(n_199),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_272),
.A2(n_193),
.B1(n_199),
.B2(n_209),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_357),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_292),
.B(n_179),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_305),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_258),
.B(n_154),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_227),
.A2(n_207),
.B1(n_198),
.B2(n_146),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_254),
.B1(n_246),
.B2(n_265),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_261),
.B(n_242),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_343),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_324),
.B(n_250),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_370),
.B(n_374),
.Y(n_423)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_230),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_375),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_232),
.Y(n_377)
);

OAI31xp33_ASAP7_75t_L g455 ( 
.A1(n_377),
.A2(n_399),
.A3(n_401),
.B(n_416),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_334),
.A2(n_255),
.B1(n_243),
.B2(n_293),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_379),
.A2(n_398),
.B1(n_407),
.B2(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_228),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_382),
.B(n_384),
.Y(n_424)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_228),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_390),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_388),
.A2(n_391),
.B1(n_329),
.B2(n_337),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_316),
.A2(n_286),
.B1(n_281),
.B2(n_267),
.Y(n_391)
);

INVx13_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_355),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_413),
.Y(n_448)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_403),
.Y(n_453)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

INVx13_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_205),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_299),
.B(n_274),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_336),
.Y(n_402)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_368),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_404),
.B(n_417),
.Y(n_440)
);

OAI22x1_ASAP7_75t_SL g405 ( 
.A1(n_313),
.A2(n_279),
.B1(n_260),
.B2(n_262),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_418),
.B1(n_359),
.B2(n_357),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_414),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_309),
.A2(n_356),
.B1(n_352),
.B2(n_354),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_323),
.B(n_264),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_411),
.Y(n_428)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_264),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_364),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_355),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_317),
.B(n_339),
.C(n_338),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_415),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_309),
.A2(n_262),
.B1(n_304),
.B2(n_266),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_330),
.B(n_266),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_309),
.A2(n_136),
.B1(n_218),
.B2(n_306),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_420),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_327),
.B1(n_358),
.B2(n_364),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_422),
.A2(n_433),
.B1(n_439),
.B2(n_373),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_358),
.B(n_345),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_429),
.A2(n_436),
.B(n_371),
.Y(n_473)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_432),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_376),
.A2(n_320),
.B1(n_332),
.B2(n_341),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_376),
.A2(n_400),
.B(n_377),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_410),
.B(n_399),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_376),
.A2(n_400),
.B(n_406),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_378),
.B(n_310),
.C(n_312),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_437),
.B(n_362),
.C(n_285),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_389),
.A2(n_332),
.B1(n_320),
.B2(n_315),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_387),
.A2(n_244),
.B1(n_257),
.B2(n_263),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_447),
.A2(n_458),
.B1(n_459),
.B2(n_396),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_378),
.B(n_347),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_450),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_347),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_414),
.B(n_342),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_452),
.B(n_340),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_375),
.Y(n_454)
);

INVx13_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_386),
.A2(n_314),
.B1(n_245),
.B2(n_294),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_408),
.A2(n_302),
.B1(n_367),
.B2(n_322),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_435),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_483),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_417),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_458),
.A2(n_418),
.B1(n_388),
.B2(n_400),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_462),
.A2(n_464),
.B(n_469),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_411),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_482),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_419),
.A2(n_405),
.B(n_416),
.C(n_403),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_467),
.A2(n_473),
.B(n_489),
.Y(n_508)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_434),
.A2(n_413),
.B(n_393),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_470),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_403),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_480),
.C(n_481),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_422),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_419),
.A2(n_372),
.B1(n_380),
.B2(n_402),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_474),
.A2(n_491),
.B1(n_427),
.B2(n_430),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_395),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_477),
.B(n_444),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_424),
.Y(n_478)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_478),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_421),
.B(n_348),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_348),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_423),
.B(n_337),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_398),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_333),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_486),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_432),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_453),
.Y(n_514)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_488),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_429),
.A2(n_397),
.B(n_340),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_419),
.A2(n_385),
.B1(n_394),
.B2(n_412),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_448),
.B(n_383),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_493),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_449),
.B(n_362),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_453),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_385),
.Y(n_495)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_495),
.Y(n_513)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_496),
.Y(n_510)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_526),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_428),
.C(n_433),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_522),
.C(n_494),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_503),
.B(n_528),
.Y(n_551)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_514),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_479),
.Y(n_515)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_515),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_451),
.B(n_455),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_516),
.Y(n_540)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_465),
.A2(n_420),
.B1(n_439),
.B2(n_453),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_519),
.A2(n_463),
.B1(n_481),
.B2(n_466),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_438),
.Y(n_520)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_438),
.C(n_427),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_469),
.A2(n_459),
.B(n_430),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_SL g552 ( 
.A1(n_524),
.A2(n_467),
.B(n_475),
.C(n_445),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_525),
.A2(n_468),
.B1(n_497),
.B2(n_485),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_474),
.A2(n_472),
.B1(n_491),
.B2(n_487),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_489),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_529),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_464),
.A2(n_444),
.B(n_446),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_446),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_530),
.B(n_532),
.Y(n_562)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_490),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_447),
.Y(n_533)
);

INVxp33_ASAP7_75t_SL g539 ( 
.A(n_533),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_505),
.B(n_478),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_535),
.B(n_537),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_536),
.A2(n_524),
.B1(n_520),
.B2(n_506),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_531),
.B(n_492),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_553),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_463),
.C(n_495),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_541),
.B(n_550),
.C(n_556),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_498),
.B(n_483),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_544),
.B(n_546),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_443),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_545),
.B(n_554),
.Y(n_580)
);

XNOR2x1_ASAP7_75t_L g546 ( 
.A(n_503),
.B(n_475),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_547),
.A2(n_543),
.B1(n_539),
.B2(n_525),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_499),
.A2(n_485),
.B1(n_467),
.B2(n_475),
.Y(n_549)
);

INVxp33_ASAP7_75t_SL g579 ( 
.A(n_549),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_502),
.B(n_528),
.C(n_533),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_524),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_467),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_504),
.B(n_443),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_467),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_555),
.B(n_560),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_445),
.C(n_318),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_507),
.B(n_457),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_558),
.B(n_559),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_SL g559 ( 
.A(n_509),
.B(n_496),
.C(n_457),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_501),
.B(n_441),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_521),
.B(n_333),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_561),
.B(n_365),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_441),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_513),
.C(n_530),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_510),
.B(n_442),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_564),
.B(n_515),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_540),
.A2(n_509),
.B(n_508),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_569),
.A2(n_574),
.B(n_365),
.Y(n_614)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_562),
.Y(n_571)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_571),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_536),
.A2(n_499),
.B1(n_526),
.B2(n_513),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_573),
.A2(n_589),
.B1(n_594),
.B2(n_392),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_540),
.A2(n_508),
.B(n_534),
.Y(n_574)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_566),
.Y(n_576)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_576),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_SL g603 ( 
.A1(n_577),
.A2(n_559),
.B(n_546),
.C(n_550),
.Y(n_603)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_565),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_578),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_581),
.B(n_496),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_582),
.B(n_556),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_500),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_583),
.B(n_588),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_539),
.A2(n_519),
.B1(n_532),
.B2(n_523),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_584),
.A2(n_592),
.B1(n_593),
.B2(n_552),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_587),
.A2(n_552),
.B1(n_555),
.B2(n_553),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_548),
.A2(n_514),
.B1(n_506),
.B2(n_534),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_590),
.B(n_318),
.Y(n_609)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_567),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_511),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_542),
.A2(n_557),
.B1(n_560),
.B2(n_563),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_542),
.A2(n_518),
.B1(n_517),
.B2(n_512),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_552),
.A2(n_517),
.B1(n_512),
.B2(n_511),
.Y(n_594)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_596),
.A2(n_599),
.B1(n_617),
.B2(n_594),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_597),
.B(n_603),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_585),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_598),
.B(n_607),
.C(n_611),
.Y(n_630)
);

BUFx12_ASAP7_75t_L g600 ( 
.A(n_579),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_600),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_538),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_601),
.B(n_612),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_SL g606 ( 
.A(n_570),
.B(n_544),
.C(n_551),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_606),
.B(n_610),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_568),
.B(n_551),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_609),
.A2(n_591),
.B1(n_578),
.B2(n_586),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_575),
.B(n_442),
.C(n_361),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_571),
.B(n_570),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_569),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_613),
.B(n_616),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_614),
.A2(n_197),
.B(n_293),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_615),
.A2(n_593),
.B1(n_577),
.B2(n_576),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_581),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_587),
.A2(n_267),
.B1(n_285),
.B2(n_381),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_605),
.Y(n_618)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_618),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_620),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_621),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_572),
.C(n_592),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_623),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_572),
.C(n_586),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_574),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_624),
.B(n_628),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_625),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_288),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_599),
.B(n_288),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_617),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_615),
.A2(n_288),
.B(n_239),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_632),
.A2(n_602),
.B(n_608),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_603),
.A2(n_231),
.B(n_277),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_635),
.B(n_603),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_604),
.B(n_231),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_636),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_637),
.B(n_602),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_638),
.A2(n_648),
.B1(n_650),
.B2(n_653),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_642),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_619),
.B(n_600),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_643),
.B(n_647),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_626),
.B(n_600),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_620),
.Y(n_648)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_634),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_633),
.B(n_603),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_652),
.B(n_624),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_640),
.A2(n_627),
.B(n_630),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_654),
.A2(n_659),
.B(n_665),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_651),
.B(n_644),
.C(n_643),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_663),
.Y(n_669)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_658),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_631),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_646),
.A2(n_622),
.B(n_619),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_661),
.A2(n_662),
.B(n_664),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_623),
.C(n_637),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_649),
.B(n_628),
.C(n_636),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_645),
.B(n_629),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_638),
.A2(n_632),
.B(n_229),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_655),
.A2(n_639),
.B1(n_642),
.B2(n_133),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_667),
.A2(n_674),
.B(n_10),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_SL g670 ( 
.A1(n_659),
.A2(n_197),
.B(n_229),
.C(n_164),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g678 ( 
.A(n_670),
.B(n_13),
.Y(n_678)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_660),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_671),
.B(n_672),
.Y(n_679)
);

AOI322xp5_ASAP7_75t_L g672 ( 
.A1(n_664),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_656),
.B(n_6),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_666),
.A2(n_6),
.B(n_9),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_675),
.A2(n_676),
.B(n_678),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_669),
.B(n_10),
.C(n_13),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_677),
.Y(n_680)
);

A2O1A1O1Ixp25_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_668),
.B(n_673),
.C(n_667),
.D(n_15),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_682),
.A2(n_13),
.B(n_14),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_683),
.B(n_684),
.C(n_681),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_680),
.B(n_14),
.Y(n_684)
);

BUFx24_ASAP7_75t_SL g686 ( 
.A(n_685),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_14),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_14),
.B(n_15),
.Y(n_688)
);


endmodule