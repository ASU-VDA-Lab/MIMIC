module fake_jpeg_27140_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_28),
.Y(n_38)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_7),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_7),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.CON(n_36),
.SN(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_7),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_20),
.B1(n_13),
.B2(n_18),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_20),
.B1(n_13),
.B2(n_19),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_31),
.B(n_15),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_14),
.B1(n_39),
.B2(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_29),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_53),
.Y(n_62)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_31),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_43),
.B1(n_53),
.B2(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_12),
.B(n_21),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_24),
.C(n_8),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_14),
.B1(n_22),
.B2(n_21),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_69),
.B1(n_58),
.B2(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_25),
.B1(n_26),
.B2(n_12),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_26),
.B1(n_12),
.B2(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_78),
.B1(n_61),
.B2(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_16),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_51),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_86),
.A2(n_21),
.B(n_22),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_19),
.B(n_11),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_11),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_81),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_68),
.A3(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_63),
.B1(n_69),
.B2(n_61),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_71),
.B1(n_56),
.B2(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_78),
.B1(n_75),
.B2(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_86),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_34),
.B(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_114),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_41),
.C(n_56),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_111),
.C(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_41),
.C(n_46),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_44),
.B1(n_41),
.B2(n_30),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_44),
.B1(n_96),
.B2(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_41),
.C(n_34),
.Y(n_117)
);

AOI21x1_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_116),
.B(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_27),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_89),
.C(n_93),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_129),
.C(n_131),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_89),
.B(n_9),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.C(n_106),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_51),
.C(n_30),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_30),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_51),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_102),
.B1(n_117),
.B2(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_139),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_30),
.C(n_27),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_122),
.C(n_131),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_124),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_130),
.C(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_143),
.B(n_118),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_161),
.B(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_162),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_143),
.B(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_135),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_121),
.B1(n_144),
.B2(n_27),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_5),
.B(n_10),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_147),
.C(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_146),
.C(n_27),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_157),
.B(n_4),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_177),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_1),
.C(n_2),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_167),
.CI(n_9),
.CON(n_181),
.SN(n_181)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_181),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_1),
.A3(n_2),
.B1(n_176),
.B2(n_179),
.C1(n_181),
.C2(n_180),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_1),
.B(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);


endmodule