module fake_jpeg_28798_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_62),
.B1(n_49),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_93),
.B1(n_66),
.B2(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_65),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_54),
.Y(n_97)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_69),
.B1(n_54),
.B2(n_62),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_77),
.B(n_61),
.C(n_68),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_21),
.B1(n_45),
.B2(n_44),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_59),
.B1(n_53),
.B2(n_69),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_24),
.B(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_107),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_54),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_111),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_60),
.B(n_53),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_83),
.C(n_80),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_67),
.B1(n_63),
.B2(n_55),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_23),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_126),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_127),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_26),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_77),
.B1(n_88),
.B2(n_2),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_18),
.B(n_40),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_15),
.C(n_38),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_131),
.B1(n_33),
.B2(n_46),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_27),
.B1(n_37),
.B2(n_36),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_22),
.B(n_25),
.C(n_29),
.D(n_30),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_148),
.C(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_112),
.Y(n_156)
);

NOR4xp25_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_129),
.C(n_115),
.D(n_122),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_141),
.B1(n_146),
.B2(n_135),
.C(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_143),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_157),
.C(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.C(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_153),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_150),
.B(n_149),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_150),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_112),
.B(n_133),
.Y(n_169)
);


endmodule