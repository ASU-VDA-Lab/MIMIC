module real_jpeg_14507_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_249, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_249;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_3),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_4),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_6),
.A2(n_30),
.B1(n_38),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_7),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_109),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_109),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_30),
.B1(n_38),
.B2(n_109),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_10),
.A2(n_44),
.B1(n_60),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_30),
.B1(n_38),
.B2(n_44),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_12),
.A2(n_60),
.B1(n_63),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_79),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_30),
.B1(n_38),
.B2(n_79),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_112),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_65),
.B(n_165),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_100),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_46),
.B(n_50),
.C(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_13),
.B(n_105),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_34),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_86),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_13),
.A2(n_63),
.B(n_73),
.C(n_220),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_30),
.B1(n_38),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_68),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_15),
.A2(n_30),
.B1(n_38),
.B2(n_68),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_16),
.A2(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_16),
.A2(n_30),
.B1(n_38),
.B2(n_70),
.Y(n_193)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_133),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_131),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_113),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_22),
.B(n_113),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.C(n_92),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_23),
.A2(n_24),
.B1(n_81),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_55),
.B2(n_56),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_57),
.C(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_27),
.B(n_41),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_28),
.A2(n_33),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_29),
.A2(n_34),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_29),
.A2(n_34),
.B(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_29),
.A2(n_34),
.B1(n_96),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_29),
.A2(n_34),
.B1(n_147),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_29),
.A2(n_34),
.B1(n_159),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_29),
.A2(n_34),
.B1(n_100),
.B2(n_205),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_29),
.A2(n_34),
.B1(n_198),
.B2(n_205),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_38),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_30),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_38),
.A2(n_51),
.B(n_100),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_43),
.A2(n_48),
.B1(n_86),
.B2(n_151),
.Y(n_168)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_46),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_45),
.A2(n_63),
.A3(n_75),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_46),
.B(n_76),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_47),
.A2(n_52),
.B1(n_150),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_48),
.A2(n_85),
.B1(n_86),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_86),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_48),
.A2(n_86),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_48),
.A2(n_86),
.B1(n_184),
.B2(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_69),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_58),
.A2(n_59),
.B1(n_108),
.B2(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_60),
.B(n_100),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_63),
.Y(n_98)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_66),
.B(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_77),
.B1(n_80),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_72),
.A2(n_77),
.B1(n_103),
.B2(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_73),
.A2(n_105),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_77),
.A2(n_141),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_81),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_91),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_92),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.C(n_106),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_93),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_101),
.B(n_106),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_233),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_176),
.B(n_232),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_160),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_137),
.B(n_160),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_152),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_138),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_145),
.C(n_146),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_175),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_172),
.C(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_226),
.B(n_231),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_225),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_194),
.B(n_213),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_202),
.B(n_212),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_200),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_221),
.C(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);


endmodule