module fake_netlist_6_4757_n_1983 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1983);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1983;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_138),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_115),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_37),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_41),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_1),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_131),
.Y(n_219)
);

BUFx2_ASAP7_75t_SL g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_39),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_30),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_15),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_127),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_75),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_61),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_47),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_55),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_67),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_91),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_40),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_155),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_24),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_2),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_64),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_85),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_177),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_124),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_42),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_139),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_126),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_27),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_82),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_160),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_68),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_129),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_189),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_14),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_151),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_33),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_89),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_105),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_5),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_128),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_50),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_143),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_132),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_121),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_136),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_174),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_125),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_17),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_93),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_7),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_39),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_101),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_122),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_43),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_188),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_137),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_63),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_20),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_32),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_166),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_112),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_25),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_84),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_142),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_48),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_60),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_167),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_141),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_49),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_32),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_186),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_67),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_66),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_157),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_62),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_185),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_16),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_3),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_37),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_64),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_99),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_13),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_7),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_27),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_9),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_123),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_49),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_100),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_180),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_8),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_52),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_103),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_178),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_110),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_62),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_175),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_149),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_1),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_69),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_10),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_42),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_164),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_55),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_24),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_53),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_45),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_60),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_61),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_8),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_107),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_28),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_0),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_76),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_15),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_33),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_41),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_104),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_90),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_74),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_48),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_54),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_87),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_11),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_117),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_36),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_81),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_102),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_88),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_159),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_86),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_119),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_19),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_96),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_36),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_65),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_109),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_79),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_52),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_281),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_281),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_195),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_199),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_202),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_241),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_281),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_211),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_217),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_281),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_219),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_226),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_227),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_281),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_204),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_281),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_251),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_376),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_272),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_228),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_272),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_316),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_254),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_213),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_235),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_388),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_238),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_239),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_252),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_307),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_267),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_288),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_241),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_340),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_244),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_210),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_210),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_293),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_203),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_218),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_317),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_192),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_245),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_254),
.B(n_0),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_218),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_225),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_225),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_229),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_229),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_232),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_232),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_233),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_377),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_386),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_248),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_233),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_249),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_237),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_250),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_237),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_256),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_192),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_240),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_260),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_193),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_261),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_263),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_340),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_240),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_342),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_277),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_264),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_269),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_271),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_277),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_378),
.B(n_2),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_257),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_257),
.B(n_3),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_273),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_378),
.B(n_6),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_283),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_316),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_283),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_286),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_274),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_286),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_292),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_205),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_292),
.B(n_6),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_300),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_205),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_278),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_282),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_207),
.B(n_11),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_300),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_302),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_284),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_433),
.B(n_203),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_391),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_203),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_398),
.B(n_287),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g499 ( 
.A(n_436),
.B(n_203),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_401),
.B(n_436),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_325),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_325),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_422),
.A2(n_268),
.B1(n_266),
.B2(n_242),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_456),
.B(n_203),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_396),
.B(n_253),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_406),
.B(n_408),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_424),
.A2(n_382),
.B1(n_375),
.B2(n_346),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_401),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_404),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_427),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_297),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_200),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_414),
.B(n_302),
.Y(n_532)
);

OA21x2_ASAP7_75t_L g533 ( 
.A1(n_417),
.A2(n_315),
.B(n_303),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_414),
.B(n_299),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_220),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_418),
.Y(n_537)
);

CKINVDCx8_ASAP7_75t_R g538 ( 
.A(n_428),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_441),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_442),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_442),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_438),
.B(n_200),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_488),
.B(n_309),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_472),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_444),
.B(n_314),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_392),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_445),
.B(n_321),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_415),
.B(n_387),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_465),
.B(n_387),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_445),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_450),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_407),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_454),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_409),
.B(n_303),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_457),
.B(n_323),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_463),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_463),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_475),
.A2(n_333),
.B(n_276),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_393),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_276),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_505),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_394),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_544),
.B(n_545),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_567),
.Y(n_580)
);

INVx8_ASAP7_75t_L g581 ( 
.A(n_536),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_544),
.A2(n_469),
.B1(n_470),
.B2(n_410),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_554),
.A2(n_483),
.B1(n_315),
.B2(n_327),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_548),
.B(n_504),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_530),
.B(n_409),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_561),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_420),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_548),
.B(n_397),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_500),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_503),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_530),
.B(n_420),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_551),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_545),
.B(n_459),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_491),
.B(n_395),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_530),
.B(n_399),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_506),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_567),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_505),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_491),
.B(n_400),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_554),
.A2(n_555),
.B1(n_497),
.B2(n_536),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_498),
.B(n_402),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_553),
.B(n_403),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_533),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_553),
.B(n_405),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_553),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_524),
.B(n_428),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_492),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_498),
.B(n_521),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_524),
.B(n_462),
.Y(n_619)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_510),
.A2(n_483),
.B(n_212),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_533),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_524),
.B(n_412),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_533),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_SL g626 ( 
.A(n_564),
.B(n_458),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_524),
.B(n_419),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_555),
.B(n_333),
.Y(n_629)
);

CKINVDCx14_ASAP7_75t_R g630 ( 
.A(n_520),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_494),
.Y(n_631)
);

NOR2x1p5_ASAP7_75t_L g632 ( 
.A(n_524),
.B(n_397),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_521),
.B(n_421),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_504),
.B(n_477),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_495),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_527),
.Y(n_636)
);

AND3x1_ASAP7_75t_L g637 ( 
.A(n_506),
.B(n_327),
.C(n_322),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_527),
.Y(n_638)
);

BUFx4f_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_341),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_527),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_564),
.B(n_220),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_502),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_504),
.B(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_503),
.B(n_478),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_509),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_509),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_511),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_503),
.B(n_341),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_511),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_561),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_534),
.B(n_429),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_538),
.B(n_462),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_523),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_505),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_497),
.A2(n_322),
.B1(n_338),
.B2(n_339),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_536),
.A2(n_338),
.B1(n_339),
.B2(n_351),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_538),
.B(n_464),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_512),
.A2(n_352),
.B1(n_347),
.B2(n_294),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_505),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_493),
.B(n_207),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_538),
.B(n_464),
.Y(n_666)
);

INVx8_ASAP7_75t_L g667 ( 
.A(n_536),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_522),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_523),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_550),
.B(n_437),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_523),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_536),
.B(n_212),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_550),
.B(n_449),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_505),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_536),
.B(n_570),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_L g679 ( 
.A(n_493),
.B(n_216),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_532),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_552),
.B(n_451),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_532),
.B(n_430),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_570),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_532),
.B(n_431),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_519),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_552),
.B(n_453),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_508),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_565),
.B(n_455),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_493),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_505),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_493),
.B(n_216),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_563),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_565),
.B(n_466),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_493),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_516),
.B(n_467),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_563),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_519),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_501),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_568),
.A2(n_351),
.B1(n_356),
.B2(n_363),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_516),
.B(n_468),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_526),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_512),
.B(n_473),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_568),
.B(n_479),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_501),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_568),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_501),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_501),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_570),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_518),
.B(n_487),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_526),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_518),
.B(n_224),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_516),
.B(n_460),
.Y(n_721)
);

NOR2x2_ASAP7_75t_L g722 ( 
.A(n_643),
.B(n_508),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_618),
.B(n_516),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_579),
.B(n_516),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_716),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_591),
.B(n_416),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_591),
.B(n_423),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_543),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_716),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_680),
.B(n_675),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_581),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_706),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_595),
.B(n_608),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_617),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_673),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_678),
.B(n_461),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_673),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_617),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_601),
.A2(n_363),
.B(n_369),
.C(n_356),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_641),
.B(n_543),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_573),
.B(n_493),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_543),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_634),
.B(n_528),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_606),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_578),
.B(n_543),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_597),
.B(n_546),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_678),
.B(n_486),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_657),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_604),
.B(n_425),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_610),
.B(n_546),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_633),
.B(n_546),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_706),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_589),
.B(n_426),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_671),
.B(n_546),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_706),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_648),
.B(n_528),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_606),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_589),
.B(n_648),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_678),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_687),
.B(n_691),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_661),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_598),
.B(n_432),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_684),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_698),
.B(n_558),
.Y(n_768)
);

NAND2x1_ASAP7_75t_L g769 ( 
.A(n_699),
.B(n_493),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_718),
.B(n_558),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_621),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_669),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_655),
.B(n_558),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_634),
.B(n_646),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_624),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_585),
.B(n_435),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_681),
.B(n_560),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_639),
.B(n_313),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_624),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_654),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_639),
.B(n_328),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_669),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_672),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_672),
.Y(n_784)
);

AND2x6_ASAP7_75t_SL g785 ( 
.A(n_643),
.B(n_369),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_580),
.B(n_584),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_580),
.B(n_560),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_584),
.B(n_596),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_639),
.B(n_335),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_596),
.B(n_560),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_600),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_585),
.B(n_447),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_674),
.B(n_682),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_684),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_601),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_560),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_631),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_573),
.A2(n_448),
.B1(n_336),
.B2(n_345),
.Y(n_798)
);

NOR2x1p5_ASAP7_75t_L g799 ( 
.A(n_588),
.B(n_196),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_573),
.A2(n_368),
.B1(n_236),
.B2(n_243),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_581),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_631),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_573),
.A2(n_374),
.B1(n_350),
.B2(n_359),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_683),
.B(n_508),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_627),
.B(n_562),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_699),
.B(n_224),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_682),
.A2(n_291),
.B1(n_236),
.B2(n_383),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_683),
.B(n_247),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_627),
.B(n_562),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_635),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_612),
.B(n_329),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_636),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_646),
.B(n_535),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_609),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_614),
.B(n_355),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_636),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_615),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_638),
.Y(n_820)
);

O2A1O1Ixp5_ASAP7_75t_L g821 ( 
.A1(n_717),
.A2(n_291),
.B(n_243),
.C(n_246),
.Y(n_821)
);

OAI22x1_ASAP7_75t_R g822 ( 
.A1(n_599),
.A2(n_295),
.B1(n_279),
.B2(n_275),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_599),
.B(n_446),
.C(n_439),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_644),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_674),
.B(n_362),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_642),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_674),
.B(n_366),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_644),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_583),
.A2(n_704),
.B1(n_660),
.B2(n_582),
.C(n_659),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_642),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_615),
.B(n_198),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_573),
.B(n_493),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_573),
.A2(n_372),
.B1(n_379),
.B2(n_381),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_710),
.B(n_562),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_623),
.B(n_201),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_206),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_573),
.B(n_556),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_674),
.B(n_525),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_572),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_629),
.A2(n_289),
.B1(n_246),
.B2(n_255),
.Y(n_840)
);

AND2x4_ASAP7_75t_SL g841 ( 
.A(n_594),
.B(n_643),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_699),
.B(n_525),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_647),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_594),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_581),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_609),
.B(n_525),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_647),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_611),
.B(n_525),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_572),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_629),
.B(n_556),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_629),
.Y(n_851)
);

NAND3x1_ASAP7_75t_L g852 ( 
.A(n_663),
.B(n_384),
.C(n_371),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_575),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_643),
.A2(n_289),
.B1(n_255),
.B2(n_262),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_611),
.B(n_525),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_613),
.B(n_525),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_613),
.B(n_525),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_575),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_577),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_588),
.B(n_208),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_586),
.B(n_209),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_629),
.A2(n_296),
.B1(n_262),
.B2(n_280),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_577),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_629),
.B(n_556),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_629),
.A2(n_296),
.B1(n_280),
.B2(n_290),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_649),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_650),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_629),
.B(n_566),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_594),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_683),
.B(n_471),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_650),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_622),
.B(n_625),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_590),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_590),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_592),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_622),
.B(n_625),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_653),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_640),
.B(n_566),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_640),
.B(n_566),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_640),
.A2(n_290),
.B1(n_301),
.B2(n_305),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_640),
.B(n_525),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_640),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_683),
.B(n_535),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_592),
.Y(n_885)
);

BUFx8_ASAP7_75t_L g886 ( 
.A(n_688),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_593),
.B(n_214),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_630),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_653),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_690),
.B(n_259),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_640),
.B(n_259),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_812),
.B(n_685),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_730),
.B(n_640),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_873),
.A2(n_667),
.B(n_581),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_816),
.B(n_685),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_764),
.B(n_645),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_877),
.A2(n_693),
.B(n_690),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_839),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_738),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_877),
.A2(n_667),
.B(n_693),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_849),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_761),
.B(n_700),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_733),
.B(n_645),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_835),
.B(n_651),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_841),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_732),
.B(n_707),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_749),
.A2(n_667),
.B(n_696),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_753),
.A2(n_697),
.B(n_696),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_758),
.A2(n_701),
.B(n_697),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_768),
.A2(n_712),
.B(n_701),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_754),
.A2(n_713),
.B(n_712),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_766),
.B(n_587),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_780),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_747),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_762),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_886),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_773),
.A2(n_576),
.B(n_574),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_853),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_774),
.B(n_685),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_834),
.A2(n_576),
.B(n_574),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_858),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_836),
.B(n_651),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_752),
.B(n_709),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_738),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_846),
.A2(n_713),
.B(n_652),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_652),
.Y(n_926)
);

NOR2x1_ASAP7_75t_L g927 ( 
.A(n_723),
.B(n_632),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_829),
.A2(n_619),
.B(n_616),
.C(n_632),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_780),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_732),
.B(n_709),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_745),
.A2(n_677),
.B(n_607),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_859),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_846),
.A2(n_855),
.B(n_848),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_748),
.A2(n_677),
.B(n_607),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_652),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_837),
.A2(n_677),
.B(n_703),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_741),
.A2(n_685),
.B(n_720),
.C(n_721),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_755),
.B(n_656),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_831),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_738),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_850),
.A2(n_711),
.B(n_703),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_865),
.A2(n_711),
.B(n_703),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_738),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_SL g944 ( 
.A1(n_741),
.A2(n_301),
.B(n_383),
.C(n_380),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_842),
.A2(n_607),
.B(n_692),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_763),
.A2(n_662),
.B1(n_666),
.B2(n_637),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_841),
.B(n_688),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_848),
.A2(n_620),
.B(n_668),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_760),
.B(n_652),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_864),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_760),
.B(n_652),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_808),
.A2(n_720),
.B(n_665),
.C(n_679),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_888),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_774),
.B(n_652),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_755),
.B(n_626),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_759),
.B(n_720),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_842),
.A2(n_607),
.B(n_692),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_838),
.A2(n_607),
.B(n_692),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_726),
.Y(n_959)
);

NAND2x1_ASAP7_75t_L g960 ( 
.A(n_731),
.B(n_603),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_759),
.B(n_720),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_869),
.A2(n_714),
.B(n_711),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_818),
.B(n_663),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_763),
.Y(n_964)
);

AO22x1_ASAP7_75t_L g965 ( 
.A1(n_805),
.A2(n_652),
.B1(n_360),
.B2(n_358),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_874),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_855),
.A2(n_620),
.B(n_603),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_727),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_774),
.B(n_714),
.Y(n_969)
);

INVx6_ASAP7_75t_L g970 ( 
.A(n_763),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_731),
.B(n_692),
.Y(n_971)
);

OAI22xp33_ASAP7_75t_L g972 ( 
.A1(n_763),
.A2(n_318),
.B1(n_306),
.B2(n_305),
.Y(n_972)
);

INVx3_ASAP7_75t_SL g973 ( 
.A(n_722),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_862),
.A2(n_714),
.B(n_715),
.C(n_306),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_SL g975 ( 
.A1(n_888),
.A2(n_320),
.B1(n_230),
.B2(n_223),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_838),
.A2(n_728),
.B(n_856),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_742),
.B(n_715),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_814),
.B(n_715),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_814),
.B(n_603),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_776),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_856),
.A2(n_692),
.B(n_664),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_875),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_318),
.B1(n_367),
.B2(n_368),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_876),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_777),
.B(n_725),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_793),
.A2(n_605),
.B1(n_602),
.B2(n_679),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_879),
.A2(n_664),
.B(n_658),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_778),
.A2(n_605),
.B1(n_602),
.B2(n_665),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_729),
.B(n_658),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_857),
.A2(n_821),
.B(n_880),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_857),
.A2(n_694),
.B(n_664),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_885),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_767),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_792),
.B(n_539),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_795),
.A2(n_694),
.B(n_670),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_818),
.B(n_308),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_884),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_795),
.A2(n_694),
.B(n_670),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_736),
.B(n_215),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_795),
.A2(n_815),
.B(n_882),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_746),
.B(n_668),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_739),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_746),
.B(n_692),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_778),
.A2(n_695),
.B(n_367),
.C(n_380),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_815),
.A2(n_676),
.B(n_695),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_815),
.A2(n_676),
.B(n_708),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_794),
.A2(n_719),
.B(n_708),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_801),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_887),
.A2(n_308),
.B(n_719),
.C(n_541),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_734),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_786),
.A2(n_705),
.B(n_702),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_746),
.B(n_342),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_767),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_L g1014 ( 
.A(n_736),
.B(n_539),
.C(n_569),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_751),
.B(n_686),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_860),
.A2(n_265),
.B(n_221),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_757),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_844),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_794),
.A2(n_705),
.B(n_702),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_765),
.B(n_686),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_890),
.A2(n_549),
.B(n_569),
.C(n_559),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_890),
.A2(n_547),
.B(n_559),
.C(n_557),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_772),
.Y(n_1023)
);

NAND2x2_ASAP7_75t_L g1024 ( 
.A(n_799),
.B(n_222),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_794),
.A2(n_689),
.B(n_499),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_801),
.B(n_845),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_782),
.B(n_689),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_788),
.A2(n_496),
.B(n_515),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_L g1029 ( 
.A(n_756),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_743),
.A2(n_507),
.B(n_499),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_809),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_743),
.A2(n_507),
.B(n_496),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_871),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_783),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_801),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_784),
.B(n_540),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_735),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_767),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_750),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_832),
.A2(n_517),
.B(n_496),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_823),
.B(n_361),
.C(n_234),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_798),
.B(n_891),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_740),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_851),
.A2(n_515),
.B(n_496),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_787),
.A2(n_517),
.B(n_515),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_883),
.A2(n_517),
.B(n_515),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_807),
.A2(n_517),
.B(n_557),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_845),
.B(n_371),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_750),
.A2(n_549),
.B1(n_547),
.B2(n_540),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_767),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_845),
.B(n_342),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_731),
.A2(n_541),
.B1(n_349),
.B2(n_348),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_737),
.B(n_478),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_790),
.A2(n_542),
.B(n_537),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_791),
.B(n_542),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_845),
.B(n_480),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_785),
.B(n_231),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_796),
.A2(n_493),
.B(n_537),
.Y(n_1058)
);

OAI321xp33_ASAP7_75t_L g1059 ( 
.A1(n_854),
.A2(n_384),
.A3(n_489),
.B1(n_480),
.B2(n_481),
.C(n_484),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_825),
.B(n_342),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_806),
.A2(n_493),
.B(n_542),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_810),
.A2(n_537),
.B(n_531),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_825),
.B(n_827),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_886),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_744),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_813),
.B(n_526),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_817),
.B(n_526),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_819),
.B(n_531),
.Y(n_1068)
);

BUFx8_ASAP7_75t_L g1069 ( 
.A(n_844),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_781),
.A2(n_789),
.B(n_769),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_852),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_827),
.B(n_481),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_781),
.A2(n_531),
.B(n_529),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_820),
.B(n_529),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_789),
.A2(n_531),
.B(n_529),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_744),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_826),
.B(n_529),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_912),
.B(n_771),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_916),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_896),
.B(n_830),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1013),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_935),
.A2(n_724),
.B(n_881),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_923),
.A2(n_724),
.B(n_878),
.C(n_872),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_926),
.A2(n_800),
.B(n_840),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1016),
.A2(n_889),
.B(n_878),
.C(n_872),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_924),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_939),
.B(n_804),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_919),
.B(n_771),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1070),
.A2(n_863),
.B(n_866),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_892),
.B(n_775),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_904),
.B(n_775),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_928),
.A2(n_889),
.B(n_779),
.C(n_868),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1063),
.A2(n_824),
.B(n_868),
.C(n_867),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_914),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_937),
.A2(n_779),
.B(n_867),
.C(n_861),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_903),
.B(n_797),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1002),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_999),
.A2(n_797),
.B(n_861),
.C(n_802),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1013),
.Y(n_1099)
);

AO21x1_ASAP7_75t_L g1100 ( 
.A1(n_983),
.A2(n_907),
.B(n_922),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_893),
.A2(n_824),
.B(n_847),
.Y(n_1101)
);

AOI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_1072),
.A2(n_803),
.B(n_811),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_895),
.B(n_357),
.C(n_270),
.Y(n_1103)
);

INVx6_ASAP7_75t_L g1104 ( 
.A(n_1069),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_894),
.A2(n_811),
.B(n_847),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_802),
.B(n_803),
.C(n_828),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_930),
.A2(n_828),
.B(n_843),
.C(n_833),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_985),
.B(n_843),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1033),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1039),
.B(n_844),
.Y(n_1110)
);

INVx3_ASAP7_75t_SL g1111 ( 
.A(n_913),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_946),
.A2(n_852),
.B1(n_870),
.B2(n_344),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_959),
.B(n_870),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_SL g1114 ( 
.A1(n_973),
.A2(n_722),
.B1(n_822),
.B2(n_343),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_949),
.A2(n_334),
.B(n_285),
.C(n_298),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1017),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_SL g1117 ( 
.A(n_1008),
.B(n_870),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_968),
.B(n_1031),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1013),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_953),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_915),
.B(n_258),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_997),
.B(n_304),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1023),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1034),
.B(n_310),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1029),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1076),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1048),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_994),
.B(n_311),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_951),
.A2(n_354),
.B1(n_324),
.B2(n_326),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1071),
.B(n_312),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_L g1131 ( 
.A(n_924),
.B(n_330),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_929),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1056),
.B(n_484),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_980),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1035),
.B(n_344),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_931),
.A2(n_934),
.B(n_917),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_947),
.A2(n_364),
.B1(n_385),
.B2(n_373),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_978),
.B(n_370),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1050),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1037),
.B(n_365),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_924),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_920),
.A2(n_490),
.B(n_73),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1053),
.B(n_353),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_1041),
.Y(n_1145)
);

OAI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1057),
.A2(n_337),
.B1(n_332),
.B2(n_331),
.C(n_19),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_SL g1147 ( 
.A(n_938),
.B(n_12),
.C(n_14),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_955),
.B(n_16),
.C(n_21),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_940),
.Y(n_1149)
);

AOI222xp33_ASAP7_75t_L g1150 ( 
.A1(n_1059),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_26),
.C2(n_29),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1010),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1043),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1060),
.A2(n_1012),
.B(n_1051),
.C(n_972),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_933),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1048),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1037),
.B(n_940),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_940),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_996),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_901),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_976),
.A2(n_31),
.B(n_38),
.C(n_40),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_954),
.A2(n_92),
.B(n_170),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_979),
.B(n_83),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_996),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_918),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1056),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1000),
.A2(n_95),
.B(n_169),
.Y(n_1166)
);

O2A1O1Ixp5_ASAP7_75t_L g1167 ( 
.A1(n_907),
.A2(n_94),
.B(n_162),
.C(n_154),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_996),
.A2(n_1049),
.B1(n_1036),
.B2(n_921),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_SL g1169 ( 
.A(n_1014),
.B(n_46),
.C(n_50),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_975),
.B(n_46),
.Y(n_1170)
);

INVx8_ASAP7_75t_L g1171 ( 
.A(n_1050),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_932),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1000),
.A2(n_179),
.B(n_80),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_902),
.B(n_51),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1050),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_990),
.A2(n_72),
.B(n_146),
.C(n_140),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_950),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_906),
.B(n_71),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_927),
.A2(n_153),
.B1(n_134),
.B2(n_133),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_984),
.B(n_114),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_992),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_969),
.B(n_113),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1007),
.A2(n_108),
.B(n_106),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1065),
.Y(n_1184)
);

O2A1O1Ixp5_ASAP7_75t_L g1185 ( 
.A1(n_974),
.A2(n_51),
.B(n_56),
.C(n_57),
.Y(n_1185)
);

AO22x1_ASAP7_75t_L g1186 ( 
.A1(n_1069),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1001),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_986),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_965),
.A2(n_59),
.B1(n_69),
.B2(n_1052),
.C(n_1004),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_898),
.B(n_966),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_982),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_900),
.A2(n_936),
.B(n_971),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_900),
.A2(n_936),
.B(n_971),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1064),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_956),
.B(n_961),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_977),
.B(n_899),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1018),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_899),
.A2(n_970),
.B1(n_943),
.B2(n_964),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1009),
.A2(n_1026),
.B(n_910),
.C(n_908),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1055),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_905),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_905),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_943),
.B(n_964),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_993),
.B(n_1038),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1015),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1020),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_970),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1042),
.A2(n_925),
.B(n_967),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1021),
.B(n_1022),
.C(n_988),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_970),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_944),
.A2(n_952),
.B1(n_908),
.B2(n_909),
.C(n_910),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_989),
.B(n_1003),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_960),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_987),
.A2(n_962),
.B(n_942),
.Y(n_1214)
);

CKINVDCx8_ASAP7_75t_R g1215 ( 
.A(n_1024),
.Y(n_1215)
);

BUFx4f_ASAP7_75t_L g1216 ( 
.A(n_897),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_987),
.A2(n_962),
.B(n_941),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1027),
.B(n_1077),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1066),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_941),
.A2(n_942),
.B(n_1028),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_991),
.A2(n_957),
.B(n_945),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1067),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1030),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_909),
.B(n_911),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1030),
.A2(n_1005),
.B1(n_1068),
.B2(n_1074),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_SL g1226 ( 
.A1(n_911),
.A2(n_1040),
.B(n_1032),
.C(n_998),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_958),
.B(n_1040),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1073),
.A2(n_1075),
.B(n_1032),
.C(n_1025),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1073),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1075),
.B(n_981),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1025),
.A2(n_995),
.B(n_998),
.C(n_1007),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1171),
.B(n_995),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1078),
.B(n_1062),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1176),
.A2(n_1047),
.B(n_1058),
.C(n_1061),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1223),
.A2(n_1045),
.B(n_1019),
.Y(n_1235)
);

OAI22x1_ASAP7_75t_L g1236 ( 
.A1(n_1112),
.A2(n_948),
.B1(n_1019),
.B2(n_1006),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1216),
.A2(n_1080),
.B1(n_1195),
.B2(n_1091),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_SL g1238 ( 
.A1(n_1160),
.A2(n_1178),
.B(n_1115),
.C(n_1180),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1180),
.A2(n_1044),
.B(n_1046),
.C(n_1054),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1224),
.A2(n_1089),
.B(n_1082),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1104),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1135),
.B(n_1117),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1084),
.A2(n_1199),
.B(n_1101),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1133),
.B(n_1090),
.Y(n_1245)
);

NAND3x1_ASAP7_75t_L g1246 ( 
.A(n_1170),
.B(n_1113),
.C(n_1110),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1132),
.B(n_1109),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1146),
.A2(n_1154),
.B1(n_1130),
.B2(n_1188),
.C(n_1169),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1120),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1116),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1136),
.A2(n_1217),
.B(n_1214),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1221),
.A2(n_1092),
.B(n_1220),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1111),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1231),
.B(n_1225),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1153),
.A2(n_1216),
.B(n_1173),
.C(n_1166),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1215),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1123),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1094),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1187),
.B(n_1138),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1211),
.A2(n_1095),
.B(n_1173),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1133),
.B(n_1134),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1118),
.B(n_1132),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1166),
.A2(n_1145),
.B(n_1189),
.C(n_1087),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1159),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1164),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1202),
.Y(n_1267)
);

AO32x2_ASAP7_75t_L g1268 ( 
.A1(n_1168),
.A2(n_1225),
.A3(n_1158),
.B1(n_1163),
.B2(n_1129),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1183),
.A2(n_1143),
.B(n_1093),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1107),
.A2(n_1083),
.B(n_1162),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1209),
.A2(n_1098),
.B(n_1106),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1194),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1201),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1138),
.B(n_1200),
.Y(n_1274)
);

INVx6_ASAP7_75t_SL g1275 ( 
.A(n_1204),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1207),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1204),
.Y(n_1277)
);

AO32x2_ASAP7_75t_L g1278 ( 
.A1(n_1168),
.A2(n_1158),
.A3(n_1163),
.B1(n_1129),
.B2(n_1137),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1201),
.B(n_1125),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1172),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1128),
.B(n_1144),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1226),
.A2(n_1096),
.B(n_1108),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1165),
.A2(n_1088),
.B1(n_1103),
.B2(n_1150),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1140),
.A2(n_1148),
.B(n_1147),
.C(n_1121),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1150),
.A2(n_1174),
.B1(n_1114),
.B2(n_1088),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1177),
.A2(n_1181),
.B1(n_1198),
.B2(n_1191),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1085),
.A2(n_1182),
.B(n_1196),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1096),
.A2(n_1102),
.B(n_1229),
.C(n_1190),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1201),
.B(n_1117),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1126),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1218),
.B(n_1124),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1142),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1155),
.B(n_1122),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1212),
.A2(n_1102),
.B(n_1227),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_1203),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1230),
.A2(n_1161),
.B(n_1156),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1179),
.A2(n_1213),
.B(n_1081),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1135),
.B(n_1185),
.C(n_1131),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1167),
.A2(n_1184),
.B(n_1152),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1213),
.A2(n_1171),
.B(n_1151),
.Y(n_1303)
);

AND2x6_ASAP7_75t_SL g1304 ( 
.A(n_1079),
.B(n_1104),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1213),
.A2(n_1171),
.B(n_1157),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1210),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1086),
.A2(n_1149),
.B(n_1157),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1186),
.A2(n_1086),
.B(n_1149),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1197),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1081),
.A2(n_1099),
.B(n_1119),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1099),
.A2(n_1119),
.B(n_1139),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_SL g1312 ( 
.A(n_1119),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1175),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1208),
.A2(n_733),
.B(n_730),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1189),
.B(n_923),
.C(n_816),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1135),
.B(n_844),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1111),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1078),
.B(n_730),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1094),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1201),
.B(n_1008),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1220),
.B(n_1214),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1153),
.A2(n_733),
.B(n_923),
.C(n_816),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1220),
.A2(n_1217),
.B(n_1214),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1111),
.Y(n_1326)
);

AOI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1146),
.A2(n_923),
.B1(n_812),
.B2(n_816),
.C(n_912),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_1197),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1097),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1201),
.B(n_1008),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1208),
.A2(n_733),
.B(n_730),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1220),
.B(n_1214),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1216),
.A2(n_733),
.B1(n_730),
.B2(n_923),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1337)
);

AND2x6_ASAP7_75t_L g1338 ( 
.A(n_1187),
.B(n_738),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1197),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1197),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1220),
.B(n_1214),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1097),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1216),
.A2(n_733),
.B1(n_730),
.B2(n_923),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1154),
.A2(n_1188),
.B1(n_733),
.B2(n_808),
.C(n_1189),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1078),
.B(n_730),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1208),
.A2(n_733),
.B(n_730),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1097),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1120),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1132),
.B(n_912),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1097),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1353)
);

AO21x1_ASAP7_75t_L g1354 ( 
.A1(n_1154),
.A2(n_733),
.B(n_1173),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1097),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1153),
.A2(n_733),
.B(n_923),
.C(n_816),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1220),
.B(n_1214),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1220),
.A2(n_1217),
.B(n_1214),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1111),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1133),
.B(n_776),
.Y(n_1360)
);

OAI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1130),
.A2(n_816),
.B(n_812),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1097),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1208),
.A2(n_733),
.B(n_1084),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1100),
.A2(n_1228),
.A3(n_1220),
.B(n_1214),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1094),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1105),
.A2(n_1193),
.B(n_1192),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1171),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1097),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1201),
.B(n_1125),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1118),
.B(n_912),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1097),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1208),
.A2(n_733),
.B(n_730),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1094),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1135),
.A2(n_923),
.B1(n_766),
.B2(n_912),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1097),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1146),
.A2(n_923),
.B(n_816),
.C(n_812),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1220),
.A2(n_1217),
.B(n_1214),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1208),
.A2(n_733),
.B(n_1084),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1153),
.A2(n_733),
.B(n_923),
.C(n_816),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1097),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1133),
.B(n_776),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1078),
.B(n_730),
.Y(n_1383)
);

NOR4xp25_ASAP7_75t_L g1384 ( 
.A(n_1154),
.B(n_1188),
.C(n_1169),
.D(n_1160),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1097),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1171),
.B(n_1201),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1078),
.B(n_730),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1223),
.A2(n_639),
.B(n_1208),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1304),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1258),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1277),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1243),
.A2(n_1315),
.B1(n_1316),
.B2(n_1336),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1243),
.A2(n_1315),
.B1(n_1316),
.B2(n_1343),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1320),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1304),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1351),
.A2(n_1361),
.B1(n_1375),
.B2(n_1300),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1265),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1280),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1366),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1361),
.A2(n_1300),
.B1(n_1292),
.B2(n_1360),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1327),
.A2(n_1248),
.B1(n_1354),
.B2(n_1286),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1286),
.A2(n_1274),
.B1(n_1371),
.B2(n_1334),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1301),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1314),
.A2(n_1373),
.B1(n_1346),
.B2(n_1260),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1250),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1266),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1331),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1342),
.Y(n_1408)
);

INVx3_ASAP7_75t_SL g1409 ( 
.A(n_1309),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1283),
.A2(n_1237),
.B1(n_1281),
.B2(n_1387),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1349),
.Y(n_1411)
);

BUFx12f_ASAP7_75t_L g1412 ( 
.A(n_1256),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1318),
.A2(n_1383),
.B1(n_1345),
.B2(n_1363),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1363),
.A2(n_1379),
.B1(n_1261),
.B2(n_1270),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1295),
.A2(n_1366),
.B1(n_1374),
.B2(n_1257),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1379),
.A2(n_1261),
.B1(n_1382),
.B2(n_1377),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1255),
.A2(n_1264),
.B1(n_1323),
.B2(n_1356),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1245),
.A2(n_1262),
.B1(n_1338),
.B2(n_1246),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1368),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1263),
.A2(n_1233),
.B1(n_1285),
.B2(n_1385),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1352),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1338),
.A2(n_1278),
.B1(n_1241),
.B2(n_1253),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1355),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1362),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1368),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1386),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1339),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1369),
.A2(n_1376),
.B1(n_1381),
.B2(n_1372),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1291),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1329),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1302),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1287),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1240),
.A2(n_1344),
.B1(n_1290),
.B2(n_1271),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1340),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1254),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1317),
.A2(n_1326),
.B1(n_1359),
.B2(n_1374),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1386),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1247),
.A2(n_1267),
.B1(n_1279),
.B2(n_1370),
.Y(n_1439)
);

CKINVDCx6p67_ASAP7_75t_R g1440 ( 
.A(n_1329),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1344),
.A2(n_1271),
.B1(n_1296),
.B2(n_1288),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1350),
.B2(n_1249),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1312),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1380),
.B(n_1284),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1277),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1278),
.A2(n_1384),
.B1(n_1244),
.B2(n_1332),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1272),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1278),
.A2(n_1384),
.B1(n_1244),
.B2(n_1365),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1276),
.B(n_1279),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1386),
.Y(n_1450)
);

BUFx4_ASAP7_75t_SL g1451 ( 
.A(n_1232),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1254),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1254),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1328),
.A2(n_1388),
.B1(n_1337),
.B2(n_1348),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1322),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1370),
.B(n_1289),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1297),
.A2(n_1299),
.B1(n_1333),
.B2(n_1321),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1273),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1353),
.A2(n_1282),
.B1(n_1338),
.B2(n_1325),
.Y(n_1459)
);

INVx5_ASAP7_75t_L g1460 ( 
.A(n_1313),
.Y(n_1460)
);

CKINVDCx6p67_ASAP7_75t_R g1461 ( 
.A(n_1232),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1306),
.B(n_1268),
.Y(n_1462)
);

BUFx4_ASAP7_75t_R g1463 ( 
.A(n_1275),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1293),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1232),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1307),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1293),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1294),
.Y(n_1468)
);

BUFx4_ASAP7_75t_SL g1469 ( 
.A(n_1310),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1298),
.B(n_1294),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1268),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1268),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1303),
.A2(n_1305),
.B1(n_1311),
.B2(n_1235),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1325),
.A2(n_1358),
.B1(n_1378),
.B2(n_1236),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1238),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1322),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1335),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1335),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1239),
.Y(n_1479)
);

CKINVDCx6p67_ASAP7_75t_R g1480 ( 
.A(n_1234),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1335),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1341),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_L g1483 ( 
.A(n_1341),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1341),
.B(n_1364),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1252),
.B(n_1378),
.Y(n_1485)
);

INVx8_ASAP7_75t_L g1486 ( 
.A(n_1358),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1251),
.A2(n_1269),
.B1(n_1242),
.B2(n_1319),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1357),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1357),
.Y(n_1489)
);

INVx8_ASAP7_75t_L g1490 ( 
.A(n_1364),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1324),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1330),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1347),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1367),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1243),
.A2(n_923),
.B1(n_766),
.B2(n_1315),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1245),
.B(n_1360),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1361),
.A2(n_923),
.B1(n_766),
.B2(n_1327),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1243),
.A2(n_923),
.B1(n_766),
.B2(n_1315),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1243),
.A2(n_923),
.B1(n_766),
.B2(n_1315),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1245),
.B(n_1360),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1368),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1320),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1361),
.A2(n_1327),
.B(n_1377),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1318),
.B(n_1345),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1258),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1375),
.A2(n_1327),
.B1(n_1361),
.B2(n_1315),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1320),
.Y(n_1509)
);

BUFx8_ASAP7_75t_L g1510 ( 
.A(n_1312),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1258),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1375),
.A2(n_1327),
.B1(n_1361),
.B2(n_1315),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1386),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1320),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1320),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1304),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1320),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1368),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1259),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1258),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1361),
.A2(n_923),
.B1(n_766),
.B2(n_1327),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1258),
.Y(n_1526)
);

CKINVDCx11_ASAP7_75t_R g1527 ( 
.A(n_1304),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1361),
.A2(n_1327),
.B1(n_1315),
.B2(n_1248),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1368),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1320),
.Y(n_1530)
);

BUFx10_ASAP7_75t_L g1531 ( 
.A(n_1304),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1258),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1304),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1481),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1417),
.A2(n_1505),
.B(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1476),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1462),
.B(n_1471),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1432),
.A2(n_1453),
.A3(n_1452),
.B(n_1436),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1465),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1405),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1486),
.B(n_1490),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1506),
.B(n_1413),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1493),
.A2(n_1432),
.B(n_1484),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1508),
.A2(n_1512),
.B1(n_1528),
.B2(n_1497),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1405),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1477),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1399),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1413),
.B(n_1497),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1496),
.B(n_1502),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1436),
.Y(n_1550)
);

INVx11_ASAP7_75t_L g1551 ( 
.A(n_1443),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1453),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1481),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1455),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1472),
.B(n_1446),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1499),
.B(n_1515),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1408),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1513),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1448),
.A2(n_1474),
.B(n_1459),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1483),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1482),
.B(n_1478),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1498),
.A2(n_1524),
.B1(n_1500),
.B2(n_1495),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1478),
.Y(n_1563)
);

AO21x1_ASAP7_75t_SL g1564 ( 
.A1(n_1401),
.A2(n_1441),
.B(n_1434),
.Y(n_1564)
);

OAI222xp33_ASAP7_75t_L g1565 ( 
.A1(n_1499),
.A2(n_1525),
.B1(n_1528),
.B2(n_1521),
.C1(n_1517),
.C2(n_1515),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1485),
.A2(n_1487),
.B(n_1454),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1422),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1488),
.B(n_1416),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1501),
.B(n_1415),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1474),
.A2(n_1459),
.B(n_1454),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1425),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1485),
.A2(n_1487),
.B(n_1473),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1517),
.A2(n_1525),
.B1(n_1521),
.B2(n_1401),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1412),
.B(n_1428),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1403),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1389),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1486),
.B(n_1490),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1513),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1416),
.B(n_1423),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1483),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1433),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1414),
.B(n_1489),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1444),
.A2(n_1402),
.B1(n_1396),
.B2(n_1410),
.C(n_1404),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1475),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1443),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1427),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1414),
.B(n_1489),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1392),
.A2(n_1393),
.B(n_1404),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1394),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1406),
.Y(n_1591)
);

NOR2x1_ASAP7_75t_R g1592 ( 
.A(n_1527),
.B(n_1533),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1412),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1407),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1427),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1479),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1597)
);

AOI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1457),
.A2(n_1470),
.B(n_1466),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1507),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_SL g1600 ( 
.A(n_1479),
.B(n_1513),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1513),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1411),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1402),
.A2(n_1410),
.B(n_1400),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1486),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1424),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1461),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1504),
.B(n_1519),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1456),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1430),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1526),
.Y(n_1610)
);

AO21x1_ASAP7_75t_SL g1611 ( 
.A1(n_1441),
.A2(n_1434),
.B(n_1420),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_SL g1612 ( 
.A(n_1395),
.B(n_1518),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1390),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1480),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1397),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1439),
.A2(n_1518),
.B1(n_1395),
.B2(n_1437),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1429),
.B(n_1523),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1398),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1464),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1443),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1429),
.A2(n_1532),
.B(n_1511),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1449),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1440),
.A2(n_1467),
.B1(n_1516),
.B2(n_1530),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1442),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1409),
.B(n_1509),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1391),
.B(n_1445),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1391),
.A2(n_1445),
.B(n_1468),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1451),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1418),
.B(n_1438),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1503),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1469),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1503),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1438),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1514),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1460),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1458),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1426),
.B(n_1529),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1460),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1426),
.B(n_1529),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1510),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1435),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1603),
.A2(n_1419),
.B(n_1421),
.C(n_1533),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1562),
.A2(n_1520),
.B(n_1460),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1581),
.B(n_1419),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1544),
.A2(n_1527),
.B(n_1463),
.Y(n_1645)
);

NOR4xp25_ASAP7_75t_SL g1646 ( 
.A(n_1569),
.B(n_1531),
.C(n_1463),
.D(n_1510),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1566),
.A2(n_1531),
.B(n_1450),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1549),
.B(n_1409),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1591),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1566),
.A2(n_1510),
.B(n_1431),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1565),
.A2(n_1431),
.B(n_1447),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1597),
.B(n_1583),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1584),
.A2(n_1589),
.B1(n_1556),
.B2(n_1574),
.C(n_1548),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1542),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1574),
.A2(n_1598),
.B(n_1624),
.Y(n_1655)
);

AND2x6_ASAP7_75t_L g1656 ( 
.A(n_1580),
.B(n_1558),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1582),
.B(n_1608),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1561),
.B(n_1572),
.Y(n_1658)
);

AND2x2_ASAP7_75t_SL g1659 ( 
.A(n_1597),
.B(n_1608),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1561),
.B(n_1576),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1547),
.B(n_1641),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1555),
.B(n_1617),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1590),
.A2(n_1616),
.B(n_1624),
.C(n_1628),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1573),
.A2(n_1598),
.B(n_1535),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1641),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1577),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1568),
.A2(n_1588),
.B1(n_1629),
.B2(n_1564),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1541),
.B(n_1578),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1573),
.A2(n_1627),
.B(n_1546),
.Y(n_1672)
);

AO32x2_ASAP7_75t_L g1673 ( 
.A1(n_1587),
.A2(n_1632),
.A3(n_1630),
.B1(n_1537),
.B2(n_1611),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1631),
.A2(n_1623),
.B(n_1636),
.C(n_1628),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1629),
.B(n_1633),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1613),
.B(n_1615),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_SL g1677 ( 
.A(n_1611),
.B(n_1564),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1619),
.B(n_1634),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_SL g1679 ( 
.A1(n_1631),
.A2(n_1614),
.B(n_1585),
.C(n_1596),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1594),
.B(n_1602),
.Y(n_1680)
);

BUFx8_ASAP7_75t_L g1681 ( 
.A(n_1586),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1586),
.A2(n_1620),
.B1(n_1640),
.B2(n_1606),
.C(n_1614),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1612),
.A2(n_1535),
.B1(n_1575),
.B2(n_1606),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1594),
.B(n_1602),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1585),
.A2(n_1640),
.B1(n_1620),
.B2(n_1551),
.Y(n_1685)
);

A2O1A1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1612),
.A2(n_1585),
.B(n_1534),
.C(n_1596),
.Y(n_1686)
);

AO21x1_ASAP7_75t_L g1687 ( 
.A1(n_1618),
.A2(n_1605),
.B(n_1609),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1596),
.A2(n_1595),
.B(n_1625),
.C(n_1560),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1540),
.B(n_1545),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1610),
.A2(n_1626),
.B1(n_1536),
.B2(n_1571),
.C(n_1567),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1637),
.A2(n_1639),
.B(n_1635),
.C(n_1638),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1627),
.A2(n_1553),
.B(n_1560),
.Y(n_1693)
);

AOI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1604),
.A2(n_1638),
.B(n_1635),
.Y(n_1694)
);

AO32x2_ASAP7_75t_L g1695 ( 
.A1(n_1559),
.A2(n_1621),
.A3(n_1538),
.B1(n_1536),
.B2(n_1552),
.Y(n_1695)
);

OAI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1570),
.A2(n_1559),
.B(n_1621),
.C(n_1610),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1695),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1695),
.B(n_1570),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1678),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1673),
.B(n_1559),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1673),
.B(n_1543),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1673),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1653),
.A2(n_1539),
.B1(n_1593),
.B2(n_1595),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1687),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1543),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1642),
.A2(n_1600),
.B(n_1592),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1662),
.B(n_1621),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1654),
.B(n_1683),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1655),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1657),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1665),
.B(n_1550),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1651),
.A2(n_1593),
.B1(n_1595),
.B2(n_1626),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1649),
.Y(n_1714)
);

OAI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1668),
.A2(n_1682),
.B1(n_1683),
.B2(n_1663),
.C1(n_1660),
.C2(n_1671),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1662),
.B(n_1538),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1657),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1651),
.A2(n_1601),
.B1(n_1579),
.B2(n_1558),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1693),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1655),
.B(n_1604),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1667),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1680),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1670),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1690),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1658),
.B(n_1538),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1645),
.A2(n_1643),
.B1(n_1646),
.B2(n_1659),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1684),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1664),
.A2(n_1626),
.B1(n_1557),
.B2(n_1599),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1669),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1714),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1702),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1717),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1700),
.B(n_1647),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1700),
.B(n_1702),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1709),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1701),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1714),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1701),
.B(n_1647),
.Y(n_1738)
);

AOI31xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1708),
.A2(n_1646),
.A3(n_1688),
.B(n_1648),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1697),
.B(n_1696),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1712),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1701),
.B(n_1675),
.Y(n_1745)
);

INVx5_ASAP7_75t_L g1746 ( 
.A(n_1723),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1698),
.B(n_1650),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1704),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1705),
.A2(n_1563),
.B(n_1554),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1698),
.B(n_1669),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1703),
.A2(n_1645),
.B1(n_1674),
.B2(n_1689),
.C(n_1685),
.Y(n_1751)
);

AOI211xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1726),
.A2(n_1679),
.B(n_1685),
.C(n_1661),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1729),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1703),
.A2(n_1656),
.B1(n_1652),
.B2(n_1681),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

OAI31xp33_ASAP7_75t_L g1756 ( 
.A1(n_1715),
.A2(n_1726),
.A3(n_1708),
.B(n_1713),
.Y(n_1756)
);

OAI211xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1710),
.A2(n_1692),
.B(n_1691),
.C(n_1676),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1725),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1736),
.B(n_1720),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1736),
.B(n_1720),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1730),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1730),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1740),
.B(n_1707),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1755),
.B(n_1711),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1737),
.Y(n_1766)
);

BUFx2_ASAP7_75t_SL g1767 ( 
.A(n_1746),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1755),
.B(n_1722),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1736),
.B(n_1724),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1731),
.B(n_1734),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1732),
.B(n_1722),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1731),
.B(n_1734),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1753),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1732),
.B(n_1727),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1757),
.B(n_1751),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1737),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1735),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1740),
.B(n_1707),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1741),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1749),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.B(n_1733),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1753),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1749),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1740),
.B(n_1716),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1753),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1733),
.B(n_1758),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1735),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1743),
.B(n_1699),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_L g1790 ( 
.A(n_1756),
.B(n_1710),
.C(n_1706),
.D(n_1728),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1778),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1778),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1788),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1770),
.B(n_1746),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1788),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1790),
.B(n_1742),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1763),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1764),
.B(n_1744),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1763),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1764),
.B(n_1744),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1764),
.B(n_1744),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1773),
.B(n_1756),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1770),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1773),
.B(n_1738),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1776),
.B(n_1771),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1761),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1770),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1776),
.B(n_1738),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1779),
.B(n_1742),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1761),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1772),
.B(n_1750),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1761),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1772),
.B(n_1750),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1771),
.B(n_1738),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1775),
.B(n_1699),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1762),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1762),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1772),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1762),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1759),
.B(n_1750),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1766),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1766),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1766),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1779),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1777),
.Y(n_1825)
);

AND2x4_ASAP7_75t_SL g1826 ( 
.A(n_1759),
.B(n_1754),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1777),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1777),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1780),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1779),
.B(n_1748),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1775),
.B(n_1745),
.Y(n_1831)
);

NOR3xp33_ASAP7_75t_L g1832 ( 
.A(n_1790),
.B(n_1751),
.C(n_1592),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1785),
.B(n_1765),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1774),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1769),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1780),
.Y(n_1836)
);

INVx3_ASAP7_75t_SL g1837 ( 
.A(n_1802),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1806),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1796),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_1718),
.B1(n_1754),
.B2(n_1713),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1804),
.A2(n_1752),
.B1(n_1739),
.B2(n_1746),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1805),
.B(n_1759),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1808),
.B(n_1760),
.Y(n_1843)
);

NAND2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1794),
.B(n_1746),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1811),
.B(n_1760),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1833),
.B(n_1785),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1833),
.B(n_1785),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1810),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1807),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1807),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1812),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1811),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1824),
.B(n_1760),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1813),
.B(n_1782),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1813),
.B(n_1782),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1721),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1791),
.B(n_1752),
.Y(n_1857)
);

AND2x2_ASAP7_75t_SL g1858 ( 
.A(n_1826),
.B(n_1723),
.Y(n_1858)
);

OAI31xp33_ASAP7_75t_L g1859 ( 
.A1(n_1826),
.A2(n_1739),
.A3(n_1748),
.B(n_1728),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1792),
.B(n_1789),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1820),
.B(n_1794),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1794),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1820),
.B(n_1782),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1797),
.A2(n_1786),
.B(n_1783),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1809),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1793),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1803),
.B(n_1786),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1795),
.B(n_1815),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1816),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1831),
.B(n_1721),
.Y(n_1870)
);

NAND2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1830),
.B(n_1746),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1809),
.B(n_1830),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1834),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1803),
.B(n_1818),
.Y(n_1874)
);

A2O1A1Ixp33_ASAP7_75t_SL g1875 ( 
.A1(n_1839),
.A2(n_1799),
.B(n_1797),
.C(n_1786),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1870),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_SL g1877 ( 
.A1(n_1841),
.A2(n_1859),
.B(n_1840),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1873),
.Y(n_1878)
);

AOI21xp33_ASAP7_75t_SL g1879 ( 
.A1(n_1837),
.A2(n_1666),
.B(n_1834),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1859),
.B(n_1746),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1840),
.A2(n_1818),
.B1(n_1718),
.B2(n_1767),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1849),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1837),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1862),
.B(n_1797),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1872),
.B(n_1798),
.Y(n_1885)
);

AOI21xp33_ASAP7_75t_L g1886 ( 
.A1(n_1857),
.A2(n_1865),
.B(n_1858),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1837),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1858),
.A2(n_1677),
.B1(n_1767),
.B2(n_1787),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1861),
.A2(n_1767),
.B1(n_1729),
.B2(n_1656),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1850),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1854),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1838),
.Y(n_1892)
);

OAI32xp33_ASAP7_75t_L g1893 ( 
.A1(n_1842),
.A2(n_1798),
.A3(n_1800),
.B1(n_1801),
.B2(n_1814),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1858),
.B(n_1799),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1866),
.B(n_1835),
.Y(n_1895)
);

OAI32xp33_ASAP7_75t_L g1896 ( 
.A1(n_1843),
.A2(n_1800),
.A3(n_1801),
.B1(n_1786),
.B2(n_1787),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1850),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1856),
.A2(n_1786),
.B(n_1783),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1854),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1868),
.A2(n_1835),
.B(n_1787),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1852),
.B(n_1789),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1883),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1887),
.B(n_1852),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1890),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1897),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1892),
.Y(n_1906)
);

AND2x4_ASAP7_75t_SL g1907 ( 
.A(n_1894),
.B(n_1861),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1882),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1892),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1876),
.B(n_1862),
.Y(n_1910)
);

OAI31xp33_ASAP7_75t_L g1911 ( 
.A1(n_1877),
.A2(n_1871),
.A3(n_1844),
.B(n_1872),
.Y(n_1911)
);

OAI221xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1900),
.A2(n_1895),
.B1(n_1885),
.B2(n_1878),
.C(n_1899),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1884),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1878),
.B(n_1845),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1879),
.B(n_1860),
.Y(n_1915)
);

NOR4xp25_ASAP7_75t_SL g1916 ( 
.A(n_1880),
.B(n_1848),
.C(n_1851),
.D(n_1838),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1879),
.B(n_1853),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1884),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1881),
.A2(n_1863),
.B1(n_1855),
.B2(n_1845),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1884),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1891),
.B(n_1863),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1891),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1908),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1911),
.B(n_1886),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1902),
.B(n_1899),
.Y(n_1925)
);

OAI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1917),
.A2(n_1888),
.B(n_1898),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1916),
.A2(n_1889),
.B1(n_1885),
.B2(n_1844),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1917),
.A2(n_1894),
.B(n_1844),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1908),
.B(n_1855),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1913),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1922),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1915),
.A2(n_1875),
.B(n_1896),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1920),
.B(n_1874),
.Y(n_1933)
);

INVxp33_ASAP7_75t_L g1934 ( 
.A(n_1915),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1925),
.B(n_1903),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1930),
.B(n_1918),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1932),
.A2(n_1912),
.B1(n_1919),
.B2(n_1910),
.C(n_1914),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1924),
.A2(n_1912),
.B1(n_1934),
.B2(n_1926),
.C(n_1896),
.Y(n_1938)
);

NOR4xp25_ASAP7_75t_L g1939 ( 
.A(n_1924),
.B(n_1905),
.C(n_1904),
.D(n_1906),
.Y(n_1939)
);

NOR2xp67_ASAP7_75t_L g1940 ( 
.A(n_1928),
.B(n_1921),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1929),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1923),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1933),
.B(n_1907),
.Y(n_1943)
);

OAI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1927),
.A2(n_1847),
.B1(n_1846),
.B2(n_1871),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1931),
.Y(n_1945)
);

BUFx10_ASAP7_75t_L g1946 ( 
.A(n_1945),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1938),
.A2(n_1901),
.B1(n_1847),
.B2(n_1846),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1935),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1937),
.A2(n_1909),
.B1(n_1873),
.B2(n_1874),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1942),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1940),
.A2(n_1893),
.B(n_1864),
.C(n_1869),
.Y(n_1951)
);

AOI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1939),
.A2(n_1893),
.B1(n_1851),
.B2(n_1869),
.C(n_1848),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1949),
.A2(n_1936),
.B1(n_1941),
.B2(n_1944),
.Y(n_1953)
);

NOR3xp33_ASAP7_75t_L g1954 ( 
.A(n_1948),
.B(n_1942),
.C(n_1943),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1950),
.Y(n_1955)
);

OAI211xp5_ASAP7_75t_SL g1956 ( 
.A1(n_1951),
.A2(n_1799),
.B(n_1786),
.C(n_1783),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1952),
.A2(n_1871),
.B(n_1864),
.Y(n_1957)
);

OAI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1947),
.A2(n_1867),
.B1(n_1774),
.B2(n_1783),
.C(n_1670),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1946),
.A2(n_1867),
.B(n_1763),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1951),
.A2(n_1774),
.B1(n_1783),
.B2(n_1670),
.C(n_1765),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1955),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1954),
.B(n_1953),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1958),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1959),
.Y(n_1964)
);

NOR2x1p5_ASAP7_75t_L g1965 ( 
.A(n_1960),
.B(n_1774),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1956),
.Y(n_1966)
);

AND3x1_ASAP7_75t_L g1967 ( 
.A(n_1962),
.B(n_1957),
.C(n_1774),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1961),
.B(n_1817),
.Y(n_1968)
);

NOR2x1p5_ASAP7_75t_L g1969 ( 
.A(n_1962),
.B(n_1681),
.Y(n_1969)
);

XNOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1965),
.B(n_1644),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1970),
.B(n_1964),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1971),
.Y(n_1972)
);

AOI311xp33_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1963),
.A3(n_1966),
.B(n_1968),
.C(n_1967),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1972),
.A2(n_1969),
.B1(n_1836),
.B2(n_1829),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1828),
.B1(n_1827),
.B2(n_1825),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1973),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1976),
.A2(n_1821),
.B(n_1819),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1975),
.A2(n_1823),
.B1(n_1822),
.B2(n_1763),
.C(n_1781),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1977),
.A2(n_1784),
.B(n_1781),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1979),
.A2(n_1978),
.B(n_1768),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1980),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1763),
.B1(n_1781),
.B2(n_1784),
.C(n_1780),
.Y(n_1982)
);

AOI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1763),
.B(n_1784),
.C(n_1781),
.Y(n_1983)
);


endmodule