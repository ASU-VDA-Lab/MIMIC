module fake_netlist_5_2072_n_1102 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1102);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1102;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_983;
wire n_725;
wire n_823;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1095;
wire n_976;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_995;
wire n_454;
wire n_961;
wire n_742;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_969;
wire n_866;
wire n_236;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_809;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_679;
wire n_710;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_952;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_67),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_162),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_84),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_60),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_95),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_55),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_46),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_47),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_88),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_5),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_112),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_107),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_14),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_2),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_75),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_100),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_161),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_136),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_124),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_118),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_126),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_26),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_19),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_80),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_4),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_82),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_166),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_233),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_220),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_217),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_228),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_202),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_217),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_220),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_224),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_207),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_214),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_230),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_201),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_204),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_244),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_244),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_245),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_245),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_201),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_306),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_239),
.B(n_223),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_278),
.B1(n_280),
.B2(n_273),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_295),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_289),
.A2(n_270),
.B1(n_205),
.B2(n_209),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_223),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_280),
.A2(n_241),
.B1(n_212),
.B2(n_213),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_283),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_221),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_269),
.B1(n_239),
.B2(n_242),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_269),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_295),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_261),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_310),
.B(n_221),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_262),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_296),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_221),
.Y(n_369)
);

INVx6_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_219),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_267),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_225),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_344),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_227),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_337),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_R g387 ( 
.A(n_337),
.B(n_319),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_329),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

NOR2x1p5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_229),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_329),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_333),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_357),
.B(n_319),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_372),
.B(n_282),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_374),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_364),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_364),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_364),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_364),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_368),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_368),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_368),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_368),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_368),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_338),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_318),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_370),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_366),
.A2(n_259),
.B1(n_237),
.B2(n_238),
.Y(n_426)
);

OR2x2_ASAP7_75t_SL g427 ( 
.A(n_370),
.B(n_318),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_370),
.Y(n_428)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_324),
.A2(n_240),
.B(n_235),
.Y(n_429)
);

CKINVDCx6p67_ASAP7_75t_R g430 ( 
.A(n_371),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_356),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_370),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_356),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_371),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_373),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_375),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_375),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_363),
.B(n_320),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_340),
.B(n_320),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_356),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_R g446 ( 
.A(n_360),
.B(n_246),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_362),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_350),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_342),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_362),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_383),
.B(n_369),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_377),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_347),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_351),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_388),
.B(n_352),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_347),
.Y(n_463)
);

AND2x4_ASAP7_75t_SL g464 ( 
.A(n_413),
.B(n_267),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_405),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_399),
.B(n_355),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_356),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_391),
.B(n_351),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_408),
.B(n_351),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_387),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_321),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_410),
.B(n_335),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_419),
.B(n_349),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_419),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_349),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_449),
.Y(n_492)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_397),
.B(n_353),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_398),
.B(n_353),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_410),
.B(n_335),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_401),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_412),
.B(n_321),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_321),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_417),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_410),
.B(n_332),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_431),
.B(n_332),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_380),
.B(n_332),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_404),
.B(n_353),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_446),
.B(n_321),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_385),
.B(n_345),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_403),
.B(n_345),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_402),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_413),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_448),
.A2(n_248),
.B1(n_258),
.B2(n_263),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_441),
.B(n_264),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_322),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_376),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_427),
.Y(n_530)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_406),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_439),
.B(n_322),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_381),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_481),
.B(n_322),
.Y(n_535)
);

AO22x2_ASAP7_75t_L g536 ( 
.A1(n_521),
.A2(n_424),
.B1(n_440),
.B2(n_389),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_481),
.B(n_322),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_390),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_520),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_487),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_389),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_330),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_490),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_490),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_469),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_508),
.B(n_330),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_496),
.B(n_330),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

AO22x2_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_268),
.B1(n_1),
.B2(n_2),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_499),
.B(n_461),
.C(n_474),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_505),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

BUFx8_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_483),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_520),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_499),
.A2(n_400),
.B1(n_395),
.B2(n_394),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_528),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_474),
.B(n_322),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_484),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_480),
.B(n_341),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

AO22x2_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_493),
.A2(n_323),
.B1(n_330),
.B2(n_341),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_480),
.B(n_341),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_457),
.B(n_461),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_450),
.B(n_323),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_454),
.A2(n_266),
.B1(n_267),
.B2(n_4),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_528),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_462),
.B(n_341),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_456),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_458),
.B(n_323),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_455),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_455),
.B(n_323),
.Y(n_587)
);

NAND3x1_ASAP7_75t_L g588 ( 
.A(n_533),
.B(n_0),
.C(n_3),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_465),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_530),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_534),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_496),
.B(n_323),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_534),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_466),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_459),
.B(n_6),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_488),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_489),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_514),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_492),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_502),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_515),
.B(n_30),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_506),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_540),
.B(n_510),
.Y(n_603)
);

NOR2x1_ASAP7_75t_R g604 ( 
.A(n_541),
.B(n_531),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_580),
.B(n_511),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_563),
.B(n_507),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_509),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_539),
.A2(n_532),
.B1(n_454),
.B2(n_494),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_502),
.B(n_504),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_581),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_535),
.A2(n_537),
.B(n_566),
.Y(n_611)
);

OAI21xp33_ASAP7_75t_L g612 ( 
.A1(n_574),
.A2(n_523),
.B(n_464),
.Y(n_612)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_600),
.A2(n_498),
.B(n_504),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_467),
.B(n_451),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_580),
.B(n_527),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_586),
.A2(n_467),
.B(n_451),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_472),
.B(n_498),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_565),
.A2(n_477),
.B(n_493),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_532),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_472),
.B(n_494),
.Y(n_620)
);

A2O1A1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_568),
.A2(n_477),
.B(n_470),
.C(n_468),
.Y(n_621)
);

HB1xp67_ASAP7_75t_SL g622 ( 
.A(n_558),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_572),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_587),
.A2(n_516),
.B(n_513),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_562),
.B(n_527),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_SL g626 ( 
.A(n_598),
.B(n_525),
.C(n_522),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_556),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_587),
.A2(n_516),
.B(n_513),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_573),
.A2(n_517),
.B(n_486),
.C(n_524),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_538),
.A2(n_517),
.B1(n_463),
.B2(n_512),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_556),
.A2(n_495),
.B(n_485),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_575),
.A2(n_500),
.B(n_497),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_584),
.A2(n_495),
.B(n_485),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_576),
.A2(n_595),
.B(n_524),
.C(n_577),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_585),
.A2(n_503),
.B(n_505),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_553),
.A2(n_501),
.B(n_471),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_542),
.B(n_475),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_564),
.B(n_471),
.C(n_531),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_559),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_545),
.A2(n_503),
.B(n_463),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_593),
.B(n_529),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_591),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_546),
.B(n_531),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_543),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_567),
.A2(n_486),
.B(n_503),
.C(n_529),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_572),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_579),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_594),
.A2(n_479),
.B(n_32),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_543),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_601),
.A2(n_479),
.B1(n_10),
.B2(n_11),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_581),
.A2(n_549),
.B(n_547),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_579),
.B(n_479),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_557),
.A2(n_33),
.B(n_31),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_569),
.A2(n_103),
.B1(n_198),
.B2(n_196),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_594),
.B(n_9),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_589),
.B(n_10),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_560),
.B(n_34),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_561),
.A2(n_38),
.B(n_35),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_582),
.A2(n_41),
.B(n_39),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_592),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_596),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_639),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_634),
.A2(n_599),
.B(n_597),
.C(n_601),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_642),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_619),
.B(n_544),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_642),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_608),
.A2(n_548),
.B1(n_550),
.B2(n_588),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_603),
.B(n_601),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_607),
.B(n_536),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_627),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_602),
.B(n_601),
.Y(n_672)
);

BUFx12f_ASAP7_75t_L g673 ( 
.A(n_642),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_606),
.A2(n_536),
.B1(n_570),
.B2(n_590),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_612),
.B(n_590),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_649),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_649),
.B(n_558),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_611),
.A2(n_570),
.B(n_552),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_605),
.B(n_610),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_629),
.A2(n_552),
.B1(n_12),
.B2(n_13),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_SL g682 ( 
.A1(n_648),
.A2(n_638),
.B(n_609),
.C(n_618),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_605),
.B(n_11),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_625),
.B(n_12),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_657),
.B(n_13),
.C(n_14),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_624),
.A2(n_110),
.B(n_195),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_621),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_622),
.Y(n_688)
);

CKINVDCx14_ASAP7_75t_R g689 ( 
.A(n_615),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_610),
.B(n_16),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_615),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_646),
.B(n_17),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_628),
.A2(n_633),
.B(n_620),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_R g694 ( 
.A(n_660),
.B(n_42),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_631),
.A2(n_114),
.B(n_192),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_SL g696 ( 
.A1(n_645),
.A2(n_113),
.B(n_191),
.C(n_189),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_644),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_641),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_637),
.B(n_18),
.Y(n_699)
);

BUFx8_ASAP7_75t_SL g700 ( 
.A(n_660),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_662),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_SL g702 ( 
.A(n_643),
.B(n_19),
.C(n_20),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_SL g703 ( 
.A1(n_640),
.A2(n_659),
.B(n_658),
.C(n_653),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_630),
.B(n_20),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_626),
.B(n_21),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_627),
.B(n_22),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_655),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_L g708 ( 
.A1(n_650),
.A2(n_22),
.B(n_23),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_656),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_636),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_617),
.A2(n_651),
.B(n_616),
.C(n_614),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_604),
.A2(n_23),
.B(n_24),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_635),
.A2(n_117),
.B(n_186),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_661),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_661),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_647),
.B(n_25),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_647),
.B(n_652),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_613),
.Y(n_719)
);

INVx3_ASAP7_75t_SL g720 ( 
.A(n_654),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_716),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_707),
.B(n_25),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_691),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_680),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_673),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_665),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_663),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_667),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_709),
.B(n_679),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_691),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_689),
.Y(n_731)
);

BUFx6f_ASAP7_75t_SL g732 ( 
.A(n_667),
.Y(n_732)
);

BUFx12f_ASAP7_75t_L g733 ( 
.A(n_688),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_667),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_26),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_690),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_701),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_714),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_676),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_700),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_697),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_714),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_714),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_692),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_715),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_715),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_671),
.B(n_678),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_671),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_706),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_677),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_666),
.B(n_27),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_715),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_683),
.Y(n_753)
);

BUFx12f_ASAP7_75t_L g754 ( 
.A(n_670),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_719),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_710),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_717),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_675),
.B(n_27),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_694),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_664),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_672),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_720),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_682),
.B(n_28),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_705),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_699),
.B(n_28),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_684),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_702),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_704),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_708),
.B(n_29),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_668),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_698),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_687),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_695),
.B(n_43),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_681),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_708),
.B(n_29),
.Y(n_777)
);

INVx6_ASAP7_75t_L g778 ( 
.A(n_685),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_696),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_693),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_713),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_724),
.B(n_686),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_726),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_729),
.B(n_711),
.Y(n_784)
);

CKINVDCx12_ASAP7_75t_R g785 ( 
.A(n_766),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_770),
.A2(n_776),
.B1(n_767),
.B2(n_778),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_724),
.B(n_712),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_727),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_781),
.A2(n_703),
.B(n_48),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_739),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_737),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_721),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_740),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_761),
.B(n_44),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_770),
.A2(n_200),
.B1(n_51),
.B2(n_52),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_721),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_778),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_756),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_780),
.A2(n_56),
.B(n_59),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_780),
.A2(n_61),
.B(n_62),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_733),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_777),
.A2(n_778),
.B1(n_771),
.B2(n_774),
.Y(n_802)
);

AO21x2_ASAP7_75t_L g803 ( 
.A1(n_764),
.A2(n_729),
.B(n_756),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_761),
.B(n_63),
.Y(n_804)
);

AO32x2_ASAP7_75t_L g805 ( 
.A1(n_764),
.A2(n_64),
.A3(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_775),
.A2(n_70),
.B(n_71),
.Y(n_806)
);

AO21x2_ASAP7_75t_L g807 ( 
.A1(n_760),
.A2(n_72),
.B(n_73),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_755),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_775),
.A2(n_74),
.B(n_76),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_728),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_760),
.A2(n_77),
.B(n_78),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_736),
.B(n_79),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_748),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_759),
.Y(n_814)
);

BUFx8_ASAP7_75t_L g815 ( 
.A(n_732),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_748),
.A2(n_747),
.B(n_735),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_736),
.B(n_81),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_735),
.A2(n_83),
.B(n_85),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_747),
.A2(n_86),
.B(n_87),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_755),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_89),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_761),
.B(n_90),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_777),
.B(n_91),
.C(n_92),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_762),
.Y(n_825)
);

AO32x2_ASAP7_75t_L g826 ( 
.A1(n_743),
.A2(n_93),
.A3(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_763),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_749),
.B(n_98),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_744),
.A2(n_99),
.B(n_101),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_763),
.Y(n_830)
);

OAI21x1_ASAP7_75t_SL g831 ( 
.A1(n_758),
.A2(n_102),
.B(n_104),
.Y(n_831)
);

BUFx4_ASAP7_75t_R g832 ( 
.A(n_772),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_755),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_758),
.A2(n_105),
.B(n_106),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_763),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_L g836 ( 
.A1(n_769),
.A2(n_109),
.B1(n_115),
.B2(n_116),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_769),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.C(n_122),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_751),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_789),
.A2(n_722),
.B(n_730),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_787),
.B(n_757),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_820),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_798),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_790),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_784),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_786),
.A2(n_754),
.B1(n_751),
.B2(n_773),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_816),
.A2(n_722),
.B(n_730),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_788),
.B(n_762),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_820),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_800),
.A2(n_762),
.B(n_779),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_786),
.A2(n_753),
.B1(n_768),
.B2(n_773),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_784),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_792),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_796),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_798),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_808),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_824),
.A2(n_726),
.B(n_723),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_799),
.A2(n_741),
.B(n_779),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_803),
.B(n_825),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_837),
.A2(n_779),
.B1(n_753),
.B2(n_773),
.Y(n_860)
);

AO21x2_ASAP7_75t_L g861 ( 
.A1(n_803),
.A2(n_753),
.B(n_723),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_791),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_782),
.B(n_743),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_799),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_793),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_821),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_829),
.A2(n_723),
.B(n_732),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_838),
.A2(n_768),
.B1(n_725),
.B2(n_731),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_833),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_799),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_815),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_835),
.Y(n_872)
);

BUFx2_ASAP7_75t_SL g873 ( 
.A(n_827),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_805),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_805),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_783),
.B(n_752),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_826),
.B(n_752),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_838),
.A2(n_745),
.B1(n_750),
.B2(n_746),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_826),
.B(n_752),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_805),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_805),
.Y(n_882)
);

BUFx2_ASAP7_75t_R g883 ( 
.A(n_801),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_810),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_845),
.B(n_802),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_R g886 ( 
.A(n_878),
.B(n_832),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_845),
.B(n_802),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_871),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_R g889 ( 
.A(n_878),
.B(n_832),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_872),
.B(n_830),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_871),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_872),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_865),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_842),
.B(n_782),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_869),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_846),
.A2(n_795),
.B1(n_837),
.B2(n_797),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_871),
.B(n_815),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_883),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_872),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_SL g900 ( 
.A1(n_840),
.A2(n_830),
.B1(n_827),
.B2(n_873),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_845),
.B(n_812),
.Y(n_901)
);

AO32x2_ASAP7_75t_L g902 ( 
.A1(n_841),
.A2(n_826),
.A3(n_785),
.B1(n_818),
.B2(n_831),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_843),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_842),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_843),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_843),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_844),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_877),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_844),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_849),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_855),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_852),
.B(n_812),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_884),
.Y(n_914)
);

NOR2x1_ASAP7_75t_L g915 ( 
.A(n_861),
.B(n_807),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_895),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_901),
.B(n_852),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_SL g918 ( 
.A1(n_900),
.A2(n_857),
.B1(n_881),
.B2(n_875),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_911),
.B(n_859),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_911),
.B(n_859),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_904),
.B(n_892),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_908),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_890),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_915),
.B(n_858),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_904),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_910),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_903),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_906),
.B(n_874),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_903),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_912),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_894),
.Y(n_931)
);

OAI221xp5_ASAP7_75t_L g932 ( 
.A1(n_896),
.A2(n_868),
.B1(n_851),
.B2(n_795),
.C(n_857),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_905),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_906),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_913),
.B(n_852),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_905),
.B(n_855),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_896),
.A2(n_822),
.B(n_881),
.C(n_875),
.Y(n_937)
);

OA21x2_ASAP7_75t_L g938 ( 
.A1(n_937),
.A2(n_870),
.B(n_864),
.Y(n_938)
);

AOI221x1_ASAP7_75t_L g939 ( 
.A1(n_937),
.A2(n_882),
.B1(n_874),
.B2(n_869),
.C(n_856),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_924),
.A2(n_870),
.B(n_864),
.Y(n_940)
);

INVx3_ASAP7_75t_SL g941 ( 
.A(n_934),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_932),
.A2(n_860),
.B(n_885),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_924),
.A2(n_870),
.B(n_864),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_925),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_931),
.B(n_909),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_922),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_918),
.B(n_887),
.C(n_822),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_921),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_927),
.A2(n_882),
.B(n_847),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_927),
.A2(n_858),
.B(n_847),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_921),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_929),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_929),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_948),
.B(n_891),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_948),
.B(n_923),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_951),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_947),
.A2(n_863),
.B1(n_888),
.B2(n_879),
.Y(n_957)
);

AOI221xp5_ASAP7_75t_L g958 ( 
.A1(n_942),
.A2(n_836),
.B1(n_930),
.B2(n_917),
.C(n_926),
.Y(n_958)
);

OAI33xp33_ASAP7_75t_L g959 ( 
.A1(n_946),
.A2(n_836),
.A3(n_916),
.B1(n_936),
.B2(n_817),
.B3(n_854),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_944),
.B(n_928),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_941),
.B(n_919),
.Y(n_961)
);

INVxp67_ASAP7_75t_SL g962 ( 
.A(n_938),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_941),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_938),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_951),
.B(n_919),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_955),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_958),
.B(n_945),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_963),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_954),
.B(n_928),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_960),
.B(n_938),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_963),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_SL g972 ( 
.A(n_957),
.B(n_898),
.C(n_893),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_954),
.B(n_891),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_968),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_966),
.B(n_956),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_965),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_973),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_969),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_972),
.B(n_961),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_972),
.B(n_897),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_967),
.B(n_938),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_974),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_976),
.B(n_970),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_977),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_952),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_959),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_897),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_975),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_978),
.B(n_962),
.Y(n_989)
);

OAI33xp33_ASAP7_75t_L g990 ( 
.A1(n_981),
.A2(n_959),
.A3(n_914),
.B1(n_964),
.B2(n_962),
.B3(n_817),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_974),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_976),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_974),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_984),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_987),
.B(n_952),
.Y(n_995)
);

NAND4xp75_ASAP7_75t_L g996 ( 
.A(n_982),
.B(n_939),
.C(n_964),
.D(n_934),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_986),
.A2(n_863),
.B1(n_818),
.B2(n_880),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_993),
.Y(n_998)
);

NOR2xp67_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_814),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_989),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_983),
.B(n_953),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_992),
.B(n_953),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_999),
.A2(n_990),
.B1(n_989),
.B2(n_988),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1000),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_994),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_985),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_1002),
.A2(n_811),
.B(n_807),
.C(n_828),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_995),
.B(n_953),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_920),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_997),
.B(n_935),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_1005),
.Y(n_1011)
);

AND3x1_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_996),
.C(n_920),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1006),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1003),
.B(n_940),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_1008),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1009),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1007),
.B(n_949),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_1005),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1011),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1019),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_940),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_943),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_943),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1016),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1012),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_1014),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1018),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1020),
.Y(n_1030)
);

NAND4xp25_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_939),
.C(n_886),
.D(n_889),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_949),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1022),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1027),
.B(n_899),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_1028),
.B(n_746),
.C(n_742),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_1026),
.B(n_834),
.C(n_794),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1034),
.B(n_1029),
.C(n_1023),
.D(n_1024),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_1030),
.A2(n_1025),
.B(n_811),
.C(n_804),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_1033),
.B(n_738),
.Y(n_1039)
);

AOI221xp5_ASAP7_75t_L g1040 ( 
.A1(n_1035),
.A2(n_794),
.B1(n_804),
.B2(n_823),
.C(n_734),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_SL g1041 ( 
.A1(n_1032),
.A2(n_873),
.B1(n_738),
.B2(n_742),
.Y(n_1041)
);

AOI211xp5_ASAP7_75t_L g1042 ( 
.A1(n_1037),
.A2(n_1036),
.B(n_1031),
.C(n_823),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_1039),
.A2(n_738),
.B(n_742),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1041),
.A2(n_950),
.B(n_899),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_1038),
.A2(n_826),
.B(n_880),
.C(n_861),
.Y(n_1045)
);

OAI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_1040),
.A2(n_746),
.B1(n_886),
.B2(n_889),
.C(n_723),
.Y(n_1046)
);

AOI211xp5_ASAP7_75t_L g1047 ( 
.A1(n_1037),
.A2(n_819),
.B(n_806),
.C(n_809),
.Y(n_1047)
);

OAI211xp5_ASAP7_75t_L g1048 ( 
.A1(n_1037),
.A2(n_866),
.B(n_949),
.C(n_856),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1037),
.A2(n_950),
.B(n_839),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1046),
.A2(n_866),
.B1(n_949),
.B2(n_856),
.Y(n_1050)
);

AOI211xp5_ASAP7_75t_L g1051 ( 
.A1(n_1043),
.A2(n_867),
.B(n_839),
.C(n_936),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_867),
.C(n_856),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1049),
.A2(n_906),
.B1(n_933),
.B2(n_863),
.Y(n_1053)
);

NOR2x1_ASAP7_75t_L g1054 ( 
.A(n_1048),
.B(n_861),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_1045),
.B(n_861),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1044),
.B(n_933),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_128),
.Y(n_1058)
);

NOR2x1p5_ASAP7_75t_L g1059 ( 
.A(n_1057),
.B(n_849),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_1058),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_L g1061 ( 
.A(n_1053),
.B(n_850),
.C(n_130),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1052),
.B(n_906),
.Y(n_1062)
);

NOR4xp75_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_841),
.C(n_134),
.D(n_135),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1054),
.B(n_876),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1056),
.A2(n_1050),
.B(n_1051),
.C(n_863),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1058),
.B(n_129),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1056),
.B(n_862),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_L g1068 ( 
.A(n_1058),
.B(n_138),
.Y(n_1068)
);

AND2x2_ASAP7_75t_SL g1069 ( 
.A(n_1058),
.B(n_848),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_1058),
.B(n_139),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1057),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1066),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1065),
.A2(n_862),
.B1(n_854),
.B2(n_876),
.C(n_848),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_1060),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1069),
.Y(n_1076)
);

XOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1070),
.B(n_1067),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_1060),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_876),
.Y(n_1079)
);

AOI221xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1064),
.A2(n_907),
.B1(n_902),
.B2(n_853),
.C(n_147),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1078),
.B(n_1059),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1076),
.B(n_1063),
.Y(n_1082)
);

AO22x2_ASAP7_75t_L g1083 ( 
.A1(n_1072),
.A2(n_1061),
.B1(n_1062),
.B2(n_907),
.Y(n_1083)
);

AND4x1_ASAP7_75t_L g1084 ( 
.A(n_1073),
.B(n_143),
.C(n_144),
.D(n_145),
.Y(n_1084)
);

XNOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1077),
.B(n_1075),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1079),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_1082),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1085),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_1081),
.A2(n_1080),
.B(n_1074),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

XNOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1090),
.B(n_1084),
.Y(n_1091)
);

INVxp33_ASAP7_75t_L g1092 ( 
.A(n_1091),
.Y(n_1092)
);

NAND4xp25_ASAP7_75t_L g1093 ( 
.A(n_1092),
.B(n_1087),
.C(n_1086),
.D(n_1089),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1092),
.Y(n_1094)
);

AOI222xp33_ASAP7_75t_L g1095 ( 
.A1(n_1094),
.A2(n_1083),
.B1(n_149),
.B2(n_150),
.C1(n_152),
.C2(n_153),
.Y(n_1095)
);

OAI222xp33_ASAP7_75t_L g1096 ( 
.A1(n_1093),
.A2(n_863),
.B1(n_154),
.B2(n_155),
.C1(n_157),
.C2(n_160),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1095),
.A2(n_1096),
.B1(n_165),
.B2(n_167),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1095),
.A2(n_148),
.B1(n_168),
.B2(n_170),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1098),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_172),
.B(n_173),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_174),
.B(n_176),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_1100),
.B1(n_177),
.B2(n_179),
.Y(n_1102)
);


endmodule