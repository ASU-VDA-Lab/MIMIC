module fake_jpeg_10094_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_4),
.Y(n_91)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_0),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_1),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_3),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_83),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_57),
.B1(n_59),
.B2(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_54),
.B1(n_51),
.B2(n_46),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_61),
.B1(n_43),
.B2(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_4),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_91),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_95),
.Y(n_102)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_5),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_28),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_42),
.B(n_32),
.C(n_33),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_29),
.C(n_34),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_98),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_115),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_100),
.B(n_111),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_100),
.B(n_110),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_102),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_96),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_104),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_108),
.B(n_106),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_122),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_107),
.B(n_105),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_109),
.Y(n_126)
);


endmodule