module fake_ariane_956_n_2084 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2084);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2084;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_1083;
wire n_337;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_62),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_144),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_73),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_136),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_7),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_108),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_63),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_31),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_84),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_72),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_118),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_62),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_181),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_2),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_82),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_92),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_77),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_170),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_99),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_23),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_142),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_81),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_121),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_93),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_109),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_70),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_106),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_71),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_122),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_63),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_107),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_70),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_95),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_18),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_149),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_172),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_163),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_12),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_169),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_133),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_69),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_151),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_120),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_152),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_17),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_45),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_161),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_51),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_153),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_143),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_195),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_115),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_148),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_43),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_66),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_60),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_102),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_180),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_87),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_123),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_54),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_188),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_89),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_57),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_5),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_124),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_71),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_178),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_141),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_74),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_139),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_52),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_129),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_34),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_19),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_67),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_79),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_11),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_110),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_191),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_26),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_61),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_54),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_125),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_45),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_39),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_167),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_43),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_113),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_137),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_37),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_135),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_104),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_12),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_53),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_192),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_112),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_38),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_26),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_37),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_29),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_100),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_157),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_83),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_90),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_6),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_13),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_29),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_28),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_96),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_159),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_74),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_103),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_30),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_53),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_21),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_86),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_150),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_35),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_22),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_164),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_28),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_44),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_140),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_24),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_47),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_21),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_61),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_134),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_58),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_42),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_97),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_126),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_19),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_40),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_68),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_25),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_94),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_24),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_77),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_51),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_158),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_216),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_219),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_252),
.B(n_0),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_209),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_206),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_278),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_315),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_222),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_209),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_211),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_252),
.B(n_0),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_392),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_390),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_390),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_242),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_239),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_225),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_255),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_197),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_255),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_372),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_222),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_260),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_260),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_224),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_226),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_266),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_235),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_266),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_244),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_247),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_222),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_348),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_298),
.B(n_1),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_249),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_242),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_202),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_250),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_257),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_258),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_202),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_272),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_275),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_202),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_267),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_269),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_275),
.B(n_1),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_273),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_288),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_208),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_208),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_279),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_208),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_221),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_288),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_304),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_290),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_304),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_369),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_306),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_291),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_221),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_303),
.B(n_4),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_293),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_296),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_221),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_306),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_200),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_309),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_302),
.B(n_6),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_348),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_236),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_309),
.B(n_9),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_316),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_236),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_299),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_271),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_301),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_308),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_236),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_271),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_200),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_234),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_312),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_205),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_271),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_316),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_314),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_199),
.B(n_201),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_317),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_232),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_348),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_338),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_338),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_205),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_346),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_397),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_455),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_346),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_357),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_357),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_357),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_453),
.B(n_305),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_408),
.B(n_204),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_R g509 ( 
.A(n_485),
.B(n_203),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_351),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_455),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_473),
.B(n_325),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_479),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_473),
.B(n_351),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_398),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_404),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_416),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_399),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_410),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_410),
.B(n_354),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_479),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_479),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_393),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_412),
.B(n_198),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_413),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_420),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_405),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_354),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_421),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_419),
.B(n_204),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_371),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_423),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_425),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_431),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_422),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_424),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_424),
.B(n_371),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_411),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_415),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_379),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_434),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_477),
.B(n_271),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_435),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_417),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_477),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_436),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_445),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_451),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_406),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_482),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_534),
.B(n_535),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_429),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_572),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_564),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_512),
.B(n_441),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_515),
.B(n_442),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_508),
.B(n_198),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_493),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_540),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_507),
.B(n_444),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_502),
.B(n_467),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_550),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_503),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_546),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_523),
.B(n_488),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_509),
.B(n_448),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_550),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_572),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_544),
.B(n_403),
.C(n_457),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_572),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_560),
.B(n_460),
.Y(n_598)
);

AND3x4_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_466),
.C(n_362),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_572),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_567),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_546),
.B(n_461),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_546),
.B(n_472),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_508),
.B(n_198),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_546),
.B(n_474),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_567),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_503),
.B(n_452),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_503),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_529),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_552),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_499),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_542),
.B(n_454),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_567),
.B(n_475),
.Y(n_617)
);

NAND3x1_ASAP7_75t_L g618 ( 
.A(n_510),
.B(n_395),
.C(n_459),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_499),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_567),
.B(n_430),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_503),
.A2(n_469),
.B1(n_407),
.B2(n_466),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_511),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_532),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_511),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_542),
.B(n_268),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_542),
.B(n_454),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_567),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_511),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_542),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_505),
.B(n_268),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_541),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_533),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_494),
.B(n_480),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_566),
.Y(n_641)
);

AO21x2_ASAP7_75t_L g642 ( 
.A1(n_497),
.A2(n_443),
.B(n_383),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_566),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_566),
.B(n_268),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_498),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_545),
.B(n_484),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_505),
.B(n_456),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_498),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_500),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_505),
.B(n_464),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_533),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_514),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_505),
.B(n_456),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_514),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_514),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_537),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_553),
.B(n_563),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_500),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_533),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_501),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_504),
.B(n_463),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_513),
.B(n_463),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_533),
.Y(n_664)
);

INVx6_ASAP7_75t_L g665 ( 
.A(n_533),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_504),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_497),
.A2(n_437),
.B1(n_440),
.B2(n_433),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_519),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_506),
.B(n_465),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_513),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_516),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_518),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_516),
.B(n_486),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_517),
.B(n_478),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_547),
.B(n_446),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_517),
.B(n_491),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_519),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_532),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_465),
.Y(n_682)
);

INVx8_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_470),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_470),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

INVx4_ASAP7_75t_SL g687 ( 
.A(n_533),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_538),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_548),
.B(n_447),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_548),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_521),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_549),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_549),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_496),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_529),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_558),
.B(n_449),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_555),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_521),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_520),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_556),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_520),
.B(n_483),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_556),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_562),
.A2(n_215),
.B1(n_323),
.B2(n_324),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_557),
.B(n_483),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_565),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_557),
.B(n_489),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_559),
.B(n_450),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_570),
.B(n_462),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_570),
.B(n_468),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_559),
.B(n_561),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_521),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_522),
.Y(n_717)
);

INVx4_ASAP7_75t_SL g718 ( 
.A(n_529),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_568),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_568),
.B(n_489),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_524),
.B(n_394),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_569),
.B(n_490),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_527),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_569),
.B(n_471),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_571),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_606),
.B(n_571),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_606),
.B(n_476),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_583),
.B(n_510),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_606),
.B(n_526),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_610),
.B(n_613),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_573),
.B(n_526),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_585),
.A2(n_554),
.B(n_551),
.C(n_543),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_672),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_579),
.B(n_539),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_683),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_637),
.A2(n_554),
.B1(n_551),
.B2(n_543),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_585),
.A2(n_539),
.B(n_530),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_637),
.A2(n_342),
.B1(n_379),
.B2(n_383),
.Y(n_738)
);

O2A1O1Ixp5_ASAP7_75t_L g739 ( 
.A1(n_585),
.A2(n_595),
.B(n_586),
.C(n_682),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_663),
.B(n_490),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_672),
.B(n_492),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_663),
.B(n_492),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_578),
.B(n_319),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_586),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_640),
.B(n_245),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_587),
.A2(n_204),
.B(n_356),
.C(n_366),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_628),
.B(n_329),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_586),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_637),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_720),
.B(n_339),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_599),
.A2(n_361),
.B1(n_276),
.B2(n_327),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_725),
.B(n_388),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_725),
.B(n_388),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_680),
.B(n_330),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_599),
.A2(n_276),
.B1(n_327),
.B2(n_361),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_725),
.B(n_241),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_218),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_720),
.B(n_353),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_720),
.B(n_367),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_691),
.B(n_331),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_682),
.B(n_356),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_682),
.B(n_356),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_703),
.B(n_218),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_287),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_599),
.A2(n_327),
.B1(n_361),
.B2(n_276),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_618),
.A2(n_366),
.B1(n_391),
.B2(n_334),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_682),
.B(n_366),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_708),
.B(n_302),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_711),
.B(n_598),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_708),
.B(n_362),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_638),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_621),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_708),
.B(n_228),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_595),
.B(n_241),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_610),
.A2(n_276),
.B1(n_361),
.B2(n_327),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_656),
.B(n_333),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_595),
.B(n_285),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_708),
.B(n_228),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_610),
.A2(n_259),
.B1(n_385),
.B2(n_369),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_643),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_656),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_643),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_639),
.B(n_285),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_639),
.B(n_360),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_591),
.B(n_336),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_683),
.Y(n_788)
);

BUFx5_ASAP7_75t_L g789 ( 
.A(n_580),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_618),
.A2(n_246),
.B1(n_277),
.B2(n_274),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_688),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_610),
.A2(n_620),
.B1(n_617),
.B2(n_676),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_688),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_588),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_645),
.A2(n_240),
.B(n_263),
.C(n_387),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_584),
.B(n_240),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_589),
.B(n_264),
.C(n_263),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_588),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_639),
.B(n_360),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_584),
.B(n_264),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_651),
.B(n_360),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_590),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_651),
.B(n_210),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_699),
.B(n_270),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_651),
.B(n_210),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_SL g806 ( 
.A1(n_612),
.A2(n_359),
.B1(n_344),
.B2(n_347),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_593),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_659),
.B(n_212),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_582),
.B(n_270),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_699),
.B(n_280),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_686),
.B(n_259),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_590),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_576),
.A2(n_530),
.B(n_527),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_700),
.B(n_280),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_576),
.A2(n_530),
.B(n_527),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_659),
.B(n_212),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_582),
.B(n_355),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_659),
.B(n_664),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_683),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_724),
.B(n_358),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_575),
.B(n_281),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_580),
.A2(n_259),
.B1(n_385),
.B2(n_369),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_589),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_676),
.B(n_281),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_676),
.B(n_284),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_705),
.A2(n_320),
.B1(n_386),
.B2(n_284),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_289),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_SL g829 ( 
.A1(n_577),
.A2(n_365),
.B1(n_364),
.B2(n_370),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_601),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_603),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_657),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_678),
.B(n_289),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_678),
.B(n_311),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_592),
.B(n_376),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_686),
.B(n_259),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_678),
.B(n_311),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_625),
.A2(n_373),
.B1(n_386),
.B2(n_322),
.C(n_384),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_580),
.A2(n_385),
.B1(n_369),
.B2(n_287),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_645),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_603),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_664),
.B(n_231),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_581),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_596),
.B(n_646),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_709),
.B(n_387),
.C(n_384),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_L g846 ( 
.A1(n_705),
.A2(n_350),
.B1(n_381),
.B2(n_340),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_664),
.B(n_671),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_678),
.B(n_320),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_709),
.B(n_696),
.Y(n_849)
);

AND2x6_ASAP7_75t_L g850 ( 
.A(n_648),
.B(n_231),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_671),
.B(n_328),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_671),
.B(n_648),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_608),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_613),
.B(n_287),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_696),
.B(n_604),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_581),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_657),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_601),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_608),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_721),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_684),
.B(n_322),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_660),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_684),
.B(n_326),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_661),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_614),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_605),
.B(n_378),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_661),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_635),
.A2(n_326),
.B1(n_381),
.B2(n_349),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_685),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_607),
.B(n_380),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_635),
.B(n_340),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_666),
.Y(n_873)
);

INVx8_ASAP7_75t_L g874 ( 
.A(n_580),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_614),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_666),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_685),
.B(n_343),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_674),
.B(n_207),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_635),
.B(n_343),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_SL g880 ( 
.A(n_674),
.B(n_368),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_633),
.B(n_349),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_714),
.B(n_350),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_650),
.B(n_373),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_650),
.B(n_375),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_616),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_650),
.B(n_375),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_580),
.B(n_374),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_620),
.A2(n_286),
.B1(n_382),
.B2(n_214),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_673),
.Y(n_889)
);

AND2x6_ASAP7_75t_SL g890 ( 
.A(n_717),
.B(n_377),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_648),
.B(n_658),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_714),
.B(n_377),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_717),
.B(n_633),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_616),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_658),
.B(n_668),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_783),
.B(n_650),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_730),
.B(n_615),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_728),
.B(n_615),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_730),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_840),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_734),
.B(n_631),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_731),
.B(n_631),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_769),
.A2(n_574),
.B1(n_620),
.B2(n_677),
.Y(n_903)
);

NAND2x1p5_ASAP7_75t_L g904 ( 
.A(n_820),
.B(n_658),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_874),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_743),
.B(n_668),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_730),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_861),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_745),
.B(n_668),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_735),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_863),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_760),
.B(n_749),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_849),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_783),
.B(n_698),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_870),
.B(n_673),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_729),
.A2(n_593),
.B1(n_594),
.B2(n_719),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_733),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_865),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_794),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_794),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_740),
.B(n_681),
.Y(n_921)
);

CKINVDCx6p67_ASAP7_75t_R g922 ( 
.A(n_824),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_742),
.B(n_681),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_868),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_874),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_792),
.A2(n_620),
.B1(n_630),
.B2(n_580),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_820),
.B(n_735),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_820),
.B(n_735),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_843),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_843),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_787),
.B(n_609),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_SL g932 ( 
.A(n_856),
.B(n_577),
.C(n_707),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_874),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_798),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_738),
.A2(n_580),
.B1(n_630),
.B2(n_713),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_798),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_880),
.B(n_594),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_733),
.B(n_712),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_873),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_856),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_752),
.A2(n_630),
.B1(n_647),
.B2(n_653),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_832),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_752),
.A2(n_753),
.B1(n_844),
.B2(n_818),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_889),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_802),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_SL g947 ( 
.A(n_777),
.B(n_667),
.C(n_662),
.Y(n_947)
);

NOR3xp33_ASAP7_75t_SL g948 ( 
.A(n_829),
.B(n_806),
.C(n_827),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_771),
.Y(n_949)
);

OR2x2_ASAP7_75t_SL g950 ( 
.A(n_727),
.B(n_665),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_772),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_773),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_874),
.B(n_690),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_741),
.B(n_670),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_846),
.B(n_722),
.C(n_710),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_860),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_771),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_793),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_779),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_753),
.A2(n_726),
.B1(n_755),
.B2(n_751),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_811),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_893),
.B(n_690),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_813),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_736),
.A2(n_695),
.B1(n_719),
.B2(n_716),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_883),
.B(n_692),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_788),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_813),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_747),
.B(n_597),
.Y(n_970)
);

INVx6_ASAP7_75t_L g971 ( 
.A(n_820),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_872),
.B(n_630),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_809),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_744),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_812),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_779),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_782),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_879),
.B(n_750),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_754),
.B(n_855),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_830),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_857),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_836),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_820),
.B(n_687),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_789),
.B(n_692),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_782),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_830),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_858),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_757),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_788),
.B(n_687),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_887),
.B(n_630),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_881),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_788),
.B(n_683),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_758),
.B(n_630),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_858),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_765),
.A2(n_630),
.B1(n_716),
.B2(n_706),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_821),
.B(n_597),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_887),
.B(n_683),
.Y(n_997)
);

CKINVDCx6p67_ASAP7_75t_R g998 ( 
.A(n_850),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_866),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_866),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_784),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_884),
.B(n_694),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_850),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_881),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_875),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_881),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_784),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_744),
.A2(n_695),
.B1(n_706),
.B2(n_704),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_838),
.A2(n_642),
.B1(n_665),
.B2(n_641),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_831),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_789),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_850),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_759),
.B(n_694),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_875),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_763),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_L g1016 ( 
.A(n_850),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_831),
.B(n_687),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_885),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_775),
.A2(n_622),
.B(n_602),
.Y(n_1019)
);

AND3x1_ASAP7_75t_SL g1020 ( 
.A(n_890),
.B(n_704),
.C(n_600),
.Y(n_1020)
);

AO22x1_ASAP7_75t_L g1021 ( 
.A1(n_850),
.A2(n_644),
.B1(n_622),
.B2(n_641),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_885),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_770),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_886),
.B(n_796),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_R g1025 ( 
.A(n_867),
.B(n_624),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_894),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_841),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_894),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_766),
.A2(n_600),
.B(n_624),
.C(n_602),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_800),
.B(n_642),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_789),
.B(n_624),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_744),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_804),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_822),
.B(n_642),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_789),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_825),
.B(n_623),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_826),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_828),
.B(n_623),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_841),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_850),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_871),
.B(n_229),
.C(n_213),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_891),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_891),
.Y(n_1043)
);

BUFx4_ASAP7_75t_SL g1044 ( 
.A(n_853),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_761),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_853),
.B(n_687),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_833),
.B(n_627),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_789),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_835),
.B(n_665),
.Y(n_1049)
);

AND2x6_ASAP7_75t_L g1050 ( 
.A(n_748),
.B(n_627),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_882),
.B(n_619),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_892),
.B(n_227),
.C(n_363),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_869),
.B(n_223),
.C(n_352),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_834),
.B(n_665),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_810),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_859),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_815),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_762),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_895),
.Y(n_1059)
);

AO22x1_ASAP7_75t_L g1060 ( 
.A1(n_797),
.A2(n_644),
.B1(n_328),
.B2(n_368),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_756),
.B(n_790),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_748),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_859),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_767),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_862),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_776),
.A2(n_619),
.B1(n_626),
.B2(n_629),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_895),
.Y(n_1067)
);

BUFx4f_ASAP7_75t_SL g1068 ( 
.A(n_756),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_807),
.B(n_718),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_837),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_848),
.B(n_626),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_789),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_789),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_748),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_774),
.B(n_629),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_739),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_764),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_780),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_888),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_864),
.B(n_634),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_877),
.Y(n_1081)
);

INVx6_ASAP7_75t_L g1082 ( 
.A(n_852),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_732),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_819),
.B(n_718),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_819),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_768),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_845),
.B(n_634),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_979),
.B(n_878),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1019),
.A2(n_814),
.B(n_816),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1019),
.A2(n_737),
.B(n_746),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_905),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_912),
.A2(n_775),
.B(n_778),
.C(n_785),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_898),
.B(n_901),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_988),
.B(n_795),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_942),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_922),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_902),
.B(n_781),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1076),
.A2(n_854),
.B(n_764),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1081),
.B(n_854),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_1034),
.A2(n_778),
.B(n_795),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_852),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1030),
.A2(n_785),
.B(n_851),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_913),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_897),
.B(n_907),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_906),
.B(n_611),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_931),
.A2(n_786),
.B(n_799),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_922),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1083),
.A2(n_851),
.B(n_805),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1015),
.B(n_652),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1083),
.A2(n_817),
.B(n_842),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_996),
.A2(n_847),
.B(n_801),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_929),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_970),
.A2(n_909),
.B(n_966),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_972),
.A2(n_847),
.B(n_801),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1024),
.B(n_823),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1076),
.A2(n_842),
.B(n_817),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1037),
.B(n_839),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1072),
.A2(n_808),
.B(n_805),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1072),
.A2(n_808),
.B(n_803),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_899),
.B(n_786),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1008),
.A2(n_803),
.B(n_799),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_1061),
.A2(n_723),
.B(n_715),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1065),
.B(n_652),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_974),
.A2(n_636),
.B(n_611),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_967),
.B(n_654),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1044),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_SL g1127 ( 
.A1(n_1042),
.A2(n_723),
.B(n_654),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_967),
.B(n_1002),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_SL g1129 ( 
.A1(n_927),
.A2(n_679),
.B(n_715),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_956),
.A2(n_903),
.B(n_978),
.C(n_923),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_984),
.A2(n_655),
.B(n_669),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_904),
.A2(n_655),
.B(n_669),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_900),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_991),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_611),
.B(n_702),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_916),
.A2(n_679),
.B(n_701),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_904),
.A2(n_693),
.B(n_689),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1002),
.B(n_689),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_904),
.A2(n_693),
.B(n_701),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1042),
.A2(n_1067),
.A3(n_1059),
.B(n_920),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_913),
.B(n_644),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_921),
.A2(n_611),
.B(n_702),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_910),
.A2(n_718),
.B(n_702),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1021),
.A2(n_718),
.B(n_702),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_910),
.A2(n_702),
.B(n_697),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_955),
.B(n_644),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1059),
.A2(n_644),
.A3(n_368),
.B(n_374),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_910),
.A2(n_697),
.B(n_636),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_908),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1029),
.A2(n_644),
.B(n_697),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_948),
.A2(n_369),
.B(n_385),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_911),
.Y(n_1152)
);

NAND2x1_ASAP7_75t_L g1153 ( 
.A(n_971),
.B(n_611),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_968),
.A2(n_644),
.B(n_697),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_929),
.B(n_217),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1079),
.A2(n_294),
.B1(n_230),
.B2(n_233),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1067),
.A2(n_374),
.A3(n_636),
.B(n_632),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_968),
.A2(n_697),
.B(n_636),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1085),
.B(n_632),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_968),
.A2(n_636),
.B(n_632),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_L g1161 ( 
.A(n_1050),
.B(n_632),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_919),
.A2(n_374),
.A3(n_632),
.B(n_234),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_930),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1075),
.A2(n_374),
.B(n_234),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_919),
.A2(n_374),
.A3(n_234),
.B(n_369),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_963),
.B(n_385),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_955),
.B(n_9),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_921),
.B(n_10),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_923),
.B(n_10),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_962),
.A2(n_385),
.B(n_13),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_920),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1074),
.A2(n_253),
.B(n_345),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1074),
.A2(n_251),
.B(n_341),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1074),
.A2(n_248),
.B(n_337),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1078),
.B(n_11),
.Y(n_1175)
);

OAI22x1_ASAP7_75t_L g1176 ( 
.A1(n_935),
.A2(n_942),
.B1(n_973),
.B2(n_938),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_918),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_SL g1178 ( 
.A1(n_940),
.A2(n_947),
.B(n_926),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_949),
.A2(n_960),
.B(n_958),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_930),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_907),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_949),
.A2(n_374),
.B(n_234),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_924),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_958),
.A2(n_374),
.B(n_234),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_960),
.A2(n_374),
.B(n_80),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1070),
.B(n_14),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_976),
.A2(n_88),
.B(n_101),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_897),
.B(n_14),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_976),
.A2(n_335),
.B(n_332),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1043),
.A2(n_321),
.B(n_318),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1017),
.B(n_116),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_934),
.A2(n_994),
.A3(n_999),
.B(n_936),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1013),
.A2(n_313),
.B(n_310),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_897),
.B(n_15),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_977),
.A2(n_119),
.B(n_130),
.Y(n_1195)
);

BUFx2_ASAP7_75t_SL g1196 ( 
.A(n_957),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_995),
.A2(n_945),
.B1(n_939),
.B2(n_943),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1004),
.B(n_15),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1051),
.A2(n_964),
.B(n_1016),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1016),
.A2(n_307),
.B(n_300),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1006),
.B(n_16),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1010),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_940),
.B(n_17),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1016),
.A2(n_297),
.B(n_295),
.Y(n_1204)
);

NAND2x1_ASAP7_75t_L g1205 ( 
.A(n_971),
.B(n_196),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1053),
.B(n_292),
.C(n_283),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_934),
.A2(n_965),
.A3(n_936),
.B(n_946),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_927),
.A2(n_282),
.B(n_265),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_915),
.B(n_20),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1043),
.A2(n_941),
.B(n_1080),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1017),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1085),
.B(n_262),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_915),
.B(n_20),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_924),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1033),
.B(n_22),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_917),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_SL g1217 ( 
.A1(n_1063),
.A2(n_943),
.B(n_939),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1080),
.A2(n_261),
.B(n_256),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_957),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_982),
.B(n_25),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_981),
.B(n_27),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1055),
.B(n_27),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_945),
.A2(n_254),
.B1(n_243),
.B2(n_238),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1057),
.A2(n_237),
.B(n_220),
.C(n_32),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_977),
.A2(n_179),
.B(n_177),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1063),
.A2(n_30),
.B(n_31),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1087),
.A2(n_32),
.B(n_33),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1079),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1082),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1023),
.B(n_41),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_905),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1007),
.A2(n_176),
.B(n_173),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_927),
.A2(n_171),
.B(n_165),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1007),
.A2(n_146),
.B(n_131),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1036),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_928),
.A2(n_50),
.B(n_52),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1022),
.A2(n_55),
.B(n_56),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1021),
.A2(n_55),
.B(n_56),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_993),
.A2(n_1022),
.B(n_1028),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1082),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1028),
.A2(n_59),
.B(n_60),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_928),
.A2(n_64),
.B(n_65),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_946),
.A2(n_64),
.B(n_65),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_961),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1025),
.A2(n_66),
.B(n_67),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1086),
.B(n_68),
.Y(n_1246)
);

NAND2x1_ASAP7_75t_L g1247 ( 
.A(n_971),
.B(n_69),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1048),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1036),
.A2(n_72),
.B(n_73),
.Y(n_1249)
);

AND2x6_ASAP7_75t_L g1250 ( 
.A(n_905),
.B(n_75),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1045),
.B(n_75),
.Y(n_1251)
);

BUFx2_ASAP7_75t_R g1252 ( 
.A(n_1107),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1164),
.A2(n_1105),
.B(n_1210),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1202),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1091),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1164),
.A2(n_1001),
.B(n_985),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1202),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1211),
.B(n_1010),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1126),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1184),
.A2(n_1005),
.B(n_1026),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1133),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_914),
.B(n_896),
.C(n_937),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1184),
.A2(n_980),
.B(n_1014),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1088),
.B(n_981),
.Y(n_1264)
);

AOI221xp5_ASAP7_75t_L g1265 ( 
.A1(n_1170),
.A2(n_932),
.B1(n_973),
.B2(n_1041),
.C(n_1060),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1094),
.A2(n_1068),
.B1(n_1064),
.B2(n_1058),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1192),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1211),
.B(n_1056),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1093),
.B(n_1038),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1149),
.Y(n_1270)
);

CKINVDCx6p67_ASAP7_75t_R g1271 ( 
.A(n_1096),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1095),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1182),
.A2(n_1089),
.B(n_1090),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1090),
.A2(n_986),
.B(n_1018),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1150),
.A2(n_1018),
.B(n_986),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1192),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1161),
.A2(n_1048),
.B(n_1073),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1150),
.A2(n_980),
.B(n_1026),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1185),
.A2(n_1014),
.B(n_987),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1152),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1185),
.A2(n_1005),
.B(n_965),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1104),
.B(n_1027),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1104),
.B(n_1027),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1103),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1158),
.A2(n_999),
.B(n_969),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1177),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1151),
.A2(n_1038),
.B1(n_1047),
.B2(n_1054),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1103),
.B(n_1056),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1128),
.B(n_950),
.Y(n_1289)
);

AOI22x1_ASAP7_75t_L g1290 ( 
.A1(n_1113),
.A2(n_1062),
.B1(n_1032),
.B2(n_1039),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1104),
.B(n_1039),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1181),
.B(n_950),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1096),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1216),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1134),
.B(n_1047),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1183),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1107),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1101),
.B(n_1085),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1130),
.B(n_1071),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1180),
.B(n_1046),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1112),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1105),
.A2(n_961),
.B(n_994),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1214),
.B(n_1071),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1134),
.B(n_951),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1101),
.A2(n_1050),
.B(n_1054),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1181),
.B(n_1017),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1122),
.A2(n_990),
.B(n_1000),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1092),
.A2(n_1050),
.B(n_1009),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1167),
.B(n_1168),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1158),
.A2(n_1000),
.B(n_969),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1192),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1141),
.B(n_1046),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1109),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1102),
.A2(n_1060),
.B(n_1012),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1171),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1249),
.A2(n_1077),
.B(n_1012),
.C(n_975),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1219),
.B(n_1046),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1091),
.B(n_1039),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1160),
.A2(n_987),
.B(n_1077),
.Y(n_1319)
);

NOR2x1_ASAP7_75t_L g1320 ( 
.A(n_1112),
.B(n_954),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1156),
.B(n_959),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1169),
.B(n_952),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1160),
.A2(n_1077),
.B(n_1062),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1228),
.A2(n_998),
.B1(n_1003),
.B2(n_1040),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1207),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1163),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1248),
.A2(n_1082),
.B1(n_998),
.B2(n_1039),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1116),
.A2(n_1066),
.B(n_1052),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1161),
.A2(n_1073),
.B(n_1011),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1246),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1163),
.B(n_1039),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1091),
.Y(n_1332)
);

AO21x1_ASAP7_75t_L g1333 ( 
.A1(n_1197),
.A2(n_1011),
.B(n_1035),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1091),
.B(n_1069),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1196),
.B(n_1069),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1098),
.A2(n_1032),
.B(n_1062),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1231),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1191),
.B(n_905),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1231),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1221),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1203),
.B(n_1082),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1207),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1178),
.B(n_1032),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1116),
.A2(n_1084),
.B(n_1069),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1207),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1145),
.A2(n_1011),
.B(n_1035),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_1035),
.B(n_1050),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1154),
.A2(n_1050),
.B(n_1003),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1231),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1144),
.A2(n_1084),
.B(n_928),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1231),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1176),
.A2(n_953),
.B1(n_1049),
.B2(n_1085),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1154),
.A2(n_1050),
.B(n_1003),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1218),
.A2(n_953),
.B1(n_1085),
.B2(n_1003),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1108),
.A2(n_1003),
.B(n_1040),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1108),
.A2(n_1040),
.B(n_953),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1110),
.A2(n_1040),
.B(n_953),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1111),
.A2(n_953),
.B(n_1084),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1110),
.A2(n_1040),
.B(n_953),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1220),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1120),
.A2(n_1020),
.B1(n_933),
.B2(n_905),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1250),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1248),
.A2(n_992),
.B1(n_925),
.B2(n_933),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1209),
.B(n_925),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1171),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1244),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1195),
.A2(n_971),
.B(n_992),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1244),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1140),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1136),
.A2(n_983),
.B(n_989),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1140),
.Y(n_1371)
);

AND2x6_ASAP7_75t_L g1372 ( 
.A(n_1120),
.B(n_925),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1140),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1250),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1166),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1140),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1245),
.A2(n_997),
.B1(n_925),
.B2(n_933),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1213),
.A2(n_1224),
.B1(n_1188),
.B2(n_1194),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1239),
.A2(n_1217),
.B(n_1106),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1186),
.B(n_76),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1198),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1153),
.B(n_925),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1191),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1238),
.A2(n_992),
.B(n_933),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1215),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1224),
.A2(n_992),
.B(n_989),
.C(n_983),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1235),
.A2(n_1247),
.B(n_1205),
.C(n_1159),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1097),
.A2(n_933),
.B1(n_989),
.B2(n_983),
.Y(n_1388)
);

AOI222xp33_ASAP7_75t_L g1389 ( 
.A1(n_1235),
.A2(n_78),
.B1(n_1240),
.B2(n_1229),
.C1(n_1175),
.C2(n_1222),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1146),
.A2(n_78),
.B1(n_1190),
.B2(n_1099),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1207),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1195),
.A2(n_1225),
.B(n_1132),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1239),
.A2(n_1114),
.B(n_1159),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1230),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1225),
.A2(n_1132),
.B(n_1131),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1179),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1250),
.A2(n_1115),
.B1(n_1189),
.B2(n_1117),
.Y(n_1397)
);

AOI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1251),
.A2(n_1223),
.B1(n_1201),
.B2(n_1206),
.C(n_1138),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1179),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1212),
.Y(n_1400)
);

AOI221xp5_ASAP7_75t_L g1401 ( 
.A1(n_1125),
.A2(n_1242),
.B1(n_1236),
.B2(n_1193),
.C(n_1226),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1123),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1131),
.A2(n_1227),
.B(n_1118),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1237),
.A2(n_1241),
.B(n_1121),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1155),
.B(n_1212),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1127),
.Y(n_1406)
);

AOI222xp33_ASAP7_75t_L g1407 ( 
.A1(n_1250),
.A2(n_1241),
.B1(n_1237),
.B2(n_1121),
.C1(n_1119),
.C2(n_1118),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1119),
.A2(n_1143),
.B(n_1234),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1187),
.A2(n_1232),
.B(n_1142),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1124),
.A2(n_1139),
.B(n_1137),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1189),
.A2(n_1100),
.B1(n_1250),
.B2(n_1204),
.Y(n_1411)
);

INVx4_ASAP7_75t_SL g1412 ( 
.A(n_1147),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1172),
.A2(n_1173),
.B(n_1174),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_SL g1414 ( 
.A(n_1129),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1243),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1135),
.A2(n_1199),
.B(n_1233),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1100),
.A2(n_1243),
.B(n_1208),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1243),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1165),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1162),
.A2(n_1157),
.B(n_1165),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1165),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1362),
.B(n_1100),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1389),
.A2(n_1189),
.B1(n_1200),
.B2(n_1147),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_1157),
.B1(n_1147),
.B2(n_1162),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1261),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1334),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1338),
.B(n_1157),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1257),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1267),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1257),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1326),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1360),
.B(n_1147),
.Y(n_1432)
);

AOI222xp33_ASAP7_75t_L g1433 ( 
.A1(n_1321),
.A2(n_1162),
.B1(n_1265),
.B2(n_1394),
.C1(n_1309),
.C2(n_1378),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1394),
.A2(n_1400),
.B1(n_1385),
.B2(n_1299),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1362),
.B(n_1374),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1392),
.A2(n_1409),
.B(n_1395),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1259),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1360),
.B(n_1330),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1269),
.B(n_1313),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1362),
.A2(n_1374),
.B1(n_1289),
.B2(n_1295),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1272),
.B(n_1303),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1381),
.A2(n_1289),
.B1(n_1405),
.B2(n_1304),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1264),
.A2(n_1343),
.B1(n_1266),
.B2(n_1316),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1343),
.A2(n_1316),
.B1(n_1398),
.B2(n_1340),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1271),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1270),
.Y(n_1447)
);

NOR3xp33_ASAP7_75t_SL g1448 ( 
.A(n_1293),
.B(n_1331),
.C(n_1288),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1284),
.B(n_1292),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1341),
.B(n_1301),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1341),
.B(n_1283),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1280),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1283),
.B(n_1326),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1362),
.A2(n_1374),
.B1(n_1340),
.B2(n_1375),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1286),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1362),
.B(n_1374),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1374),
.A2(n_1375),
.B1(n_1292),
.B2(n_1361),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1306),
.B(n_1322),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1306),
.B(n_1322),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1383),
.B(n_1334),
.Y(n_1460)
);

OAI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1320),
.A2(n_1401),
.B1(n_1262),
.B2(n_1390),
.C(n_1308),
.Y(n_1461)
);

NOR2xp67_ASAP7_75t_SL g1462 ( 
.A(n_1293),
.B(n_1297),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1252),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1271),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1296),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_L g1466 ( 
.A(n_1297),
.B(n_1254),
.Y(n_1466)
);

OAI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1397),
.A2(n_1407),
.B(n_1305),
.C(n_1298),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1338),
.B(n_1383),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1315),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1365),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1287),
.A2(n_1298),
.B1(n_1354),
.B2(n_1299),
.Y(n_1471)
);

AND2x2_ASAP7_75t_SL g1472 ( 
.A(n_1370),
.B(n_1418),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1324),
.A2(n_1282),
.B1(n_1294),
.B2(n_1402),
.Y(n_1473)
);

OAI222xp33_ASAP7_75t_L g1474 ( 
.A1(n_1352),
.A2(n_1303),
.B1(n_1411),
.B2(n_1366),
.C1(n_1368),
.C2(n_1338),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1337),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1312),
.B(n_1254),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1414),
.A2(n_1418),
.B1(n_1370),
.B2(n_1358),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1392),
.A2(n_1409),
.B(n_1395),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1312),
.B(n_1282),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1276),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1364),
.A2(n_1258),
.B1(n_1386),
.B2(n_1268),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1334),
.B(n_1268),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1332),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1369),
.Y(n_1485)
);

CKINVDCx16_ASAP7_75t_R g1486 ( 
.A(n_1300),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1273),
.A2(n_1403),
.B(n_1417),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1268),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1312),
.A2(n_1300),
.B1(n_1418),
.B2(n_1317),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1277),
.A2(n_1413),
.B(n_1329),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1370),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1300),
.A2(n_1418),
.B1(n_1317),
.B2(n_1328),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_1317),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1258),
.A2(n_1377),
.B1(n_1290),
.B2(n_1291),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1335),
.B(n_1332),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1328),
.A2(n_1371),
.B1(n_1373),
.B2(n_1376),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1276),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1311),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1327),
.B(n_1333),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1403),
.A2(n_1273),
.B(n_1416),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1311),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1291),
.B(n_1337),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1325),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1338),
.A2(n_1363),
.B1(n_1388),
.B2(n_1328),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1325),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1372),
.B2(n_1415),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1349),
.Y(n_1507)
);

OR2x4_ASAP7_75t_L g1508 ( 
.A(n_1349),
.B(n_1259),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1259),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1333),
.A2(n_1346),
.B(n_1387),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1372),
.B2(n_1307),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1255),
.A2(n_1339),
.B1(n_1318),
.B2(n_1351),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1349),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1274),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1372),
.A2(n_1307),
.B1(n_1420),
.B2(n_1419),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1372),
.A2(n_1307),
.B1(n_1420),
.B2(n_1421),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1351),
.B(n_1255),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1255),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1339),
.A2(n_1318),
.B1(n_1349),
.B2(n_1382),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1339),
.B(n_1372),
.Y(n_1520)
);

AOI222xp33_ASAP7_75t_L g1521 ( 
.A1(n_1372),
.A2(n_1412),
.B1(n_1399),
.B2(n_1396),
.C1(n_1384),
.C2(n_1275),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1379),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1420),
.A2(n_1344),
.B1(n_1302),
.B2(n_1274),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1387),
.A2(n_1396),
.B1(n_1399),
.B2(n_1253),
.C(n_1379),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1406),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1274),
.Y(n_1526)
);

BUFx8_ASAP7_75t_SL g1527 ( 
.A(n_1406),
.Y(n_1527)
);

BUFx10_ASAP7_75t_L g1528 ( 
.A(n_1382),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1379),
.B(n_1350),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1344),
.A2(n_1302),
.B1(n_1412),
.B2(n_1253),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1412),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1404),
.A2(n_1344),
.B1(n_1302),
.B2(n_1256),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1404),
.A2(n_1314),
.B1(n_1256),
.B2(n_1410),
.C(n_1260),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1393),
.B(n_1404),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1275),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1253),
.A2(n_1393),
.B1(n_1260),
.B2(n_1279),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1393),
.B(n_1323),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1260),
.A2(n_1256),
.B1(n_1410),
.B2(n_1348),
.Y(n_1538)
);

INVx6_ASAP7_75t_L g1539 ( 
.A(n_1323),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1279),
.A2(n_1281),
.B1(n_1278),
.B2(n_1263),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1278),
.B(n_1285),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1285),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1310),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1348),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1310),
.B(n_1336),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1263),
.Y(n_1546)
);

INVx6_ASAP7_75t_L g1547 ( 
.A(n_1319),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1353),
.A2(n_1367),
.B1(n_1356),
.B2(n_1359),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1281),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1319),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_SL g1551 ( 
.A(n_1416),
.B(n_1336),
.C(n_1408),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1408),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1353),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1356),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1367),
.B(n_1357),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1357),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1359),
.A2(n_1355),
.B1(n_1347),
.B2(n_1410),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1355),
.B(n_1347),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1346),
.A2(n_769),
.B1(n_399),
.B2(n_415),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1380),
.A2(n_944),
.B1(n_769),
.B2(n_979),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1389),
.A2(n_599),
.B1(n_769),
.B2(n_947),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1272),
.B(n_1284),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1334),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1261),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1380),
.A2(n_769),
.B1(n_979),
.B2(n_760),
.C(n_743),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1269),
.B(n_979),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1261),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1389),
.A2(n_599),
.B1(n_769),
.B2(n_947),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1269),
.B(n_979),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1261),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1257),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1261),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1389),
.A2(n_599),
.B1(n_769),
.B2(n_947),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1293),
.Y(n_1576)
);

OAI21xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1389),
.A2(n_1249),
.B(n_944),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1269),
.B(n_979),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1261),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1261),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1389),
.A2(n_599),
.B1(n_769),
.B2(n_947),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1284),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1389),
.A2(n_599),
.B1(n_769),
.B2(n_947),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1383),
.B(n_1299),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1272),
.B(n_1284),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1394),
.A2(n_769),
.B1(n_979),
.B2(n_743),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1583),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1577),
.A2(n_1560),
.B1(n_1445),
.B2(n_1444),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1561),
.A2(n_1569),
.B1(n_1575),
.B2(n_1581),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1586),
.A2(n_1566),
.B1(n_1583),
.B2(n_1569),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1461),
.A2(n_1567),
.B1(n_1570),
.B2(n_1578),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1442),
.B(n_1458),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1446),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1467),
.A2(n_1584),
.B1(n_1471),
.B2(n_1443),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1446),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1584),
.B(n_1435),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1510),
.A2(n_1490),
.B(n_1478),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1434),
.A2(n_1559),
.B1(n_1508),
.B2(n_1448),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1433),
.A2(n_1434),
.B1(n_1457),
.B2(n_1423),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1428),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1499),
.A2(n_1441),
.B(n_1456),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1584),
.A2(n_1432),
.B1(n_1472),
.B2(n_1486),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1582),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1459),
.B(n_1440),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1423),
.A2(n_1499),
.B(n_1477),
.C(n_1491),
.Y(n_1605)
);

BUFx10_ASAP7_75t_L g1606 ( 
.A(n_1508),
.Y(n_1606)
);

OAI33xp33_ASAP7_75t_L g1607 ( 
.A1(n_1449),
.A2(n_1465),
.A3(n_1447),
.B1(n_1425),
.B2(n_1574),
.B3(n_1565),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1562),
.B(n_1585),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1450),
.B(n_1451),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1475),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1500),
.A2(n_1436),
.B(n_1540),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1457),
.A2(n_1474),
.B1(n_1584),
.B2(n_1454),
.C1(n_1473),
.C2(n_1572),
.Y(n_1612)
);

INVx3_ASAP7_75t_SL g1613 ( 
.A(n_1464),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1435),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1430),
.B(n_1452),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1463),
.A2(n_1454),
.B1(n_1473),
.B2(n_1493),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1439),
.A2(n_1431),
.B1(n_1509),
.B2(n_1437),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1453),
.B(n_1476),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1438),
.B(n_1564),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1428),
.Y(n_1620)
);

BUFx12f_ASAP7_75t_L g1621 ( 
.A(n_1475),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1438),
.B(n_1564),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1424),
.A2(n_1580),
.B1(n_1568),
.B2(n_1579),
.C(n_1455),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1469),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1573),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1509),
.A2(n_1481),
.B1(n_1525),
.B2(n_1488),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1576),
.A2(n_1513),
.B1(n_1573),
.B2(n_1527),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1504),
.A2(n_1493),
.B1(n_1470),
.B2(n_1460),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1529),
.A2(n_1522),
.B(n_1494),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1571),
.B(n_1482),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1571),
.B(n_1482),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1479),
.B(n_1483),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1517),
.Y(n_1633)
);

OAI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1518),
.A2(n_1524),
.B(n_1537),
.C(n_1466),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1456),
.A2(n_1558),
.B(n_1538),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1460),
.A2(n_1527),
.B1(n_1576),
.B2(n_1485),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1484),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1497),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1489),
.A2(n_1506),
.B1(n_1520),
.B2(n_1468),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1460),
.A2(n_1492),
.B1(n_1506),
.B2(n_1427),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1480),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1489),
.A2(n_1520),
.B1(n_1468),
.B2(n_1563),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1498),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1551),
.A2(n_1552),
.B(n_1545),
.C(n_1533),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1462),
.A2(n_1468),
.B1(n_1563),
.B2(n_1426),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1529),
.A2(n_1515),
.B(n_1516),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1540),
.A2(n_1536),
.B(n_1541),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1427),
.B(n_1426),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1501),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1538),
.A2(n_1514),
.B(n_1526),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1532),
.A2(n_1534),
.B1(n_1492),
.B2(n_1537),
.C(n_1496),
.Y(n_1651)
);

OAI211xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1557),
.A2(n_1521),
.B(n_1507),
.C(n_1536),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1496),
.A2(n_1516),
.B1(n_1515),
.B2(n_1523),
.C(n_1511),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1505),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1542),
.A2(n_1543),
.B(n_1512),
.C(n_1530),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1519),
.B(n_1548),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1502),
.B(n_1495),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1549),
.A2(n_1546),
.B(n_1422),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1495),
.B(n_1472),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1422),
.A2(n_1539),
.B1(n_1427),
.B2(n_1511),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1554),
.B(n_1544),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1531),
.A2(n_1514),
.B1(n_1503),
.B2(n_1530),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1531),
.A2(n_1556),
.B1(n_1523),
.B2(n_1547),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1555),
.A2(n_1554),
.B(n_1549),
.C(n_1550),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1546),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1531),
.A2(n_1556),
.B1(n_1547),
.B2(n_1539),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1528),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1547),
.A2(n_1539),
.B1(n_1550),
.B2(n_1535),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1553),
.A2(n_1544),
.B1(n_1535),
.B2(n_1487),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1528),
.A2(n_1569),
.B1(n_1575),
.B2(n_1561),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1487),
.B(n_1458),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1429),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1577),
.A2(n_1560),
.B1(n_1445),
.B2(n_769),
.Y(n_1674)
);

OAI21xp33_ASAP7_75t_L g1675 ( 
.A1(n_1566),
.A2(n_1586),
.B(n_1560),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_SL g1676 ( 
.A(n_1509),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1566),
.A2(n_1560),
.B1(n_769),
.B2(n_979),
.C(n_743),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1577),
.A2(n_1560),
.B1(n_1445),
.B2(n_769),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1428),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1446),
.Y(n_1681)
);

OAI211xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1586),
.A2(n_1566),
.B(n_583),
.C(n_574),
.Y(n_1682)
);

CKINVDCx11_ASAP7_75t_R g1683 ( 
.A(n_1446),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1428),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1586),
.A2(n_1566),
.B1(n_1560),
.B2(n_1561),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1566),
.A2(n_1560),
.B1(n_769),
.B2(n_979),
.C(n_743),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1566),
.B(n_1586),
.C(n_1560),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1429),
.Y(n_1689)
);

OAI322xp33_ASAP7_75t_L g1690 ( 
.A1(n_1560),
.A2(n_1586),
.A3(n_219),
.B1(n_1228),
.B2(n_403),
.C1(n_769),
.C2(n_390),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1509),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1566),
.A2(n_769),
.B1(n_1586),
.B2(n_1560),
.C(n_1569),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1586),
.A2(n_1566),
.B1(n_1560),
.B2(n_1561),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1582),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1566),
.A2(n_1560),
.B1(n_769),
.B2(n_979),
.C(n_743),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1577),
.A2(n_1566),
.B(n_1569),
.C(n_1561),
.Y(n_1696)
);

AOI221x1_ASAP7_75t_L g1697 ( 
.A1(n_1560),
.A2(n_1443),
.B1(n_1235),
.B2(n_1445),
.C(n_1176),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1560),
.B(n_1566),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1586),
.A2(n_1566),
.B(n_583),
.C(n_574),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1577),
.A2(n_1560),
.B1(n_1445),
.B2(n_769),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1584),
.B(n_1435),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1428),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1567),
.B(n_1570),
.Y(n_1705)
);

OAI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1566),
.A2(n_769),
.B1(n_1586),
.B2(n_1560),
.C(n_1569),
.Y(n_1706)
);

OAI211xp5_ASAP7_75t_L g1707 ( 
.A1(n_1566),
.A2(n_1586),
.B(n_1560),
.C(n_1228),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1577),
.A2(n_1560),
.B1(n_1445),
.B2(n_769),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1428),
.Y(n_1709)
);

AO22x1_ASAP7_75t_L g1710 ( 
.A1(n_1584),
.A2(n_1560),
.B1(n_1445),
.B2(n_582),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1586),
.A2(n_1566),
.B1(n_1560),
.B2(n_1561),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1582),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1586),
.A2(n_1566),
.B1(n_1560),
.B2(n_1561),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1561),
.A2(n_1575),
.B1(n_1581),
.B2(n_1569),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1567),
.B(n_1570),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1588),
.A2(n_1599),
.B1(n_1678),
.B2(n_1701),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1671),
.B(n_1603),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1637),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1694),
.B(n_1713),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1661),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1665),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1624),
.Y(n_1725)
);

AO31x2_ASAP7_75t_L g1726 ( 
.A1(n_1605),
.A2(n_1669),
.A3(n_1697),
.B(n_1660),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1705),
.B(n_1716),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1608),
.B(n_1633),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1604),
.B(n_1615),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1597),
.B(n_1651),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1597),
.B(n_1611),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1656),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1623),
.B(n_1591),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1658),
.B(n_1673),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1613),
.B(n_1691),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1596),
.B(n_1614),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1638),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1620),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1596),
.B(n_1614),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1643),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1649),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1654),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1656),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1596),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1609),
.B(n_1662),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1634),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1613),
.B(n_1675),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1646),
.A2(n_1629),
.B(n_1605),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1592),
.B(n_1659),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1601),
.B(n_1698),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1618),
.B(n_1614),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1702),
.B(n_1639),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1702),
.B(n_1664),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1632),
.B(n_1625),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1668),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1663),
.B(n_1672),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1689),
.B(n_1628),
.Y(n_1761)
);

CKINVDCx16_ASAP7_75t_R g1762 ( 
.A(n_1676),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1644),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1628),
.B(n_1640),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1698),
.B(n_1674),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1600),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1600),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1708),
.B(n_1688),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1655),
.Y(n_1769)
);

AOI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1710),
.A2(n_1693),
.B(n_1714),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1762),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1738),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1752),
.A2(n_1695),
.B(n_1686),
.C(n_1677),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1734),
.A2(n_1690),
.B1(n_1696),
.B2(n_1590),
.C(n_1711),
.Y(n_1774)
);

AOI31xp33_ASAP7_75t_L g1775 ( 
.A1(n_1752),
.A2(n_1685),
.A3(n_1696),
.B(n_1715),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1738),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1734),
.A2(n_1587),
.B1(n_1589),
.B2(n_1712),
.C(n_1703),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1741),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1749),
.A2(n_1599),
.B1(n_1594),
.B2(n_1715),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1737),
.B(n_1680),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1769),
.A2(n_1706),
.B1(n_1692),
.B2(n_1712),
.C(n_1687),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1769),
.A2(n_1587),
.B1(n_1589),
.B2(n_1679),
.C(n_1703),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1717),
.A2(n_1679),
.B1(n_1699),
.B2(n_1687),
.C(n_1707),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1765),
.A2(n_1699),
.B(n_1700),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_SL g1785 ( 
.A(n_1765),
.B(n_1670),
.C(n_1598),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1768),
.A2(n_1670),
.B1(n_1636),
.B2(n_1616),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1742),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1742),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1762),
.B(n_1610),
.Y(n_1790)
);

OAI33xp33_ASAP7_75t_L g1791 ( 
.A1(n_1768),
.A2(n_1763),
.A3(n_1744),
.B1(n_1732),
.B2(n_1721),
.B3(n_1728),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1724),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1747),
.A2(n_1682),
.B1(n_1636),
.B2(n_1626),
.C(n_1652),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1718),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1739),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1749),
.A2(n_1612),
.B1(n_1607),
.B2(n_1640),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1747),
.A2(n_1683),
.B(n_1617),
.C(n_1709),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1735),
.B(n_1684),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1770),
.A2(n_1645),
.B1(n_1602),
.B2(n_1627),
.Y(n_1799)
);

OAI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1732),
.A2(n_1657),
.B1(n_1642),
.B2(n_1667),
.C(n_1684),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1735),
.B(n_1709),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1718),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1753),
.B(n_1622),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1728),
.B(n_1666),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1745),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1721),
.B(n_1619),
.Y(n_1806)
);

OAI33xp33_ASAP7_75t_L g1807 ( 
.A1(n_1763),
.A2(n_1595),
.A3(n_1681),
.B1(n_1667),
.B2(n_1683),
.B3(n_1621),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1744),
.B(n_1631),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_R g1809 ( 
.A(n_1770),
.B(n_1595),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1743),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1749),
.A2(n_1606),
.B1(n_1610),
.B2(n_1621),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1767),
.Y(n_1812)
);

NAND4xp25_ASAP7_75t_L g1813 ( 
.A(n_1748),
.B(n_1593),
.C(n_1681),
.D(n_1630),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1767),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1745),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1745),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1753),
.B(n_1606),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1751),
.B(n_1729),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1736),
.A2(n_1766),
.B(n_1725),
.C(n_1719),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1757),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1730),
.A2(n_1720),
.B1(n_1722),
.B2(n_1764),
.C(n_1727),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1794),
.B(n_1729),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1805),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1805),
.B(n_1737),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1776),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1776),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1820),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1778),
.B(n_1730),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1778),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1798),
.B(n_1730),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1803),
.B(n_1753),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1774),
.B(n_1750),
.C(n_1720),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1803),
.B(n_1733),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1801),
.B(n_1733),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1802),
.B(n_1751),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1733),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1820),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1818),
.B(n_1756),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1818),
.B(n_1756),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1792),
.Y(n_1843)
);

INVx4_ASAP7_75t_L g1844 ( 
.A(n_1771),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1786),
.Y(n_1845)
);

NOR2x1p5_ASAP7_75t_L g1846 ( 
.A(n_1813),
.B(n_1771),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1788),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1789),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1790),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1780),
.B(n_1723),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1812),
.B(n_1726),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1792),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1780),
.B(n_1731),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1814),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1780),
.B(n_1731),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1810),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1832),
.B(n_1816),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1822),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1806),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1843),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1830),
.B(n_1806),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1822),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1843),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1840),
.B(n_1795),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1826),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1843),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1826),
.B(n_1821),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1827),
.B(n_1775),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1827),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1828),
.B(n_1775),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1853),
.B(n_1737),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1829),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1828),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1832),
.B(n_1817),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1832),
.B(n_1817),
.Y(n_1875)
);

OAI31xp33_ASAP7_75t_L g1876 ( 
.A1(n_1834),
.A2(n_1777),
.A3(n_1793),
.B(n_1783),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1853),
.B(n_1740),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1842),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1835),
.B(n_1833),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1849),
.B(n_1807),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1840),
.B(n_1808),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1831),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1845),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1804),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1854),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1835),
.B(n_1833),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1849),
.B(n_1813),
.Y(n_1888)
);

NAND2x1_ASAP7_75t_SL g1889 ( 
.A(n_1825),
.B(n_1755),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1849),
.Y(n_1890)
);

NAND2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1844),
.B(n_1750),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1845),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1852),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1847),
.B(n_1725),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1847),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1852),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1867),
.B(n_1851),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1868),
.B(n_1834),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1858),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1900)
);

CKINVDCx14_ASAP7_75t_R g1901 ( 
.A(n_1881),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1860),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1880),
.B(n_1853),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1888),
.B(n_1791),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1890),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1887),
.B(n_1836),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1890),
.B(n_1844),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1887),
.B(n_1836),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1891),
.B(n_1838),
.Y(n_1909)
);

NAND2xp33_ASAP7_75t_R g1910 ( 
.A(n_1868),
.B(n_1809),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1886),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1888),
.B(n_1844),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1851),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1875),
.B(n_1838),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1860),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1858),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1860),
.Y(n_1917)
);

OAI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1891),
.A2(n_1889),
.B(n_1851),
.Y(n_1918)
);

AOI221x1_ASAP7_75t_SL g1919 ( 
.A1(n_1870),
.A2(n_1867),
.B1(n_1876),
.B2(n_1787),
.C(n_1773),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1863),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1886),
.B(n_1823),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1872),
.B(n_1823),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1872),
.B(n_1823),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1875),
.B(n_1838),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1876),
.A2(n_1811),
.B(n_1797),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1862),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1875),
.B(n_1855),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1862),
.B(n_1856),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1865),
.B(n_1856),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_L g1930 ( 
.A(n_1864),
.B(n_1846),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_R g1931 ( 
.A(n_1864),
.B(n_1844),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1865),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1871),
.B(n_1855),
.Y(n_1933)
);

NAND2xp33_ASAP7_75t_SL g1934 ( 
.A(n_1889),
.B(n_1846),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1871),
.B(n_1855),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1869),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1891),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1871),
.B(n_1850),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1869),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1891),
.B(n_1785),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1873),
.B(n_1848),
.Y(n_1941)
);

OAI321xp33_ASAP7_75t_L g1942 ( 
.A1(n_1898),
.A2(n_1897),
.A3(n_1913),
.B1(n_1912),
.B2(n_1904),
.C(n_1919),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1902),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1904),
.A2(n_1796),
.B1(n_1779),
.B2(n_1750),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1902),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1902),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1931),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1899),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1919),
.B(n_1885),
.Y(n_1949)
);

AOI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1940),
.A2(n_1781),
.A3(n_1782),
.B1(n_1799),
.B2(n_1764),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1899),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1898),
.B(n_1885),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1914),
.B(n_1871),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1901),
.B(n_1844),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1911),
.B(n_1859),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_SL g1956 ( 
.A1(n_1930),
.A2(n_1784),
.B(n_1879),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1916),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1930),
.A2(n_1859),
.B1(n_1861),
.B2(n_1877),
.Y(n_1958)
);

AOI222xp33_ASAP7_75t_L g1959 ( 
.A1(n_1940),
.A2(n_1764),
.B1(n_1720),
.B2(n_1722),
.C1(n_1746),
.C2(n_1758),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1925),
.B(n_1841),
.Y(n_1960)
);

AND2x2_ASAP7_75t_SL g1961 ( 
.A(n_1905),
.B(n_1750),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1921),
.B(n_1861),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1916),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1926),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1926),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1932),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1915),
.Y(n_1967)
);

OAI322xp33_ASAP7_75t_L g1968 ( 
.A1(n_1897),
.A2(n_1829),
.A3(n_1839),
.B1(n_1882),
.B2(n_1841),
.C1(n_1837),
.C2(n_1873),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1914),
.B(n_1877),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1932),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1936),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1911),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1925),
.A2(n_1839),
.B(n_1819),
.C(n_1879),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_L g1974 ( 
.A(n_1934),
.B(n_1879),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1905),
.B(n_1882),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1905),
.B(n_1874),
.Y(n_1976)
);

OAI321xp33_ASAP7_75t_L g1977 ( 
.A1(n_1913),
.A2(n_1800),
.A3(n_1804),
.B1(n_1758),
.B2(n_1754),
.C(n_1722),
.Y(n_1977)
);

AOI222xp33_ASAP7_75t_L g1978 ( 
.A1(n_1922),
.A2(n_1746),
.B1(n_1761),
.B2(n_1759),
.C1(n_1760),
.C2(n_1866),
.Y(n_1978)
);

NOR4xp25_ASAP7_75t_L g1979 ( 
.A(n_1942),
.B(n_1937),
.C(n_1921),
.D(n_1923),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1961),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1973),
.B(n_1907),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1953),
.B(n_1924),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1961),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1949),
.B(n_1905),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1960),
.B(n_1922),
.Y(n_1985)
);

OAI31xp33_ASAP7_75t_L g1986 ( 
.A1(n_1956),
.A2(n_1937),
.A3(n_1909),
.B(n_1923),
.Y(n_1986)
);

AOI32xp33_ASAP7_75t_L g1987 ( 
.A1(n_1977),
.A2(n_1952),
.A3(n_1958),
.B1(n_1974),
.B2(n_1918),
.Y(n_1987)
);

AO22x1_ASAP7_75t_L g1988 ( 
.A1(n_1972),
.A2(n_1909),
.B1(n_1910),
.B2(n_1903),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1948),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1962),
.B(n_1928),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1948),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1953),
.B(n_1924),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1968),
.A2(n_1909),
.B1(n_1939),
.B2(n_1936),
.C(n_1915),
.Y(n_1993)
);

AOI222xp33_ASAP7_75t_L g1994 ( 
.A1(n_1944),
.A2(n_1918),
.B1(n_1920),
.B2(n_1917),
.C1(n_1915),
.C2(n_1939),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1951),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1947),
.A2(n_1903),
.B1(n_1877),
.B2(n_1927),
.Y(n_1996)
);

NOR2x1_ASAP7_75t_L g1997 ( 
.A(n_1954),
.B(n_1903),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1969),
.B(n_1927),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1951),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1950),
.B(n_1900),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1943),
.A2(n_1918),
.B(n_1917),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1974),
.A2(n_1941),
.B(n_1928),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1943),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1965),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1975),
.Y(n_2005)
);

XOR2x2_ASAP7_75t_L g2006 ( 
.A(n_2000),
.B(n_1750),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_2001),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1991),
.Y(n_2008)
);

NAND2x1_ASAP7_75t_L g2009 ( 
.A(n_1997),
.B(n_1969),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1979),
.B(n_1955),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_L g2011 ( 
.A(n_1984),
.B(n_1987),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1991),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1980),
.B(n_1962),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1995),
.Y(n_2014)
);

AOI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_1994),
.A2(n_1967),
.B(n_1946),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_2003),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1995),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1981),
.B(n_1976),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1980),
.B(n_1900),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1999),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1999),
.Y(n_2021)
);

OAI31xp33_ASAP7_75t_L g2022 ( 
.A1(n_1986),
.A2(n_1945),
.A3(n_1967),
.B(n_1946),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2004),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1982),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2004),
.Y(n_2025)
);

NAND4xp25_ASAP7_75t_L g2026 ( 
.A(n_2018),
.B(n_2010),
.C(n_2024),
.D(n_2013),
.Y(n_2026)
);

NOR3xp33_ASAP7_75t_SL g2027 ( 
.A(n_2018),
.B(n_1996),
.C(n_1985),
.Y(n_2027)
);

NOR3xp33_ASAP7_75t_SL g2028 ( 
.A(n_2019),
.B(n_2002),
.C(n_1988),
.Y(n_2028)
);

NOR4xp25_ASAP7_75t_L g2029 ( 
.A(n_2011),
.B(n_2005),
.C(n_1983),
.D(n_1989),
.Y(n_2029)
);

NAND4xp25_ASAP7_75t_L g2030 ( 
.A(n_2024),
.B(n_1993),
.C(n_1990),
.D(n_1988),
.Y(n_2030)
);

NAND4xp25_ASAP7_75t_SL g2031 ( 
.A(n_2022),
.B(n_1998),
.C(n_1982),
.D(n_1992),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2007),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2007),
.Y(n_2033)
);

NAND3xp33_ASAP7_75t_L g2034 ( 
.A(n_2011),
.B(n_1983),
.C(n_2003),
.Y(n_2034)
);

NOR4xp25_ASAP7_75t_L g2035 ( 
.A(n_2016),
.B(n_1990),
.C(n_1965),
.D(n_1966),
.Y(n_2035)
);

NAND3xp33_ASAP7_75t_L g2036 ( 
.A(n_2015),
.B(n_1959),
.C(n_1957),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_SL g2037 ( 
.A(n_2016),
.B(n_1992),
.Y(n_2037)
);

NOR3xp33_ASAP7_75t_L g2038 ( 
.A(n_2009),
.B(n_2025),
.C(n_2023),
.Y(n_2038)
);

AOI222xp33_ASAP7_75t_L g2039 ( 
.A1(n_2036),
.A2(n_2006),
.B1(n_2021),
.B2(n_2008),
.C1(n_2020),
.C2(n_2014),
.Y(n_2039)
);

AOI222xp33_ASAP7_75t_L g2040 ( 
.A1(n_2034),
.A2(n_2017),
.B1(n_2012),
.B2(n_1945),
.C1(n_1966),
.C2(n_1971),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2026),
.A2(n_2001),
.B1(n_1978),
.B2(n_1917),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_R g2042 ( 
.A(n_2028),
.B(n_2001),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2037),
.B(n_1998),
.Y(n_2043)
);

AOI222xp33_ASAP7_75t_L g2044 ( 
.A1(n_2032),
.A2(n_2033),
.B1(n_2029),
.B2(n_2035),
.C1(n_2030),
.C2(n_1970),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_2031),
.A2(n_2038),
.B1(n_2027),
.B2(n_1963),
.C(n_1964),
.Y(n_2045)
);

OAI211xp5_ASAP7_75t_SL g2046 ( 
.A1(n_2028),
.A2(n_1941),
.B(n_1929),
.C(n_1920),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_2026),
.B(n_1906),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2037),
.B(n_1906),
.Y(n_2048)
);

NAND2xp67_ASAP7_75t_SL g2049 ( 
.A(n_2029),
.B(n_1933),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2043),
.B(n_1908),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2042),
.Y(n_2051)
);

NAND2xp33_ASAP7_75t_R g2052 ( 
.A(n_2047),
.B(n_1903),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2048),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_2046),
.A2(n_1920),
.B(n_1908),
.Y(n_2054)
);

BUFx12f_ASAP7_75t_L g2055 ( 
.A(n_2049),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_2041),
.A2(n_1929),
.B1(n_1896),
.B2(n_1866),
.C(n_1863),
.Y(n_2056)
);

AND3x4_ASAP7_75t_L g2057 ( 
.A(n_2052),
.B(n_2055),
.C(n_2039),
.Y(n_2057)
);

NAND4xp75_ASAP7_75t_L g2058 ( 
.A(n_2053),
.B(n_2045),
.C(n_2044),
.D(n_2040),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_2051),
.B(n_1933),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2050),
.B(n_1878),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2054),
.B(n_2056),
.C(n_1866),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_SL g2062 ( 
.A1(n_2053),
.A2(n_1854),
.B1(n_1935),
.B2(n_1938),
.C(n_1895),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2051),
.A2(n_1935),
.B(n_1938),
.Y(n_2063)
);

NOR2x1p5_ASAP7_75t_L g2064 ( 
.A(n_2058),
.B(n_1824),
.Y(n_2064)
);

NOR2x2_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_1754),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2059),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_2062),
.B(n_2063),
.Y(n_2067)
);

INVxp33_ASAP7_75t_SL g2068 ( 
.A(n_2060),
.Y(n_2068)
);

OAI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2061),
.A2(n_1896),
.B1(n_1893),
.B2(n_1863),
.C(n_1883),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2066),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2067),
.B(n_1878),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2068),
.B(n_1883),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2064),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2070),
.Y(n_2074)
);

XNOR2xp5_ASAP7_75t_L g2075 ( 
.A(n_2074),
.B(n_2073),
.Y(n_2075)
);

XNOR2xp5_ASAP7_75t_L g2076 ( 
.A(n_2075),
.B(n_2071),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2075),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2076),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2077),
.B(n_2072),
.Y(n_2079)
);

INVxp67_ASAP7_75t_L g2080 ( 
.A(n_2078),
.Y(n_2080)
);

OAI222xp33_ASAP7_75t_L g2081 ( 
.A1(n_2079),
.A2(n_2069),
.B1(n_2065),
.B2(n_1884),
.C1(n_1892),
.C2(n_1895),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2080),
.Y(n_2082)
);

AOI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2082),
.A2(n_2081),
.B1(n_1892),
.B2(n_1884),
.C(n_1896),
.Y(n_2083)
);

AOI211xp5_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_1894),
.B(n_1874),
.C(n_1857),
.Y(n_2084)
);


endmodule