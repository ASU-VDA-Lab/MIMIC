module fake_jpeg_5358_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_54),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_59),
.Y(n_66)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_39),
.B1(n_17),
.B2(n_20),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_65),
.A2(n_67),
.B1(n_100),
.B2(n_95),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_21),
.B(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_20),
.B1(n_17),
.B2(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_69),
.B1(n_82),
.B2(n_106),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_20),
.B1(n_39),
.B2(n_21),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_72),
.Y(n_140)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_87),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_18),
.B1(n_34),
.B2(n_30),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_79),
.B1(n_14),
.B2(n_12),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_18),
.B1(n_34),
.B2(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_38),
.B1(n_22),
.B2(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_45),
.A2(n_38),
.B1(n_22),
.B2(n_24),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_109),
.B1(n_95),
.B2(n_107),
.Y(n_110)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_90),
.Y(n_124)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_26),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_103),
.Y(n_125)
);

AO22x2_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_0),
.B2(n_1),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_26),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_37),
.B1(n_23),
.B2(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_0),
.Y(n_122)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_33),
.C(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_10),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_43),
.A2(n_37),
.B1(n_23),
.B2(n_27),
.Y(n_106)
);

NAND2xp67_ASAP7_75t_SL g107 ( 
.A(n_62),
.B(n_8),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_95),
.B1(n_9),
.B2(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_33),
.B1(n_37),
.B2(n_2),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_138),
.B1(n_145),
.B2(n_136),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_136),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_78),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_109),
.B1(n_93),
.B2(n_74),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_101),
.B(n_81),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_139),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_113),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_67),
.A2(n_9),
.B1(n_8),
.B2(n_3),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_1),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_119),
.Y(n_169)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_66),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_66),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_120),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_97),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_136),
.B1(n_130),
.B2(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_162),
.B1(n_172),
.B2(n_180),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_96),
.B(n_105),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_170),
.B1(n_181),
.B2(n_134),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_175),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_80),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_71),
.C(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_81),
.B(n_75),
.C(n_64),
.Y(n_174)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_171),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_129),
.A2(n_85),
.B1(n_78),
.B2(n_84),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_74),
.B1(n_92),
.B2(n_84),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_114),
.B1(n_131),
.B2(n_117),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_186),
.B1(n_202),
.B2(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_126),
.B1(n_85),
.B2(n_140),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_122),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_195),
.B(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_173),
.B1(n_172),
.B2(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_206),
.C(n_167),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_118),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_104),
.B(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_116),
.B1(n_104),
.B2(n_127),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_204),
.B1(n_209),
.B2(n_166),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_142),
.B1(n_119),
.B2(n_135),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_3),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_208),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_144),
.B1(n_5),
.B2(n_6),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_7),
.C(n_155),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_174),
.B1(n_150),
.B2(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_150),
.A2(n_181),
.B1(n_149),
.B2(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_152),
.B(n_148),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_219),
.B1(n_221),
.B2(n_223),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_229),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_179),
.B1(n_156),
.B2(n_148),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_155),
.B1(n_169),
.B2(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_194),
.C(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_155),
.B1(n_168),
.B2(n_167),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_231),
.B1(n_233),
.B2(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_156),
.B1(n_176),
.B2(n_171),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_176),
.B(n_175),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_175),
.B1(n_178),
.B2(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_212),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_190),
.B(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_195),
.B1(n_206),
.B2(n_211),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_246),
.B1(n_255),
.B2(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_185),
.B1(n_182),
.B2(n_190),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_258),
.C(n_227),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_205),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_253),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_225),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_203),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_217),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_260),
.B1(n_184),
.B2(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_214),
.C(n_210),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

NAND4xp25_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_234),
.C(n_231),
.D(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_196),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_262),
.A2(n_237),
.B1(n_233),
.B2(n_226),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_272),
.B1(n_241),
.B2(n_244),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.C(n_274),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_250),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_267),
.A2(n_250),
.B(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_239),
.C(n_227),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_245),
.A2(n_222),
.B1(n_228),
.B2(n_231),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_222),
.C(n_225),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_223),
.A3(n_228),
.B1(n_232),
.B2(n_215),
.C1(n_234),
.C2(n_220),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_249),
.C(n_256),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_233),
.C(n_184),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_260),
.C(n_242),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_241),
.B1(n_245),
.B2(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_277),
.B1(n_265),
.B2(n_266),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_289),
.B(n_290),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_261),
.B1(n_247),
.B2(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_261),
.B1(n_247),
.B2(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.C(n_274),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_252),
.B1(n_255),
.B2(n_187),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_278),
.B1(n_267),
.B2(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_300),
.Y(n_306)
);

NAND2xp67_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_255),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_302),
.B(n_291),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_263),
.B(n_270),
.C(n_264),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_283),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_268),
.C(n_187),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_213),
.B1(n_220),
.B2(n_288),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_284),
.B(n_286),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_280),
.B1(n_282),
.B2(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_295),
.B(n_294),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_285),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_293),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_303),
.B(n_310),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_315),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.C(n_312),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_318),
.C(n_314),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_306),
.Y(n_325)
);


endmodule