module fake_jpeg_10979_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_14),
.B1(n_31),
.B2(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_37),
.C(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_42),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_38),
.B1(n_34),
.B2(n_4),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_76),
.B1(n_8),
.B2(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_15),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_38),
.C(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_32),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_57),
.B(n_65),
.C(n_54),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_12),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_85),
.A3(n_87),
.B1(n_88),
.B2(n_89),
.C1(n_77),
.C2(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_11),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_16),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_96),
.C(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_74),
.B1(n_66),
.B2(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_85),
.B1(n_83),
.B2(n_23),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

NAND2x1p5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_83),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_94),
.A3(n_95),
.B1(n_92),
.B2(n_96),
.C(n_26),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_19),
.C(n_20),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_25),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_100),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_94),
.Y(n_106)
);


endmodule