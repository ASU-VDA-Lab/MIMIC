module fake_jpeg_20587_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_3),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_18),
.B(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_2),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_75),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_69),
.B1(n_43),
.B2(n_3),
.Y(n_78)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_40),
.B1(n_54),
.B2(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_44),
.B1(n_52),
.B2(n_49),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_82),
.B1(n_74),
.B2(n_68),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_50),
.B(n_45),
.C(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_85),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_19),
.B1(n_35),
.B2(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_4),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_84),
.C(n_9),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_77),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_102),
.B(n_92),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_84),
.C(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_90),
.B(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_102),
.B1(n_99),
.B2(n_91),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_106),
.B1(n_107),
.B2(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_111),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_23),
.C(n_24),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_27),
.B(n_28),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_29),
.Y(n_115)
);


endmodule