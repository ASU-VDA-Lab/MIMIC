module real_jpeg_21100_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_2),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_31),
.B1(n_48),
.B2(n_49),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_135),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_135),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_135),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_4),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_167),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_167),
.Y(n_223)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_6),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_161),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_161),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_7),
.B(n_24),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_14),
.B(n_49),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_165),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_80),
.B1(n_174),
.B2(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_7),
.B(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_7),
.B(n_27),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_7),
.A2(n_27),
.B(n_247),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_8),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_94),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.C(n_76),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_20),
.B(n_67),
.CI(n_76),
.CON(n_139),
.SN(n_139)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_21),
.A2(n_22),
.B1(n_96),
.B2(n_109),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_22),
.B(n_39),
.C(n_55),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_23),
.A2(n_28),
.B1(n_90),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_23),
.A2(n_90),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_23),
.A2(n_90),
.B1(n_134),
.B2(n_179),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_24),
.B(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_24),
.A2(n_35),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_25),
.A2(n_36),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_25),
.A2(n_42),
.A3(n_59),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_27),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_58),
.Y(n_60)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g164 ( 
.A(n_30),
.B(n_165),
.CON(n_164),
.SN(n_164)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_40),
.B1(n_101),
.B2(n_107),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_41),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_41),
.A2(n_47),
.B1(n_86),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_41),
.A2(n_51),
.B(n_87),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_41),
.A2(n_47),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_41),
.A2(n_47),
.B1(n_218),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_41),
.A2(n_47),
.B1(n_238),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_41),
.A2(n_71),
.B(n_254),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_43),
.A2(n_50),
.B(n_165),
.C(n_214),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g248 ( 
.A(n_43),
.B(n_58),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_47),
.A2(n_73),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_47),
.B(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_48),
.B(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_65),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_56),
.A2(n_103),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_56),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_56),
.A2(n_65),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_57),
.A2(n_61),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_57),
.A2(n_61),
.B1(n_196),
.B2(n_251),
.Y(n_250)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_69),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_66),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_68),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_89),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_78),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_80),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_80),
.A2(n_150),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_80),
.A2(n_82),
.B1(n_208),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_80),
.A2(n_128),
.B(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_81),
.A2(n_129),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_81),
.A2(n_84),
.B(n_152),
.Y(n_245)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_127),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_85),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_108),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_104),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_316),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_139),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_115),
.B(n_139),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_116),
.B(n_120),
.Y(n_314)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_121),
.A2(n_122),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.C(n_137),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_123),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_124),
.B(n_130),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_173),
.B(n_174),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_139),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_310),
.B(n_315),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_298),
.B(n_309),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_199),
.B(n_277),
.C(n_297),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_184),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_144),
.B(n_184),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_168),
.B2(n_183),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_147),
.B(n_155),
.C(n_183),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_148),
.B(n_154),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_163),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_174),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_169),
.B(n_176),
.C(n_181),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_194),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_276),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_271),
.B(n_275),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_259),
.B(n_270),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_241),
.B(n_258),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_230),
.B(n_240),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_219),
.B(n_229),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_215),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_232),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_249),
.B1(n_256),
.B2(n_257),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_295),
.B2(n_296),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_285),
.C(n_296),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_294),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_292),
.C(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_306),
.C(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);


endmodule