module fake_jpeg_1246_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_57),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_62),
.B1(n_65),
.B2(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_93),
.B1(n_56),
.B2(n_75),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_62),
.B1(n_70),
.B2(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_64),
.B1(n_79),
.B2(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_61),
.C(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_96),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_55),
.B(n_67),
.C(n_68),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_111),
.B1(n_51),
.B2(n_48),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_83),
.B1(n_79),
.B2(n_61),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_110),
.B1(n_114),
.B2(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_32),
.B(n_40),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_42),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_56),
.B1(n_73),
.B2(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_71),
.B1(n_69),
.B2(n_68),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_71),
.B1(n_69),
.B2(n_75),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_94),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_131),
.C(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_132),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_136),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_14),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_130),
.B1(n_12),
.B2(n_13),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_44),
.C(n_43),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_109),
.A3(n_106),
.B1(n_101),
.B2(n_10),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_134),
.B(n_16),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_6),
.B(n_7),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_149),
.B1(n_157),
.B2(n_131),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_38),
.B1(n_35),
.B2(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_151),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_15),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_26),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_16),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_24),
.B1(n_18),
.B2(n_19),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_22),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_122),
.C(n_123),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_169),
.C(n_126),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_177),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_141),
.C(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_133),
.B(n_123),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_153),
.C(n_137),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_185),
.C(n_186),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_188),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_163),
.B1(n_174),
.B2(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_164),
.C(n_170),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_151),
.C(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_144),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_176),
.C(n_163),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_166),
.B1(n_165),
.B2(n_167),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_189),
.B(n_162),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_161),
.C(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_203),
.B1(n_181),
.B2(n_187),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_208),
.B1(n_201),
.B2(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_190),
.B(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_207),
.A2(n_171),
.B1(n_147),
.B2(n_20),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_193),
.C(n_143),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_209),
.C(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_210),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_17),
.B(n_18),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_17),
.B(n_20),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_21),
.Y(n_216)
);


endmodule