module real_aes_8755_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_1), .A2(n_156), .B(n_168), .C(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g275 ( .A(n_2), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_3), .A2(n_183), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_4), .B(n_179), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g182 ( .A1(n_5), .A2(n_183), .B(n_184), .Y(n_182) );
AND2x6_ASAP7_75t_L g156 ( .A(n_6), .B(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_8), .B(n_42), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_8), .B(n_42), .Y(n_129) );
INVx1_ASAP7_75t_L g482 ( .A(n_9), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_10), .B(n_189), .Y(n_470) );
INVx1_ASAP7_75t_L g191 ( .A(n_11), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_12), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g153 ( .A(n_13), .Y(n_153) );
INVx1_ASAP7_75t_L g257 ( .A(n_14), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_15), .A2(n_192), .B(n_258), .C(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_16), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_16), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_17), .B(n_179), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_18), .B(n_202), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_19), .B(n_183), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_524), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_21), .A2(n_159), .B(n_243), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_22), .B(n_179), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_23), .B(n_189), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_24), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_25), .B(n_189), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_26), .Y(n_541) );
INVx1_ASAP7_75t_L g531 ( .A(n_27), .Y(n_531) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_28), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_29), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_30), .B(n_189), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_31), .A2(n_66), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_31), .Y(n_739) );
INVx1_ASAP7_75t_L g520 ( .A(n_32), .Y(n_520) );
INVx1_ASAP7_75t_L g167 ( .A(n_33), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_34), .A2(n_104), .B1(n_117), .B2(n_742), .Y(n_103) );
INVx2_ASAP7_75t_L g161 ( .A(n_35), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_36), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_37), .A2(n_193), .B(n_243), .C(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g521 ( .A(n_38), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_39), .A2(n_156), .B(n_168), .C(n_213), .Y(n_212) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_40), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_168), .B(n_530), .C(n_534), .Y(n_529) );
INVx1_ASAP7_75t_L g165 ( .A(n_43), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_44), .A2(n_188), .B(n_218), .C(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_45), .B(n_189), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_46), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_47), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_48), .Y(n_517) );
INVx1_ASAP7_75t_L g497 ( .A(n_49), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_50), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_51), .B(n_183), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_52), .A2(n_159), .B1(n_162), .B2(n_168), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_53), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_54), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_55), .A2(n_188), .B(n_190), .C(n_193), .Y(n_187) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_56), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_57), .Y(n_232) );
INVx1_ASAP7_75t_L g185 ( .A(n_58), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_59), .A2(n_736), .B1(n_737), .B2(n_740), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_59), .Y(n_740) );
INVx1_ASAP7_75t_L g157 ( .A(n_60), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_61), .A2(n_77), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_61), .Y(n_138) );
INVx1_ASAP7_75t_L g152 ( .A(n_62), .Y(n_152) );
INVx1_ASAP7_75t_SL g510 ( .A(n_63), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_64), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_65), .B(n_179), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_66), .Y(n_738) );
INVx1_ASAP7_75t_L g544 ( .A(n_67), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_SL g201 ( .A1(n_68), .A2(n_193), .B(n_202), .C(n_203), .Y(n_201) );
INVxp67_ASAP7_75t_L g204 ( .A(n_69), .Y(n_204) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_71), .A2(n_183), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_72), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_73), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_74), .A2(n_183), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g225 ( .A(n_75), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_251), .B(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_77), .Y(n_137) );
INVx1_ASAP7_75t_L g489 ( .A(n_78), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_79), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_80), .A2(n_156), .B(n_168), .C(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_81), .A2(n_183), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g492 ( .A(n_82), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
INVx1_ASAP7_75t_L g468 ( .A(n_85), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_86), .B(n_202), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_87), .A2(n_156), .B(n_168), .C(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g113 ( .A(n_88), .Y(n_113) );
OR2x2_ASAP7_75t_L g126 ( .A(n_88), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g723 ( .A(n_88), .B(n_128), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_89), .A2(n_168), .B(n_543), .C(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_90), .B(n_196), .Y(n_195) );
AOI222xp33_ASAP7_75t_SL g131 ( .A1(n_91), .A2(n_132), .B1(n_133), .B2(n_139), .C1(n_724), .C2(n_728), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_92), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_93), .A2(n_156), .B(n_168), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_94), .Y(n_247) );
INVx1_ASAP7_75t_L g200 ( .A(n_95), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_96), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_97), .B(n_215), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_98), .B(n_181), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_99), .B(n_181), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_101), .A2(n_183), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g500 ( .A(n_102), .Y(n_500) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g742 ( .A(n_106), .Y(n_742) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g128 ( .A(n_112), .B(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g455 ( .A(n_113), .B(n_128), .Y(n_455) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_113), .B(n_127), .Y(n_730) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_131), .B1(n_731), .B2(n_732), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g731 ( .A(n_122), .Y(n_731) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_124), .A2(n_733), .B(n_741), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_130), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_126), .Y(n_741) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_453), .B1(n_456), .B2(n_723), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_141), .A2(n_453), .B1(n_725), .B2(n_726), .Y(n_724) );
AND3x1_ASAP7_75t_L g141 ( .A(n_142), .B(n_378), .C(n_427), .Y(n_141) );
NOR3xp33_ASAP7_75t_SL g142 ( .A(n_143), .B(n_285), .C(n_323), .Y(n_142) );
OAI222xp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_206), .B1(n_260), .B2(n_266), .C1(n_280), .C2(n_283), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_177), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_145), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_145), .B(n_328), .Y(n_419) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g296 ( .A(n_146), .B(n_197), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_146), .B(n_178), .Y(n_304) );
AND2x2_ASAP7_75t_L g339 ( .A(n_146), .B(n_316), .Y(n_339) );
OR2x2_ASAP7_75t_L g363 ( .A(n_146), .B(n_178), .Y(n_363) );
OR2x2_ASAP7_75t_L g371 ( .A(n_146), .B(n_270), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_146), .B(n_197), .Y(n_374) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g268 ( .A(n_147), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_147), .B(n_197), .Y(n_282) );
AND2x2_ASAP7_75t_L g332 ( .A(n_147), .B(n_270), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_147), .B(n_178), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_147), .B(n_431), .Y(n_452) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_154), .B(n_175), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_148), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_148), .A2(n_271), .B(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_150), .B(n_151), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B1(n_171), .B2(n_172), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_186), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_155), .A2(n_186), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_155), .A2(n_186), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_155), .A2(n_186), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_155), .A2(n_186), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_155), .A2(n_186), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_155), .A2(n_186), .B(n_517), .C(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g546 ( .A(n_155), .Y(n_546) );
INVx4_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_156), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g183 ( .A(n_156), .B(n_173), .Y(n_183) );
BUFx3_ASAP7_75t_L g534 ( .A(n_156), .Y(n_534) );
INVx2_ASAP7_75t_L g277 ( .A(n_159), .Y(n_277) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g169 ( .A(n_161), .Y(n_169) );
INVx1_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_162) );
INVx2_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
INVx4_ASAP7_75t_L g255 ( .A(n_163), .Y(n_255) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
AND2x2_ASAP7_75t_L g173 ( .A(n_164), .B(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_164), .Y(n_189) );
INVx3_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx1_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
INVx2_ASAP7_75t_L g469 ( .A(n_166), .Y(n_469) );
INVx5_ASAP7_75t_L g186 ( .A(n_168), .Y(n_186) );
AND2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
BUFx3_ASAP7_75t_L g219 ( .A(n_169), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_172), .A2(n_225), .B(n_226), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_172), .A2(n_272), .B(n_273), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_172), .A2(n_465), .B(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_172), .A2(n_196), .B(n_528), .C(n_529), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_172), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g522 ( .A(n_174), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_177), .A2(n_371), .B(n_372), .C(n_375), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_177), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_177), .B(n_315), .Y(n_437) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_197), .Y(n_177) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_178), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g295 ( .A(n_178), .Y(n_295) );
AND2x2_ASAP7_75t_L g322 ( .A(n_178), .B(n_316), .Y(n_322) );
INVx1_ASAP7_75t_SL g330 ( .A(n_178), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_178), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g431 ( .A(n_178), .Y(n_431) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_195), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g221 ( .A(n_180), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_180), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_180), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_180), .A2(n_540), .B(n_547), .Y(n_539) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_198), .B(n_205), .Y(n_197) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_181), .Y(n_486) );
BUFx2_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx4_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_192), .B(n_204), .Y(n_203) );
INVx5_ASAP7_75t_L g215 ( .A(n_192), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_192), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_194), .Y(n_244) );
INVx1_ASAP7_75t_L g233 ( .A(n_196), .Y(n_233) );
INVx2_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_196), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_196), .A2(n_477), .B(n_483), .Y(n_476) );
BUFx2_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
INVx1_ASAP7_75t_L g329 ( .A(n_197), .Y(n_329) );
INVx3_ASAP7_75t_L g354 ( .A(n_197), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_206), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_234), .Y(n_206) );
INVx1_ASAP7_75t_L g350 ( .A(n_207), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g356 ( .A1(n_207), .A2(n_295), .A3(n_357), .B1(n_358), .B2(n_359), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_207), .A2(n_361), .B1(n_364), .B2(n_369), .Y(n_360) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g298 ( .A(n_208), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g376 ( .A(n_208), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g446 ( .A(n_208), .B(n_392), .Y(n_446) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_223), .Y(n_208) );
AND2x2_ASAP7_75t_L g261 ( .A(n_209), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
INVx1_ASAP7_75t_L g310 ( .A(n_209), .Y(n_310) );
OR2x2_ASAP7_75t_L g318 ( .A(n_209), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_209), .B(n_299), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_209), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g346 ( .A(n_209), .B(n_264), .Y(n_346) );
INVx3_ASAP7_75t_L g368 ( .A(n_209), .Y(n_368) );
AND2x2_ASAP7_75t_L g393 ( .A(n_209), .B(n_265), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_209), .B(n_358), .Y(n_441) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_216), .B(n_217), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_215), .A2(n_275), .B(n_276), .C(n_277), .Y(n_274) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_215), .A2(n_255), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_215), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g467 ( .A1(n_217), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_217), .A2(n_469), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
INVx1_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AND2x2_ASAP7_75t_L g397 ( .A(n_223), .B(n_235), .Y(n_397) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_230), .B(n_231), .Y(n_223) );
INVx1_ASAP7_75t_L g514 ( .A(n_230), .Y(n_514) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_230), .A2(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_233), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_233), .B(n_279), .Y(n_278) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_233), .A2(n_464), .B(n_471), .Y(n_463) );
INVx2_ASAP7_75t_L g439 ( .A(n_234), .Y(n_439) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_248), .Y(n_234) );
INVx1_ASAP7_75t_L g284 ( .A(n_235), .Y(n_284) );
AND2x2_ASAP7_75t_L g311 ( .A(n_235), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_235), .B(n_265), .Y(n_319) );
AND2x2_ASAP7_75t_L g377 ( .A(n_235), .B(n_300), .Y(n_377) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
AND2x2_ASAP7_75t_L g290 ( .A(n_236), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_236), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_236), .B(n_265), .Y(n_365) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
INVx1_ASAP7_75t_L g524 ( .A(n_237), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_237), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_243), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_248), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_248), .B(n_265), .Y(n_358) );
AND2x2_ASAP7_75t_L g367 ( .A(n_248), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g392 ( .A(n_248), .Y(n_392) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g264 ( .A(n_249), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_255), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_255), .B(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_270), .B1(n_429), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_262), .A2(n_373), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_263), .B(n_368), .Y(n_385) );
INVx1_ASAP7_75t_L g410 ( .A(n_263), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_264), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g337 ( .A(n_264), .B(n_290), .Y(n_337) );
INVx2_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_266), .A2(n_418), .B1(n_435), .B2(n_438), .C(n_440), .Y(n_434) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_267), .B(n_316), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_268), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g359 ( .A(n_268), .B(n_305), .Y(n_359) );
INVx3_ASAP7_75t_SL g400 ( .A(n_268), .Y(n_400) );
AND2x2_ASAP7_75t_L g344 ( .A(n_269), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g373 ( .A(n_269), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_269), .B(n_282), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_269), .B(n_328), .Y(n_414) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g316 ( .A(n_270), .Y(n_316) );
OAI322xp33_ASAP7_75t_L g411 ( .A1(n_270), .A2(n_342), .A3(n_364), .B1(n_412), .B2(n_414), .C1(n_415), .C2(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_281), .A2(n_284), .B(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_SL g361 ( .A(n_282), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g383 ( .A(n_282), .B(n_295), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_282), .B(n_322), .Y(n_398) );
INVxp67_ASAP7_75t_L g349 ( .A(n_284), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_284), .A2(n_356), .B(n_360), .C(n_370), .Y(n_355) );
OAI221xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_294), .B1(n_297), .B2(n_301), .C(n_306), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_293), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g426 ( .A(n_293), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_294), .A2(n_443), .B1(n_448), .B2(n_449), .C(n_451), .Y(n_442) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_295), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_295), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_295), .B(n_373), .Y(n_380) );
AND2x2_ASAP7_75t_L g422 ( .A(n_295), .B(n_400), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_296), .B(n_321), .Y(n_320) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_296), .A2(n_308), .B1(n_418), .B2(n_419), .Y(n_417) );
OR2x2_ASAP7_75t_L g448 ( .A(n_296), .B(n_316), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g425 ( .A(n_299), .Y(n_425) );
AND2x2_ASAP7_75t_L g450 ( .A(n_299), .B(n_393), .Y(n_450) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_304), .B(n_315), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_317), .B2(n_320), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g381 ( .A(n_309), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_309), .B(n_349), .Y(n_416) );
AOI322xp5_ASAP7_75t_L g340 ( .A1(n_311), .A2(n_341), .A3(n_343), .B1(n_344), .B2(n_346), .C1(n_347), .C2(n_351), .Y(n_340) );
INVxp67_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_314), .A2(n_319), .B1(n_336), .B2(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_315), .B(n_328), .Y(n_415) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_316), .B(n_354), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_316), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g412 ( .A(n_318), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_340), .C(n_355), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_331), .B2(n_333), .C(n_335), .Y(n_324) );
AND2x2_ASAP7_75t_L g331 ( .A(n_327), .B(n_332), .Y(n_331) );
INVx3_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g341 ( .A(n_332), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_334), .Y(n_413) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_339), .B(n_353), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_342), .B(n_400), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_343), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g418 ( .A(n_346), .Y(n_418) );
AND2x2_ASAP7_75t_L g433 ( .A(n_346), .B(n_410), .Y(n_433) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_357), .A2(n_428), .B(n_434), .C(n_442), .Y(n_427) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g396 ( .A(n_367), .B(n_397), .Y(n_396) );
NAND2x1_ASAP7_75t_SL g438 ( .A(n_368), .B(n_439), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_371), .Y(n_408) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
AND2x2_ASAP7_75t_L g407 ( .A(n_377), .B(n_393), .Y(n_407) );
NOR5xp2_ASAP7_75t_L g378 ( .A(n_379), .B(n_394), .C(n_411), .D(n_417), .E(n_420), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_386), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_383), .B(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g409 ( .A(n_393), .B(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_398), .B1(n_399), .B2(n_401), .C(n_404), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
AOI211xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_423), .B(n_425), .C(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g725 ( .A(n_456), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_456), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_678), .Y(n_456) );
NAND5xp2_ASAP7_75t_L g457 ( .A(n_458), .B(n_590), .C(n_628), .D(n_649), .E(n_666), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_562), .C(n_583), .Y(n_458) );
OAI221xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_502), .B1(n_525), .B2(n_549), .C(n_553), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_473), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_462), .B(n_551), .Y(n_570) );
OR2x2_ASAP7_75t_L g597 ( .A(n_462), .B(n_485), .Y(n_597) );
AND2x2_ASAP7_75t_L g611 ( .A(n_462), .B(n_485), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_462), .B(n_476), .Y(n_625) );
AND2x2_ASAP7_75t_L g663 ( .A(n_462), .B(n_627), .Y(n_663) );
AND2x2_ASAP7_75t_L g692 ( .A(n_462), .B(n_602), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_462), .B(n_574), .Y(n_709) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g589 ( .A(n_463), .B(n_484), .Y(n_589) );
BUFx3_ASAP7_75t_L g614 ( .A(n_463), .Y(n_614) );
AND2x2_ASAP7_75t_L g643 ( .A(n_463), .B(n_485), .Y(n_643) );
AND3x2_ASAP7_75t_L g656 ( .A(n_463), .B(n_657), .C(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g579 ( .A(n_473), .Y(n_579) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AOI32xp33_ASAP7_75t_L g634 ( .A1(n_474), .A2(n_586), .A3(n_635), .B1(n_638), .B2(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g561 ( .A(n_475), .B(n_484), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_475), .B(n_589), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_475), .B(n_611), .Y(n_639) );
OR2x2_ASAP7_75t_L g645 ( .A(n_475), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_475), .B(n_600), .Y(n_670) );
OR2x2_ASAP7_75t_L g688 ( .A(n_475), .B(n_513), .Y(n_688) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g552 ( .A(n_476), .B(n_494), .Y(n_552) );
INVx2_ASAP7_75t_L g574 ( .A(n_476), .Y(n_574) );
OR2x2_ASAP7_75t_L g596 ( .A(n_476), .B(n_494), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_476), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_476), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_476), .B(n_551), .Y(n_657) );
INVx1_ASAP7_75t_SL g708 ( .A(n_484), .Y(n_708) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
INVx1_ASAP7_75t_SL g551 ( .A(n_485), .Y(n_551) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_485), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_485), .B(n_637), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_485), .B(n_574), .C(n_692), .Y(n_703) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_486), .A2(n_495), .B(n_501), .Y(n_494) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_486), .A2(n_505), .B(n_511), .Y(n_504) );
INVx2_ASAP7_75t_L g602 ( .A(n_494), .Y(n_602) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_494), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx1_ASAP7_75t_L g638 ( .A(n_503), .Y(n_638) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g556 ( .A(n_504), .B(n_538), .Y(n_556) );
INVx2_ASAP7_75t_L g573 ( .A(n_504), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_539), .Y(n_578) );
AND2x2_ASAP7_75t_L g593 ( .A(n_504), .B(n_526), .Y(n_593) );
AND2x2_ASAP7_75t_L g605 ( .A(n_504), .B(n_577), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_512), .B(n_621), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_512), .B(n_578), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_512), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_512), .B(n_572), .Y(n_700) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g537 ( .A(n_513), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_513), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g582 ( .A(n_513), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g608 ( .A(n_513), .B(n_538), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_513), .B(n_648), .Y(n_647) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_523), .Y(n_513) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx2_ASAP7_75t_L g533 ( .A(n_522), .Y(n_533) );
INVx1_ASAP7_75t_L g568 ( .A(n_523), .Y(n_568) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_526), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
INVx3_ASAP7_75t_SL g577 ( .A(n_526), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_526), .B(n_564), .Y(n_630) );
OR2x2_ASAP7_75t_L g640 ( .A(n_526), .B(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_526), .B(n_608), .Y(n_668) );
OR2x2_ASAP7_75t_L g698 ( .A(n_526), .B(n_538), .Y(n_698) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_539), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_526), .B(n_578), .Y(n_715) );
AND2x2_ASAP7_75t_L g722 ( .A(n_526), .B(n_604), .Y(n_722) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_535), .Y(n_526) );
INVx1_ASAP7_75t_SL g665 ( .A(n_537), .Y(n_665) );
AND2x2_ASAP7_75t_L g604 ( .A(n_538), .B(n_566), .Y(n_604) );
AND2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_573), .Y(n_618) );
AND2x2_ASAP7_75t_L g621 ( .A(n_538), .B(n_577), .Y(n_621) );
INVx1_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g560 ( .A(n_539), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_550), .A2(n_596), .B(n_720), .C(n_721), .Y(n_719) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g626 ( .A(n_551), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_552), .B(n_569), .Y(n_584) );
AND2x2_ASAP7_75t_L g610 ( .A(n_552), .B(n_611), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_557), .B(n_561), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_555), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_556), .B(n_577), .Y(n_622) );
AND2x2_ASAP7_75t_L g713 ( .A(n_556), .B(n_564), .Y(n_713) );
INVxp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g586 ( .A(n_560), .B(n_573), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_560), .B(n_571), .Y(n_587) );
OAI322xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_570), .A3(n_571), .B1(n_574), .B2(n_575), .C1(n_579), .C2(n_580), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .Y(n_563) );
AND2x2_ASAP7_75t_L g674 ( .A(n_564), .B(n_586), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_564), .B(n_638), .Y(n_720) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g617 ( .A(n_566), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g683 ( .A(n_570), .B(n_596), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_571), .B(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_572), .B(n_604), .Y(n_661) );
AND2x2_ASAP7_75t_L g607 ( .A(n_573), .B(n_577), .Y(n_607) );
AND2x2_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_574), .A2(n_653), .B(n_713), .C(n_714), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_575), .A2(n_588), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_577), .B(n_604), .Y(n_644) );
AND2x2_ASAP7_75t_L g650 ( .A(n_577), .B(n_618), .Y(n_650) );
AND2x2_ASAP7_75t_L g684 ( .A(n_577), .B(n_586), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_578), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g694 ( .A(n_578), .Y(n_694) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_582), .A2(n_610), .B1(n_612), .B2(n_617), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_585), .B1(n_587), .B2(n_588), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_584), .A2(n_620), .B1(n_622), .B2(n_623), .Y(n_619) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_589), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_699), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B(n_598), .C(n_619), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g660 ( .A(n_596), .B(n_613), .Y(n_660) );
INVx1_ASAP7_75t_L g711 ( .A(n_596), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_606), .C(n_609), .Y(n_598) );
INVx2_ASAP7_75t_SL g653 ( .A(n_597), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g718 ( .A(n_600), .Y(n_718) );
AND2x2_ASAP7_75t_L g642 ( .A(n_601), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g627 ( .A(n_602), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g689 ( .A(n_605), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_613), .B(n_715), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_617), .A2(n_629), .B(n_631), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g706 ( .A(n_620), .Y(n_706) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_624), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g637 ( .A(n_627), .Y(n_637) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_640), .B1(n_641), .B2(n_644), .C1(n_645), .C2(n_647), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g673 ( .A(n_637), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_640), .B(n_694), .Y(n_693) );
NAND2xp33_ASAP7_75t_SL g671 ( .A(n_641), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g646 ( .A(n_643), .Y(n_646) );
AND2x2_ASAP7_75t_L g710 ( .A(n_643), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g676 ( .A(n_646), .B(n_673), .Y(n_676) );
INVx1_ASAP7_75t_L g705 ( .A(n_647), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_654), .C(n_659), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_653), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g704 ( .A1(n_656), .A2(n_684), .A3(n_689), .B1(n_705), .B2(n_706), .C1(n_707), .C2(n_710), .Y(n_704) );
AND2x2_ASAP7_75t_L g691 ( .A(n_657), .B(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_664), .Y(n_659) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_671), .B2(n_674), .C(n_675), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND5xp2_ASAP7_75t_L g678 ( .A(n_679), .B(n_690), .C(n_704), .D(n_712), .E(n_716), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_684), .B(n_685), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp33_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_692), .A2(n_717), .B(n_718), .C(n_719), .Y(n_716) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_694), .A2(n_700), .A3(n_701), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_723), .Y(n_727) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
endmodule