module fake_jpeg_4886_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx12_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_1),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_18),
.C(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_8),
.B1(n_12),
.B2(n_7),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.C(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_20),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_19),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_19),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_32),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_25),
.B(n_42),
.Y(n_44)
);


endmodule