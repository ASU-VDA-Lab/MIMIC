module fake_jpeg_1977_n_219 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_219);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_11),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_54),
.Y(n_108)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_74),
.B1(n_52),
.B2(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_62),
.B1(n_53),
.B2(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_65),
.B(n_75),
.C(n_68),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_73),
.C(n_70),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_71),
.C(n_56),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_115),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_113),
.B1(n_62),
.B2(n_53),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_60),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_61),
.B(n_60),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_71),
.B(n_59),
.Y(n_125)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_83),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_73),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_129),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_96),
.B1(n_88),
.B2(n_76),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_132),
.B1(n_135),
.B2(n_106),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_80),
.B1(n_86),
.B2(n_52),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_86),
.B(n_63),
.C(n_76),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_69),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_80),
.B1(n_74),
.B2(n_67),
.Y(n_135)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_131),
.B1(n_128),
.B2(n_116),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_144),
.B1(n_63),
.B2(n_2),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_86),
.B1(n_103),
.B2(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_154),
.B1(n_35),
.B2(n_33),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_102),
.C(n_114),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_102),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_63),
.B(n_48),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_41),
.C(n_40),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_30),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_120),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_173),
.B1(n_178),
.B2(n_154),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_0),
.B(n_2),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_168),
.B(n_169),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_39),
.B(n_38),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_37),
.B(n_36),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_3),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_171),
.B1(n_176),
.B2(n_10),
.C(n_12),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_3),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_31),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_13),
.C(n_14),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_140),
.B1(n_152),
.B2(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_181),
.B1(n_185),
.B2(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_154),
.B1(n_137),
.B2(n_138),
.Y(n_185)
);

XOR2x1_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_12),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_167),
.C(n_29),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

AO221x1_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_172),
.B1(n_169),
.B2(n_166),
.C(n_174),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.C(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_159),
.C(n_175),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_19),
.C(n_20),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_204)
);

AOI321xp33_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_189),
.A3(n_190),
.B1(n_192),
.B2(n_28),
.C(n_26),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_206),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_207),
.B1(n_196),
.B2(n_195),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_25),
.C(n_18),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_197),
.C(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_208),
.C(n_21),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_210),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_213),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_212),
.C(n_209),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_213),
.C2(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_218),
.Y(n_219)
);


endmodule