module real_jpeg_4354_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_1),
.Y(n_134)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_3),
.A2(n_64),
.B1(n_186),
.B2(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_5),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_6),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_6),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_6),
.A2(n_144),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_6),
.A2(n_144),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_6),
.A2(n_144),
.B1(n_173),
.B2(n_364),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_7),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_10),
.A2(n_83),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_10),
.A2(n_83),
.B1(n_209),
.B2(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_10),
.A2(n_83),
.B1(n_258),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_11),
.A2(n_44),
.B1(n_247),
.B2(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_11),
.B(n_176),
.C(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_11),
.B(n_130),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_11),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_11),
.B(n_189),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_11),
.B(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_12),
.A2(n_257),
.B1(n_258),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_13),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_14),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_187),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_14),
.A2(n_187),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_15),
.A2(n_75),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_16),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_16),
.A2(n_94),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_16),
.A2(n_94),
.B1(n_174),
.B2(n_209),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_16),
.A2(n_51),
.B1(n_94),
.B2(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_269),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_268),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_222),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_21),
.B(n_222),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_157),
.C(n_205),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_22),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_77),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_23),
.B(n_78),
.C(n_111),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_24),
.A2(n_46),
.B1(n_47),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_24),
.Y(n_278)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_33),
.B1(n_36),
.B2(n_43),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_25),
.A2(n_35),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_28),
.Y(n_236)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_43),
.A2(n_44),
.B(n_98),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_44),
.B(n_88),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_44),
.A2(n_48),
.B(n_316),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g369 ( 
.A1(n_44),
.A2(n_370),
.B(n_371),
.Y(n_369)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_45),
.Y(n_240)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_55),
.B1(n_65),
.B2(n_69),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_48),
.A2(n_197),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_48),
.A2(n_311),
.B(n_316),
.Y(n_310)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_49),
.A2(n_70),
.B1(n_196),
.B2(n_203),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_49),
.A2(n_56),
.B1(n_283),
.B2(n_288),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_49),
.B(n_318),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_49),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_50),
.Y(n_352)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_53),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_54),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_59),
.Y(n_199)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_59),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_59),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_59),
.Y(n_319)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_59),
.Y(n_339)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_62),
.A2(n_176),
.B1(n_178),
.B2(n_180),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_63),
.Y(n_265)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_68),
.Y(n_332)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_68),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_110),
.B2(n_111),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_92),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_80),
.A2(n_88),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_87),
.B(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_90),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_99),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_100),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_100),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_139),
.B(n_149),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g228 ( 
.A1(n_112),
.A2(n_130),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_112),
.B(n_229),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_112),
.A2(n_149),
.B(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_113),
.A2(n_140),
.B1(n_156),
.B2(n_217),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_130),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_117),
.Y(n_383)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_119),
.Y(n_389)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_129),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_129),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_130),
.Y(n_156)
);

AO22x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_137),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_134),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_136),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_136),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_136),
.Y(n_306)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_156),
.A2(n_217),
.B(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_157),
.A2(n_158),
.B1(n_205),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_195),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_159),
.B(n_195),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_182),
.B1(n_188),
.B2(n_190),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_160),
.A2(n_301),
.B(n_303),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_160),
.A2(n_188),
.B1(n_323),
.B2(n_363),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_160),
.A2(n_303),
.B(n_363),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_161),
.A2(n_189),
.B1(n_191),
.B2(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_175),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_165),
.Y(n_366)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_175),
.A2(n_207),
.B(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_188),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_186),
.Y(n_324)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_189),
.B(n_208),
.Y(n_303)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_205),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_216),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_206),
.B(n_216),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g381 ( 
.A(n_209),
.Y(n_381)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_211),
.A2(n_212),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_244),
.B1(n_266),
.B2(n_267),
.Y(n_224)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_294),
.B(n_408),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_291),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_272),
.B(n_291),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.C(n_279),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_273),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_279),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.C(n_290),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_280),
.B(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_282),
.B(n_290),
.Y(n_399)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_283),
.Y(n_377)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_402),
.B(n_407),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_391),
.B(n_401),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_357),
.B(n_390),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_327),
.B(n_356),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_309),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_309),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_300),
.A2(n_304),
.B1(n_305),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_320),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_321),
.C(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_311),
.Y(n_349)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_325),
.B2(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_346),
.B(n_355),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_334),
.B(n_345),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_344),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_340),
.B(n_343),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_353),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_353),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_359),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_375),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_367),
.B2(n_368),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_367),
.C(n_375),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI32xp33_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_380),
.A3(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_379)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_379),
.Y(n_397)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_400),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_397),
.C(n_400),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_398),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_403),
.B(n_404),
.Y(n_407)
);


endmodule