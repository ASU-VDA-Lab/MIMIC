module fake_jpeg_21815_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_18),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_17),
.B1(n_25),
.B2(n_15),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_46),
.B(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_17),
.B1(n_15),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_17),
.B1(n_15),
.B2(n_30),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_56),
.B1(n_37),
.B2(n_41),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_24),
.B1(n_16),
.B2(n_27),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_21),
.B1(n_31),
.B2(n_10),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_65),
.B1(n_30),
.B2(n_38),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_42),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_19),
.B1(n_21),
.B2(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_70),
.Y(n_95)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_68),
.Y(n_93)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_63),
.B1(n_50),
.B2(n_61),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_88),
.B1(n_61),
.B2(n_31),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_41),
.B1(n_35),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_23),
.B1(n_59),
.B2(n_9),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_39),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_39),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_60),
.B1(n_42),
.B2(n_50),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_97),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_104),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_58),
.C(n_52),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_106),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_42),
.B1(n_46),
.B2(n_49),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_56),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_0),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_50),
.B1(n_61),
.B2(n_58),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_64),
.B1(n_45),
.B2(n_53),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_39),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_21),
.B1(n_33),
.B2(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_21),
.B(n_59),
.C(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_84),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_111),
.Y(n_121)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_13),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_117),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_77),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_82),
.B1(n_69),
.B2(n_72),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_127),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_83),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_98),
.B1(n_97),
.B2(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_83),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_79),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_83),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_127),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_99),
.C(n_80),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.C(n_147),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_102),
.C(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_101),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_156),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_90),
.B1(n_82),
.B2(n_110),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_148),
.B1(n_159),
.B2(n_3),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_90),
.C(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_81),
.B1(n_89),
.B2(n_23),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_81),
.C(n_23),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_160),
.C(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_133),
.Y(n_151)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_1),
.B(n_2),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_125),
.B(n_118),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_81),
.C(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_114),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_3),
.C(n_4),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_169),
.B(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_119),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

HB1xp67_ASAP7_75t_SL g170 ( 
.A(n_137),
.Y(n_170)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_171),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_115),
.B1(n_122),
.B2(n_113),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_157),
.B1(n_159),
.B2(n_150),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_113),
.B(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_180),
.C(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_131),
.B1(n_136),
.B2(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_182),
.B1(n_154),
.B2(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_131),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_131),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_163),
.B1(n_162),
.B2(n_175),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_198),
.C(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_140),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_202),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_189),
.B1(n_195),
.B2(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_152),
.B1(n_145),
.B2(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_141),
.B1(n_139),
.B2(n_8),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_14),
.C(n_7),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_14),
.C(n_7),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_14),
.C(n_7),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_166),
.B(n_6),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_209),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_165),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_212),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_171),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_178),
.B(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_216),
.B1(n_218),
.B2(n_174),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_178),
.B(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_178),
.B1(n_179),
.B2(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_167),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_187),
.B1(n_192),
.B2(n_189),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_200),
.B1(n_177),
.B2(n_168),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_183),
.B(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_202),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_197),
.Y(n_226)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_234),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_233),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_208),
.C(n_184),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_241),
.C(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_196),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_169),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_199),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_251),
.C(n_253),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_222),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_252),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_229),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_258),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_250),
.B(n_247),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_233),
.C(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_235),
.B(n_236),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_214),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_257),
.C(n_8),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_266),
.B(n_11),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_270),
.A2(n_271),
.B(n_6),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_265),
.B(n_11),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_272),
.B(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_6),
.C(n_12),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_12),
.Y(n_275)
);


endmodule