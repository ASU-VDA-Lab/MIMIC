module fake_jpeg_6161_n_58 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_15),
.B2(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_2),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_11),
.Y(n_23)
);

AND2x4_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_20),
.B(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_34),
.B(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_21),
.B1(n_9),
.B2(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_13),
.B1(n_11),
.B2(n_14),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_9),
.C(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_30),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_14),
.C(n_10),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_10),
.C(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_45),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_17),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_24),
.B(n_17),
.C(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_17),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_37),
.C(n_24),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_50),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_45),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_48),
.C(n_51),
.Y(n_53)
);

AOI31xp67_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.A3(n_44),
.B(n_6),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_47),
.C(n_44),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

AOI221xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_4),
.B1(n_7),
.B2(n_44),
.C(n_55),
.Y(n_58)
);


endmodule