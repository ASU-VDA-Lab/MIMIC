module fake_jpeg_820_n_220 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_39),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_77),
.Y(n_88)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_71),
.B1(n_72),
.B2(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_64),
.B1(n_51),
.B2(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_90),
.B1(n_54),
.B2(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_71),
.B1(n_53),
.B2(n_55),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_63),
.B(n_58),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_68),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_50),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_107),
.B1(n_82),
.B2(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_65),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_93),
.C(n_82),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_21),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_125),
.B(n_129),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_58),
.A3(n_57),
.B1(n_63),
.B2(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_127),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_75),
.B1(n_78),
.B2(n_76),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_75),
.B(n_57),
.C(n_58),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_70),
.B(n_67),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_0),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_49),
.B(n_47),
.C(n_46),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_94),
.B1(n_109),
.B2(n_2),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_145),
.B1(n_151),
.B2(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_1),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_1),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_3),
.B(n_4),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_11),
.B(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_7),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_127),
.B1(n_128),
.B2(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_132),
.B1(n_22),
.B2(n_28),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_10),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_16),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_160),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_171),
.B1(n_17),
.B2(n_18),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_170),
.Y(n_182)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_16),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_143),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_188),
.B1(n_158),
.B2(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_143),
.C(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_183),
.C(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_32),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_189),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_37),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_17),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_168),
.C(n_162),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_161),
.B1(n_164),
.B2(n_170),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_200),
.B(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_178),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_180),
.B1(n_192),
.B2(n_193),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_180),
.B1(n_163),
.B2(n_31),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_207),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_206),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_206),
.A3(n_208),
.B1(n_213),
.B2(n_41),
.C1(n_19),
.C2(n_44),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_20),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_40),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_42),
.Y(n_220)
);


endmodule