module fake_jpeg_24381_n_68 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_21),
.Y(n_27)
);

CKINVDCx9p33_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_0),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_9),
.C(n_15),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_14),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_37),
.B(n_11),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_13),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_13),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_31),
.Y(n_43)
);

XNOR2x1_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_20),
.B1(n_28),
.B2(n_1),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.C(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_17),
.B1(n_16),
.B2(n_24),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_17),
.B1(n_30),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_28),
.Y(n_59)
);

BUFx12f_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B(n_52),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_62),
.B(n_5),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_55),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_2),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_65),
.Y(n_68)
);


endmodule