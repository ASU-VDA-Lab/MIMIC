module fake_jpeg_4810_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_38),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_37),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_25),
.B1(n_30),
.B2(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_23),
.B1(n_28),
.B2(n_21),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_55),
.B1(n_15),
.B2(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_15),
.B1(n_30),
.B2(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_66),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_22),
.B(n_25),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_82),
.B(n_43),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_68),
.B1(n_49),
.B2(n_24),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_25),
.B1(n_18),
.B2(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_39),
.B1(n_27),
.B2(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_59),
.B1(n_45),
.B2(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_29),
.B1(n_19),
.B2(n_30),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_2),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_31),
.B1(n_24),
.B2(n_27),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_93),
.B1(n_96),
.B2(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_89),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_91),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_58),
.Y(n_90)
);

XOR2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_82),
.B1(n_81),
.B2(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_74),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_123),
.B1(n_90),
.B2(n_92),
.C(n_89),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_115),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_70),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_113),
.B(n_93),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_65),
.B(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_60),
.B1(n_64),
.B2(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_77),
.B1(n_49),
.B2(n_64),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_74),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_121),
.Y(n_144)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_137),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_134),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_135),
.Y(n_154)
);

XOR2x1_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_31),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_86),
.CI(n_74),
.CON(n_137),
.SN(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_116),
.B(n_109),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_45),
.C(n_27),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_145),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_124),
.B1(n_77),
.B2(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_77),
.C(n_27),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_152),
.B1(n_145),
.B2(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_112),
.B1(n_104),
.B2(n_117),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_163),
.B1(n_133),
.B2(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_104),
.B1(n_122),
.B2(n_120),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_115),
.A3(n_31),
.B1(n_66),
.B2(n_121),
.C1(n_57),
.C2(n_50),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_142),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_72),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_137),
.B1(n_128),
.B2(n_143),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_57),
.B1(n_50),
.B2(n_60),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_156),
.B1(n_162),
.B2(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_138),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_177),
.B1(n_178),
.B2(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_130),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_147),
.C(n_167),
.Y(n_186)
);

AOI321xp33_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_156),
.A3(n_152),
.B1(n_149),
.B2(n_153),
.C(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_41),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_185),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_17),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_166),
.C(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_191),
.C(n_20),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_20),
.C(n_57),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_2),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_13),
.B(n_4),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_196),
.C(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_66),
.C(n_18),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_18),
.B1(n_17),
.B2(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_6),
.C(n_7),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_181),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_208),
.Y(n_211)
);

OAI221xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_183),
.B1(n_192),
.B2(n_188),
.C(n_185),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_202),
.B(n_8),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_195),
.B(n_184),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_209),
.B(n_9),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_205),
.A2(n_194),
.B1(n_195),
.B2(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_214),
.Y(n_220)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_9),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.C(n_210),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_206),
.C(n_214),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_11),
.C(n_12),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_11),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_217),
.C(n_220),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.B(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_12),
.Y(n_227)
);


endmodule