module fake_jpeg_18737_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_25),
.B1(n_16),
.B2(n_32),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_70),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_44),
.B1(n_45),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_36),
.B1(n_23),
.B2(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_92),
.Y(n_115)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_46),
.B1(n_49),
.B2(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_41),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_56),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_98),
.Y(n_126)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_41),
.B1(n_58),
.B2(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_80),
.B1(n_65),
.B2(n_81),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_113),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_116),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_52),
.B1(n_47),
.B2(n_36),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_123),
.B1(n_66),
.B2(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_47),
.Y(n_116)
);

NOR2x1p5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_40),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_142),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_16),
.B(n_23),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_139),
.B1(n_118),
.B2(n_113),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_119),
.B1(n_101),
.B2(n_108),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_115),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_143),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_85),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_30),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_74),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_122),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_108),
.C(n_74),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_155),
.C(n_146),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_119),
.B1(n_91),
.B2(n_99),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_158),
.B1(n_177),
.B2(n_64),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_105),
.C(n_97),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_95),
.B1(n_89),
.B2(n_49),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_118),
.B1(n_100),
.B2(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_59),
.B1(n_102),
.B2(n_40),
.Y(n_200)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_178),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_174),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_82),
.B(n_68),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_173),
.B(n_124),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_169),
.B(n_171),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_94),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_57),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_59),
.B1(n_49),
.B2(n_57),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_182),
.B(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_192),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_126),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_173),
.B(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_188),
.B(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_199),
.B1(n_168),
.B2(n_176),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_131),
.Y(n_192)
);

AOI22x1_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_102),
.B1(n_137),
.B2(n_30),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_150),
.B(n_31),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_131),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_163),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_31),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_64),
.B1(n_12),
.B2(n_14),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_208),
.B1(n_176),
.B2(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_162),
.A2(n_73),
.B1(n_34),
.B2(n_17),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_206),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_11),
.B1(n_14),
.B2(n_10),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_73),
.C(n_27),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_27),
.C(n_34),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_170),
.A3(n_168),
.B1(n_151),
.B2(n_159),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_171),
.B(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_213),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_231),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_208),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_30),
.C(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_222),
.B(n_236),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_194),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_234),
.B(n_237),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_189),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_34),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_195),
.B1(n_181),
.B2(n_184),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_240),
.B1(n_226),
.B2(n_236),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_215),
.B1(n_195),
.B2(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_181),
.B1(n_183),
.B2(n_200),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_209),
.C(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_247),
.C(n_253),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_211),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_196),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_252),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_187),
.C(n_185),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_199),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_207),
.C(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_203),
.C(n_201),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_234),
.C(n_226),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_237),
.B(n_228),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_233),
.B(n_229),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_1),
.B(n_2),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_219),
.B1(n_213),
.B2(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_269),
.B1(n_251),
.B2(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_232),
.B1(n_237),
.B2(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_238),
.C(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_273),
.B1(n_276),
.B2(n_1),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_216),
.B1(n_223),
.B2(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_227),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_223),
.B1(n_20),
.B2(n_18),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_263),
.C(n_261),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_242),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

OAI22x1_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_256),
.B1(n_251),
.B2(n_3),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_8),
.B(n_9),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_289),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_290),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_9),
.B(n_11),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_269),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_266),
.B1(n_274),
.B2(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_7),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_20),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_267),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_263),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_290),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_297),
.C(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_270),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_7),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_313),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_281),
.B(n_283),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_311),
.B(n_10),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_280),
.B(n_7),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_18),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_319),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_302),
.B1(n_298),
.B2(n_296),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_9),
.B(n_18),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_322),
.B(n_31),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_17),
.B(n_31),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.B(n_315),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_309),
.B(n_307),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.A3(n_323),
.B1(n_17),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_316),
.B(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_31),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_2),
.B(n_4),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_2),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_5),
.C(n_6),
.Y(n_334)
);


endmodule