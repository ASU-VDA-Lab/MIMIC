module fake_jpeg_9637_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

OR2x2_ASAP7_75t_SL g14 ( 
.A(n_0),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_29),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_28),
.B(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_17),
.Y(n_40)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_58),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_34),
.B1(n_28),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_59),
.B1(n_19),
.B2(n_24),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_14),
.B(n_19),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_14),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_60),
.Y(n_63)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_17),
.B1(n_16),
.B2(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_19),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_72),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_60),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_57),
.C(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_78),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_81),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_50),
.C(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_86),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_67),
.B(n_16),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_44),
.C(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_74),
.B1(n_68),
.B2(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_89),
.B1(n_96),
.B2(n_23),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_82),
.B1(n_43),
.B2(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_61),
.B(n_74),
.C(n_67),
.D(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_87),
.C(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_97),
.B1(n_13),
.B2(n_15),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_17),
.B(n_20),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_96),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_75),
.C(n_69),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_107),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_75),
.B1(n_13),
.B2(n_15),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_22),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_43),
.B1(n_23),
.B2(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_105),
.B1(n_36),
.B2(n_2),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_49),
.C(n_42),
.Y(n_107)
);

OA21x2_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_94),
.B(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_113),
.B(n_100),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_112),
.C(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_111),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_36),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_5),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_106),
.B(n_102),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_1),
.B(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_5),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_109),
.B1(n_115),
.B2(n_7),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_115),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_36),
.C1(n_123),
.C2(n_124),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_130),
.B(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_132),
.Y(n_134)
);


endmodule