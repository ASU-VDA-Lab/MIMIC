module fake_netlist_5_1429_n_46 (n_8, n_10, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_46);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_46;

wire n_29;
wire n_16;
wire n_43;
wire n_12;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_42;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_38;
wire n_35;
wire n_32;
wire n_41;
wire n_11;
wire n_17;
wire n_19;
wire n_37;
wire n_26;
wire n_15;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;
wire n_39;

INVx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_11),
.B(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_19),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_29),
.Y(n_33)
);

AOI222xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_21),
.C1(n_20),
.C2(n_30),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_31),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_30),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_32),
.B(n_34),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_15),
.Y(n_39)
);

NOR2x1p5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_15),
.Y(n_40)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_22),
.B1(n_1),
.B2(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_20),
.B1(n_21),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_21),
.B1(n_12),
.B2(n_22),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_12),
.C(n_21),
.Y(n_45)
);

AOI221xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_41),
.B1(n_43),
.B2(n_12),
.C(n_5),
.Y(n_46)
);


endmodule