module fake_jpeg_23325_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_204;
wire n_81;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_49),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_21),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_29),
.B(n_32),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_57),
.B(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_33),
.B1(n_37),
.B2(n_24),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_68),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_73),
.B1(n_45),
.B2(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_30),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_29),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_78),
.B(n_82),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_34),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_55),
.C(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_34),
.B1(n_18),
.B2(n_28),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_37),
.B1(n_34),
.B2(n_24),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_97),
.B1(n_32),
.B2(n_31),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_95),
.B1(n_34),
.B2(n_73),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_79),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_97),
.B1(n_66),
.B2(n_87),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_60),
.B1(n_48),
.B2(n_44),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_115),
.B1(n_119),
.B2(n_66),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_44),
.B1(n_49),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_116),
.B1(n_117),
.B2(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

AO22x2_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_18),
.B1(n_40),
.B2(n_38),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_71),
.B1(n_35),
.B2(n_41),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_18),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_88),
.B(n_75),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_35),
.B1(n_31),
.B2(n_74),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_98),
.C(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_136),
.C(n_117),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_143),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_26),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_105),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_76),
.B(n_78),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_134),
.B(n_140),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_116),
.A3(n_99),
.B1(n_36),
.B2(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_78),
.B1(n_84),
.B2(n_35),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_84),
.B1(n_35),
.B2(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_118),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_64),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_15),
.B1(n_77),
.B2(n_96),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_19),
.B1(n_92),
.B2(n_66),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_86),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_26),
.B(n_27),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_110),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_153),
.C(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_156),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_102),
.Y(n_153)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_116),
.B1(n_102),
.B2(n_103),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_162),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_116),
.B(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_117),
.C(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_166),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_69),
.B1(n_61),
.B2(n_63),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_169),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_133),
.B1(n_144),
.B2(n_125),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_181),
.B1(n_194),
.B2(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_122),
.B1(n_121),
.B2(n_128),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_189),
.B1(n_160),
.B2(n_146),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_121),
.B1(n_130),
.B2(n_142),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_188),
.B(n_191),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_161),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_142),
.B1(n_136),
.B2(n_69),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_155),
.B1(n_63),
.B2(n_61),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_140),
.B(n_67),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_113),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_202),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_212),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_181),
.B1(n_187),
.B2(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_204),
.B1(n_210),
.B2(n_177),
.Y(n_224)
);

XNOR2x2_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_150),
.C(n_175),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_206),
.C(n_216),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_156),
.B1(n_163),
.B2(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_170),
.C(n_164),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_172),
.A2(n_162),
.B1(n_160),
.B2(n_165),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_174),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_191),
.B(n_173),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_159),
.B1(n_162),
.B2(n_167),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_153),
.C(n_155),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_162),
.B1(n_72),
.B2(n_73),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_173),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_183),
.C(n_182),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_227),
.C(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_228),
.B(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_188),
.C(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_177),
.B1(n_179),
.B2(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_196),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_185),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_202),
.C(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_81),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_10),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_205),
.C(n_211),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_21),
.C(n_22),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_26),
.B1(n_81),
.B2(n_22),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_67),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_212),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_67),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_251),
.C(n_254),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_20),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_20),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_8),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_10),
.B(n_1),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_9),
.Y(n_262)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_40),
.C(n_38),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_14),
.B1(n_25),
.B2(n_16),
.C(n_3),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_36),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_235),
.B(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_237),
.B1(n_220),
.B2(n_25),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_264),
.B1(n_249),
.B2(n_247),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_262),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_250),
.A2(n_40),
.B1(n_17),
.B2(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_267),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_38),
.B1(n_0),
.B2(n_17),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_36),
.C(n_0),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_268),
.C(n_254),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_36),
.C(n_0),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_239),
.B(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_272),
.C(n_277),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_238),
.B(n_240),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_276),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_259),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_17),
.Y(n_277)
);

OAI21x1_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_7),
.B(n_1),
.Y(n_278)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_9),
.B(n_2),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_279),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

AOI31xp67_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_263),
.A3(n_268),
.B(n_4),
.Y(n_287)
);

OAI322xp33_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_288),
.A3(n_10),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_8),
.B(n_2),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_9),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_280),
.B(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_277),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_6),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_7),
.B(n_11),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_11),
.B(n_12),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_294),
.A3(n_281),
.B1(n_293),
.B2(n_11),
.C(n_12),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_0),
.A3(n_12),
.B1(n_28),
.B2(n_296),
.C1(n_295),
.C2(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_28),
.Y(n_305)
);


endmodule