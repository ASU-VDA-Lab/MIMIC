module fake_jpeg_30694_n_199 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_24),
.B1(n_33),
.B2(n_27),
.Y(n_65)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_18),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_21),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_26),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_52),
.B1(n_53),
.B2(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_67),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_65),
.B1(n_45),
.B2(n_41),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_24),
.B1(n_32),
.B2(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_68),
.B1(n_74),
.B2(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_32),
.B1(n_17),
.B2(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_36),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_33),
.B1(n_27),
.B2(n_23),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_30),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_90),
.B1(n_95),
.B2(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_50),
.B(n_31),
.C(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_52),
.B1(n_46),
.B2(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_42),
.B1(n_44),
.B2(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_61),
.B(n_10),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_45),
.B(n_41),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_103),
.B1(n_92),
.B2(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_42),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_70),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_93),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_77),
.B1(n_75),
.B2(n_71),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_80),
.B1(n_77),
.B2(n_75),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_71),
.B1(n_79),
.B2(n_72),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_79),
.B1(n_72),
.B2(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_95),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_131),
.C(n_108),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_115),
.B1(n_118),
.B2(n_88),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_93),
.B(n_99),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_107),
.B(n_94),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_134),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_104),
.B1(n_97),
.B2(n_115),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_94),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_114),
.B1(n_86),
.B2(n_72),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_123),
.C(n_130),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_156),
.C(n_141),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_127),
.B(n_125),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_140),
.B(n_137),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_145),
.B1(n_148),
.B2(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_85),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_29),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_45),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_147),
.A3(n_140),
.B1(n_138),
.B2(n_141),
.C1(n_137),
.C2(n_87),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_164),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_169),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_11),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_84),
.B1(n_98),
.B2(n_81),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_155),
.B1(n_151),
.B2(n_89),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_159),
.C(n_153),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_41),
.C(n_29),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_84),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_9),
.B(n_2),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_163),
.B1(n_165),
.B2(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_174),
.C(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_175),
.B1(n_171),
.B2(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_165),
.B1(n_166),
.B2(n_4),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_170),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.CI(n_29),
.CON(n_192),
.SN(n_192)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_191),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_189),
.A2(n_180),
.B1(n_6),
.B2(n_5),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_188),
.B(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_192),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_186),
.B(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_192),
.C(n_190),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_29),
.Y(n_199)
);


endmodule