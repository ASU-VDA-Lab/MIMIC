module real_aes_16188_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_0), .A2(n_70), .B1(n_610), .B2(n_613), .Y(n_609) );
OAI22xp33_ASAP7_75t_SL g651 ( .A1(n_0), .A2(n_239), .B1(n_652), .B2(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_2), .A2(n_186), .B1(n_352), .B2(n_591), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1066 ( .A(n_2), .Y(n_1066) );
INVx1_ASAP7_75t_L g671 ( .A(n_3), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g707 ( .A1(n_3), .A2(n_80), .B1(n_299), .B2(n_354), .C(n_564), .Y(n_707) );
INVx1_ASAP7_75t_L g1041 ( .A(n_4), .Y(n_1041) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_4), .A2(n_132), .B1(n_482), .B2(n_648), .C(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g589 ( .A(n_5), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_6), .A2(n_14), .B1(n_860), .B2(n_863), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_6), .A2(n_14), .B1(n_892), .B2(n_895), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_7), .A2(n_173), .B1(n_349), .B2(n_352), .C(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g458 ( .A(n_7), .Y(n_458) );
INVx1_ASAP7_75t_L g263 ( .A(n_8), .Y(n_263) );
AND2x2_ASAP7_75t_L g375 ( .A(n_8), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g387 ( .A(n_8), .B(n_203), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_8), .B(n_273), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g1404 ( .A1(n_9), .A2(n_191), .B1(n_265), .B2(n_1405), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_9), .A2(n_191), .B1(n_965), .B2(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g826 ( .A(n_10), .Y(n_826) );
INVx1_ASAP7_75t_L g491 ( .A(n_11), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_11), .A2(n_226), .B1(n_296), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g1452 ( .A(n_12), .Y(n_1452) );
AOI22xp5_ASAP7_75t_L g1471 ( .A1(n_12), .A2(n_25), .B1(n_630), .B2(n_1472), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_13), .B(n_1193), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_13), .B(n_99), .Y(n_1195) );
INVx2_ASAP7_75t_L g1199 ( .A(n_13), .Y(n_1199) );
INVxp67_ASAP7_75t_SL g921 ( .A(n_15), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_15), .A2(n_150), .B1(n_538), .B2(n_955), .Y(n_954) );
XNOR2x2_ASAP7_75t_L g1034 ( .A(n_16), .B(n_1035), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1209 ( .A1(n_17), .A2(n_164), .B1(n_1200), .B2(n_1210), .Y(n_1209) );
AOI22xp5_ASAP7_75t_L g1233 ( .A1(n_18), .A2(n_151), .B1(n_1194), .B2(n_1200), .Y(n_1233) );
INVx1_ASAP7_75t_L g1154 ( .A(n_19), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_20), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_21), .A2(n_181), .B1(n_1190), .B2(n_1197), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_22), .Y(n_1097) );
XOR2x2_ASAP7_75t_L g903 ( .A(n_23), .B(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g468 ( .A(n_24), .Y(n_468) );
INVx1_ASAP7_75t_L g1461 ( .A(n_25), .Y(n_1461) );
OAI22xp5_ASAP7_75t_SL g547 ( .A1(n_26), .A2(n_548), .B1(n_549), .B2(n_657), .Y(n_547) );
INVx1_ASAP7_75t_L g657 ( .A(n_26), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_26), .A2(n_548), .B1(n_549), .B2(n_657), .Y(n_727) );
INVx1_ASAP7_75t_L g1042 ( .A(n_27), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_27), .A2(n_68), .B1(n_1062), .B2(n_1063), .C(n_1065), .Y(n_1061) );
INVx1_ASAP7_75t_L g1458 ( .A(n_28), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_28), .A2(n_155), .B1(n_482), .B2(n_630), .Y(n_1474) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_29), .A2(n_235), .B1(n_976), .B2(n_977), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_29), .A2(n_235), .B1(n_1025), .B2(n_1027), .Y(n_1024) );
AOI211xp5_ASAP7_75t_L g324 ( .A1(n_30), .A2(n_325), .B(n_327), .C(n_333), .Y(n_324) );
INVx1_ASAP7_75t_L g447 ( .A(n_30), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_31), .A2(n_59), .B1(n_296), .B2(n_301), .C(n_307), .Y(n_1052) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_31), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_32), .A2(n_107), .B1(n_1190), .B2(n_1197), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g1222 ( .A1(n_33), .A2(n_188), .B1(n_1190), .B2(n_1200), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1232 ( .A1(n_34), .A2(n_94), .B1(n_1190), .B2(n_1197), .Y(n_1232) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_35), .A2(n_471), .B(n_474), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_35), .A2(n_43), .B1(n_535), .B2(n_536), .C(n_537), .Y(n_534) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_36), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g948 ( .A1(n_36), .A2(n_39), .B1(n_518), .B2(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g1003 ( .A(n_37), .Y(n_1003) );
INVx1_ASAP7_75t_L g289 ( .A(n_38), .Y(n_289) );
INVx1_ASAP7_75t_L g306 ( .A(n_38), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_39), .A2(n_150), .B1(n_670), .B2(n_687), .C(n_691), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_40), .A2(n_137), .B1(n_392), .B2(n_487), .Y(n_689) );
INVx1_ASAP7_75t_L g711 ( .A(n_40), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_41), .A2(n_219), .B1(n_296), .B2(n_301), .C(n_307), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_41), .A2(n_115), .B1(n_416), .B2(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g493 ( .A(n_42), .Y(n_493) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_43), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g1092 ( .A(n_44), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_45), .A2(n_147), .B1(n_558), .B2(n_561), .C(n_565), .Y(n_557) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_45), .A2(n_617), .B(n_621), .C(n_632), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_46), .Y(n_1102) );
INVx1_ASAP7_75t_L g1145 ( .A(n_47), .Y(n_1145) );
INVx1_ASAP7_75t_L g1380 ( .A(n_48), .Y(n_1380) );
INVx1_ASAP7_75t_L g852 ( .A(n_49), .Y(n_852) );
INVx1_ASAP7_75t_L g1389 ( .A(n_50), .Y(n_1389) );
INVx1_ASAP7_75t_L g256 ( .A(n_51), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_52), .A2(n_194), .B1(n_313), .B2(n_320), .Y(n_1051) );
INVx1_ASAP7_75t_L g1060 ( .A(n_52), .Y(n_1060) );
INVx2_ASAP7_75t_L g292 ( .A(n_53), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_54), .A2(n_76), .B1(n_1197), .B2(n_1210), .Y(n_1223) );
XNOR2x2_ASAP7_75t_L g1371 ( .A(n_54), .B(n_1372), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_54), .A2(n_1431), .B1(n_1434), .B2(n_1479), .Y(n_1430) );
OAI221xp5_ASAP7_75t_L g1441 ( .A1(n_55), .A2(n_100), .B1(n_313), .B2(n_320), .C(n_1442), .Y(n_1441) );
INVxp67_ASAP7_75t_SL g1466 ( .A(n_55), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_56), .A2(n_202), .B1(n_863), .B2(n_1415), .Y(n_1414) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_56), .A2(n_202), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_57), .A2(n_166), .B1(n_343), .B2(n_346), .Y(n_1038) );
INVx1_ASAP7_75t_L g1058 ( .A(n_57), .Y(n_1058) );
INVx1_ASAP7_75t_L g996 ( .A(n_58), .Y(n_996) );
INVx1_ASAP7_75t_L g1075 ( .A(n_59), .Y(n_1075) );
INVx1_ASAP7_75t_L g815 ( .A(n_60), .Y(n_815) );
INVx1_ASAP7_75t_L g822 ( .A(n_61), .Y(n_822) );
INVx1_ASAP7_75t_L g814 ( .A(n_62), .Y(n_814) );
INVx1_ASAP7_75t_L g1109 ( .A(n_63), .Y(n_1109) );
AOI21xp33_ASAP7_75t_L g1149 ( .A1(n_64), .A2(n_524), .B(n_525), .Y(n_1149) );
INVxp67_ASAP7_75t_L g1168 ( .A(n_64), .Y(n_1168) );
INVx1_ASAP7_75t_L g1381 ( .A(n_65), .Y(n_1381) );
OAI211xp5_ASAP7_75t_L g846 ( .A1(n_66), .A2(n_847), .B(n_848), .C(n_851), .Y(n_846) );
INVx1_ASAP7_75t_L g890 ( .A(n_66), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_67), .A2(n_159), .B1(n_687), .B2(n_688), .C(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g712 ( .A(n_67), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_68), .A2(n_187), .B1(n_352), .B2(n_1044), .C(n_1046), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_69), .A2(n_119), .B1(n_1190), .B2(n_1197), .Y(n_1218) );
INVx1_ASAP7_75t_L g997 ( .A(n_71), .Y(n_997) );
OAI222xp33_ASAP7_75t_L g1115 ( .A1(n_72), .A2(n_116), .B1(n_214), .B2(n_317), .C1(n_334), .C2(n_1014), .Y(n_1115) );
INVx1_ASAP7_75t_L g1127 ( .A(n_72), .Y(n_1127) );
INVx1_ASAP7_75t_L g817 ( .A(n_73), .Y(n_817) );
INVx1_ASAP7_75t_L g1459 ( .A(n_74), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_74), .A2(n_205), .B1(n_392), .B2(n_487), .Y(n_1473) );
XOR2x2_ASAP7_75t_L g277 ( .A(n_75), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g989 ( .A(n_77), .Y(n_989) );
INVx1_ASAP7_75t_L g1376 ( .A(n_78), .Y(n_1376) );
OAI211xp5_ASAP7_75t_L g1406 ( .A1(n_79), .A2(n_1407), .B(n_1409), .C(n_1413), .Y(n_1406) );
INVx1_ASAP7_75t_L g1422 ( .A(n_79), .Y(n_1422) );
INVx1_ASAP7_75t_L g682 ( .A(n_80), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_81), .Y(n_1448) );
INVx1_ASAP7_75t_L g931 ( .A(n_82), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_83), .A2(n_161), .B1(n_343), .B2(n_346), .Y(n_1155) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_83), .Y(n_1157) );
AOI22xp5_ASAP7_75t_L g1227 ( .A1(n_84), .A2(n_117), .B1(n_1190), .B2(n_1197), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_85), .A2(n_115), .B1(n_343), .B2(n_346), .Y(n_342) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_85), .A2(n_368), .B(n_380), .C(n_401), .Y(n_367) );
INVx1_ASAP7_75t_L g1101 ( .A(n_86), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1118 ( .A1(n_86), .A2(n_134), .B1(n_352), .B2(n_1119), .C(n_1121), .Y(n_1118) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_87), .A2(n_246), .B1(n_429), .B2(n_645), .C(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g696 ( .A(n_87), .Y(n_696) );
INVx1_ASAP7_75t_L g341 ( .A(n_88), .Y(n_341) );
AOI22xp5_ASAP7_75t_SL g1226 ( .A1(n_89), .A2(n_236), .B1(n_1200), .B2(n_1210), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_90), .Y(n_258) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_90), .B(n_256), .Y(n_1191) );
INVx1_ASAP7_75t_L g824 ( .A(n_91), .Y(n_824) );
INVx1_ASAP7_75t_L g357 ( .A(n_92), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_93), .Y(n_775) );
OA22x2_ASAP7_75t_L g959 ( .A1(n_94), .A2(n_960), .B1(n_1031), .B2(n_1032), .Y(n_959) );
INVxp67_ASAP7_75t_L g1032 ( .A(n_94), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_95), .A2(n_141), .B1(n_761), .B2(n_763), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_95), .A2(n_96), .B1(n_488), .B2(n_675), .Y(n_798) );
INVx1_ASAP7_75t_L g776 ( .A(n_96), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_97), .A2(n_109), .B1(n_1194), .B2(n_1200), .Y(n_1206) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_98), .A2(n_162), .B1(n_480), .B2(n_482), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_98), .A2(n_148), .B1(n_325), .B2(n_522), .C(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g1193 ( .A(n_99), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_99), .B(n_1199), .Y(n_1201) );
INVx1_ASAP7_75t_L g1477 ( .A(n_100), .Y(n_1477) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_101), .A2(n_732), .B1(n_733), .B2(n_805), .Y(n_731) );
INVx1_ASAP7_75t_L g805 ( .A(n_101), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_102), .Y(n_936) );
INVx1_ASAP7_75t_L g355 ( .A(n_103), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_104), .A2(n_244), .B1(n_1190), .B2(n_1194), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_105), .A2(n_237), .B1(n_926), .B2(n_927), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_105), .A2(n_138), .B1(n_522), .B2(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g984 ( .A(n_106), .Y(n_984) );
INVx1_ASAP7_75t_L g677 ( .A(n_108), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_108), .A2(n_606), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g294 ( .A(n_110), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_110), .B(n_292), .Y(n_316) );
INVx1_ASAP7_75t_L g360 ( .A(n_110), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g964 ( .A1(n_111), .A2(n_247), .B1(n_965), .B2(n_967), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_111), .A2(n_247), .B1(n_265), .B2(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1110 ( .A(n_112), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_112), .A2(n_139), .B1(n_296), .B2(n_301), .Y(n_1116) );
INVx1_ASAP7_75t_L g1147 ( .A(n_113), .Y(n_1147) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_114), .A2(n_209), .B1(n_1190), .B2(n_1197), .Y(n_1211) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_116), .A2(n_139), .B1(n_410), .B2(n_1104), .C(n_1106), .Y(n_1103) );
INVx1_ASAP7_75t_L g1081 ( .A(n_117), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_118), .A2(n_229), .B1(n_486), .B2(n_488), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_118), .A2(n_193), .B1(n_325), .B2(n_518), .C(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_119), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_119), .Y(n_661) );
INVx1_ASAP7_75t_L g1462 ( .A(n_120), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_120), .A2(n_167), .B1(n_668), .B2(n_1476), .Y(n_1475) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_121), .A2(n_158), .B1(n_867), .B2(n_868), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_121), .A2(n_158), .B1(n_875), .B2(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g1050 ( .A(n_122), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_123), .A2(n_168), .B1(n_486), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g722 ( .A(n_123), .Y(n_722) );
INVx1_ASAP7_75t_L g818 ( .A(n_124), .Y(n_818) );
INVx1_ASAP7_75t_L g994 ( .A(n_125), .Y(n_994) );
XOR2x2_ASAP7_75t_L g1129 ( .A(n_126), .B(n_1130), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_127), .A2(n_228), .B1(n_1200), .B2(n_1217), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_128), .A2(n_129), .B1(n_313), .B2(n_320), .Y(n_312) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_128), .Y(n_402) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_129), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_130), .A2(n_192), .B1(n_486), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_130), .A2(n_229), .B1(n_518), .B2(n_520), .Y(n_517) );
AOI221xp5_ASAP7_75t_SL g686 ( .A1(n_131), .A2(n_149), .B1(n_649), .B2(n_687), .C(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g715 ( .A(n_131), .Y(n_715) );
INVx1_ASAP7_75t_L g1047 ( .A(n_132), .Y(n_1047) );
INVx1_ASAP7_75t_L g911 ( .A(n_133), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_133), .A2(n_237), .B1(n_951), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1088 ( .A(n_134), .Y(n_1088) );
BUFx3_ASAP7_75t_L g286 ( .A(n_135), .Y(n_286) );
INVx1_ASAP7_75t_L g581 ( .A(n_136), .Y(n_581) );
INVx1_ASAP7_75t_L g724 ( .A(n_137), .Y(n_724) );
INVx1_ASAP7_75t_L g913 ( .A(n_138), .Y(n_913) );
INVx1_ASAP7_75t_L g1133 ( .A(n_140), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_141), .A2(n_210), .B1(n_693), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g330 ( .A(n_142), .Y(n_330) );
INVx1_ASAP7_75t_L g1377 ( .A(n_143), .Y(n_1377) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_144), .Y(n_270) );
INVx1_ASAP7_75t_L g475 ( .A(n_145), .Y(n_475) );
OAI21xp5_ASAP7_75t_SL g933 ( .A1(n_146), .A2(n_610), .B(n_934), .Y(n_933) );
OAI221xp5_ASAP7_75t_SL g634 ( .A1(n_147), .A2(n_179), .B1(n_635), .B2(n_638), .C(n_642), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_148), .A2(n_193), .B1(n_503), .B2(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g721 ( .A(n_149), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g1140 ( .A1(n_152), .A2(n_518), .B(n_528), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g1165 ( .A(n_152), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_153), .Y(n_684) );
INVx1_ASAP7_75t_L g1386 ( .A(n_154), .Y(n_1386) );
INVx1_ASAP7_75t_L g1451 ( .A(n_155), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_156), .A2(n_220), .B1(n_591), .B2(n_592), .Y(n_590) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_156), .Y(n_646) );
INVx1_ASAP7_75t_L g751 ( .A(n_157), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g793 ( .A1(n_157), .A2(n_794), .B1(n_795), .B2(n_799), .C(n_800), .Y(n_793) );
INVx1_ASAP7_75t_L g725 ( .A(n_159), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_160), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1176 ( .A1(n_161), .A2(n_189), .B1(n_410), .B2(n_1104), .C(n_1106), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_162), .A2(n_192), .B1(n_520), .B2(n_530), .Y(n_529) );
OAI211xp5_ASAP7_75t_SL g968 ( .A1(n_163), .A2(n_880), .B(n_969), .C(n_971), .Y(n_968) );
INVx1_ASAP7_75t_L g1021 ( .A(n_163), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_165), .A2(n_171), .B1(n_1194), .B2(n_1200), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_166), .Y(n_1073) );
INVx1_ASAP7_75t_L g1456 ( .A(n_167), .Y(n_1456) );
INVx1_ASAP7_75t_L g718 ( .A(n_168), .Y(n_718) );
INVx1_ASAP7_75t_L g973 ( .A(n_169), .Y(n_973) );
INVx1_ASAP7_75t_L g1153 ( .A(n_170), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_172), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_172), .A2(n_212), .B1(n_628), .B2(n_648), .C(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g434 ( .A(n_173), .Y(n_434) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_174), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_175), .Y(n_739) );
OAI222xp33_ASAP7_75t_L g906 ( .A1(n_176), .A2(n_234), .B1(n_638), .B2(n_907), .C1(n_908), .C2(n_916), .Y(n_906) );
INVx1_ASAP7_75t_L g939 ( .A(n_176), .Y(n_939) );
INVx1_ASAP7_75t_L g1142 ( .A(n_177), .Y(n_1142) );
INVx1_ASAP7_75t_L g1444 ( .A(n_178), .Y(n_1444) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_178), .A2(n_180), .B1(n_416), .B2(n_420), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_179), .Y(n_551) );
INVx1_ASAP7_75t_L g1447 ( .A(n_180), .Y(n_1447) );
INVx1_ASAP7_75t_L g336 ( .A(n_182), .Y(n_336) );
INVx1_ASAP7_75t_L g974 ( .A(n_183), .Y(n_974) );
OAI211xp5_ASAP7_75t_SL g1016 ( .A1(n_183), .A2(n_848), .B(n_1017), .C(n_1019), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_184), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_185), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_185), .A2(n_320), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
INVx1_ASAP7_75t_L g1070 ( .A(n_186), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_187), .Y(n_1071) );
OAI221xp5_ASAP7_75t_L g1134 ( .A1(n_189), .A2(n_208), .B1(n_296), .B2(n_301), .C(n_307), .Y(n_1134) );
INVx1_ASAP7_75t_L g929 ( .A(n_190), .Y(n_929) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_194), .Y(n_1054) );
INVx1_ASAP7_75t_L g1412 ( .A(n_195), .Y(n_1412) );
OAI211xp5_ASAP7_75t_L g1419 ( .A1(n_195), .A2(n_880), .B(n_1420), .C(n_1421), .Y(n_1419) );
OAI211xp5_ASAP7_75t_L g1445 ( .A1(n_196), .A2(n_283), .B(n_307), .C(n_1446), .Y(n_1445) );
INVxp33_ASAP7_75t_SL g1468 ( .A(n_196), .Y(n_1468) );
INVx1_ASAP7_75t_L g281 ( .A(n_197), .Y(n_281) );
INVx1_ASAP7_75t_L g583 ( .A(n_198), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_198), .A2(n_220), .B1(n_628), .B2(n_630), .C(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g735 ( .A(n_199), .Y(n_735) );
INVxp67_ASAP7_75t_SL g740 ( .A(n_200), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_200), .A2(n_307), .B1(n_313), .B2(n_766), .C(n_773), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_201), .Y(n_1090) );
BUFx3_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
INVx1_ASAP7_75t_L g376 ( .A(n_203), .Y(n_376) );
INVx1_ASAP7_75t_L g1410 ( .A(n_204), .Y(n_1410) );
INVx1_ASAP7_75t_L g1454 ( .A(n_205), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_206), .A2(n_1436), .B1(n_1437), .B2(n_1478), .Y(n_1435) );
CKINVDCx5p33_ASAP7_75t_R g1436 ( .A(n_206), .Y(n_1436) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_207), .A2(n_525), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g788 ( .A(n_207), .Y(n_788) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_208), .Y(n_1178) );
INVx1_ASAP7_75t_L g772 ( .A(n_210), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_211), .Y(n_747) );
INVx1_ASAP7_75t_L g585 ( .A(n_212), .Y(n_585) );
OAI211xp5_ASAP7_75t_L g922 ( .A1(n_213), .A2(n_654), .B(n_923), .C(n_928), .Y(n_922) );
INVx1_ASAP7_75t_L g943 ( .A(n_213), .Y(n_943) );
INVx1_ASAP7_75t_L g1112 ( .A(n_214), .Y(n_1112) );
INVx2_ASAP7_75t_L g366 ( .A(n_215), .Y(n_366) );
INVx1_ASAP7_75t_L g373 ( .A(n_215), .Y(n_373) );
INVx1_ASAP7_75t_L g384 ( .A(n_215), .Y(n_384) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_216), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g1048 ( .A(n_217), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_218), .A2(n_225), .B1(n_322), .B2(n_762), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_218), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_219), .Y(n_400) );
INVx1_ASAP7_75t_L g608 ( .A(n_221), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_222), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_223), .A2(n_227), .B1(n_1197), .B2(n_1200), .Y(n_1196) );
INVx1_ASAP7_75t_L g1137 ( .A(n_224), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g1163 ( .A(n_225), .Y(n_1163) );
INVx1_ASAP7_75t_L g476 ( .A(n_226), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_230), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g1390 ( .A(n_231), .Y(n_1390) );
OAI21xp33_ASAP7_75t_SL g1439 ( .A1(n_232), .A2(n_368), .B(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1443 ( .A(n_232), .Y(n_1443) );
INVx1_ASAP7_75t_L g827 ( .A(n_233), .Y(n_827) );
INVx1_ASAP7_75t_L g941 ( .A(n_234), .Y(n_941) );
INVx1_ASAP7_75t_L g572 ( .A(n_238), .Y(n_572) );
OAI322xp33_ASAP7_75t_SL g567 ( .A1(n_239), .A2(n_568), .A3(n_575), .B1(n_578), .B2(n_584), .C1(n_593), .C2(n_598), .Y(n_567) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_240), .Y(n_464) );
INVx1_ASAP7_75t_L g855 ( .A(n_241), .Y(n_855) );
OAI211xp5_ASAP7_75t_L g879 ( .A1(n_241), .A2(n_582), .B(n_880), .C(n_882), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_242), .Y(n_669) );
INVx1_ASAP7_75t_L g993 ( .A(n_243), .Y(n_993) );
INVx1_ASAP7_75t_L g750 ( .A(n_245), .Y(n_750) );
INVx1_ASAP7_75t_L g700 ( .A(n_246), .Y(n_700) );
INVx1_ASAP7_75t_L g1384 ( .A(n_248), .Y(n_1384) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_274), .B(n_1183), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_259), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_253), .B(n_262), .Y(n_1429) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1433 ( .A(n_255), .B(n_258), .Y(n_1433) );
INVx1_ASAP7_75t_L g1481 ( .A(n_255), .Y(n_1481) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g1484 ( .A(n_258), .B(n_1481), .Y(n_1484) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g871 ( .A(n_262), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g452 ( .A(n_263), .B(n_273), .Y(n_452) );
AND2x4_ASAP7_75t_L g650 ( .A(n_263), .B(n_272), .Y(n_650) );
INVx1_ASAP7_75t_L g867 ( .A(n_264), .Y(n_867) );
AND2x4_ASAP7_75t_SL g1428 ( .A(n_264), .B(n_1429), .Y(n_1428) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
OR2x6_ASAP7_75t_L g861 ( .A(n_266), .B(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g988 ( .A(n_266), .Y(n_988) );
BUFx4f_ASAP7_75t_L g1089 ( .A(n_266), .Y(n_1089) );
INVxp67_ASAP7_75t_L g1100 ( .A(n_266), .Y(n_1100) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx4f_ASAP7_75t_L g438 ( .A(n_267), .Y(n_438) );
INVx3_ASAP7_75t_L g456 ( .A(n_267), .Y(n_456) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g378 ( .A(n_269), .Y(n_378) );
INVx2_ASAP7_75t_L g395 ( .A(n_269), .Y(n_395) );
NAND2x1_ASAP7_75t_L g399 ( .A(n_269), .B(n_270), .Y(n_399) );
AND2x2_ASAP7_75t_L g406 ( .A(n_269), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g423 ( .A(n_269), .Y(n_423) );
AND2x2_ASAP7_75t_L g484 ( .A(n_269), .B(n_270), .Y(n_484) );
INVx1_ASAP7_75t_L g379 ( .A(n_270), .Y(n_379) );
AND2x2_ASAP7_75t_L g394 ( .A(n_270), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g407 ( .A(n_270), .Y(n_407) );
BUFx2_ASAP7_75t_L g419 ( .A(n_270), .Y(n_419) );
OR2x2_ASAP7_75t_L g432 ( .A(n_270), .B(n_378), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_270), .B(n_395), .Y(n_442) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g850 ( .A(n_272), .Y(n_850) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g854 ( .A(n_273), .Y(n_854) );
AND2x4_ASAP7_75t_L g858 ( .A(n_273), .B(n_422), .Y(n_858) );
XNOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_728), .Y(n_274) );
OAI22xp33_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_277), .B1(n_459), .B2(n_460), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI211x1_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_361), .B(n_367), .C(n_408), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_323), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_295), .C(n_312), .Y(n_280) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_281), .A2(n_381), .B1(n_388), .B2(n_389), .C1(n_396), .C2(n_400), .Y(n_380) );
INVx2_ASAP7_75t_L g541 ( .A(n_282), .Y(n_541) );
AOI211xp5_ASAP7_75t_SL g1049 ( .A1(n_282), .A2(n_1050), .B(n_1051), .C(n_1052), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_282), .A2(n_532), .B1(n_1109), .B2(n_1115), .C(n_1116), .Y(n_1114) );
AOI211xp5_ASAP7_75t_L g1132 ( .A1(n_282), .A2(n_1133), .B(n_1134), .C(n_1135), .Y(n_1132) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x6_ASAP7_75t_L g613 ( .A(n_283), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g737 ( .A(n_283), .B(n_614), .Y(n_737) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
AND2x2_ASAP7_75t_L g344 ( .A(n_284), .B(n_345), .Y(n_344) );
INVx8_ASAP7_75t_L g519 ( .A(n_284), .Y(n_519) );
BUFx3_ASAP7_75t_L g762 ( .A(n_284), .Y(n_762) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AND2x4_ASAP7_75t_L g318 ( .A(n_285), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_286), .Y(n_300) );
AND2x4_ASAP7_75t_L g326 ( .A(n_286), .B(n_305), .Y(n_326) );
OR2x2_ASAP7_75t_L g335 ( .A(n_286), .B(n_288), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_286), .B(n_306), .Y(n_340) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
AND2x6_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g302 ( .A(n_290), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
AND2x4_ASAP7_75t_L g560 ( .A(n_290), .B(n_383), .Y(n_560) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_291), .B(n_360), .Y(n_359) );
NAND3x1_ASAP7_75t_L g596 ( .A(n_291), .B(n_360), .C(n_597), .Y(n_596) );
OR2x4_ASAP7_75t_L g875 ( .A(n_291), .B(n_335), .Y(n_875) );
INVx1_ASAP7_75t_L g878 ( .A(n_291), .Y(n_878) );
AND2x4_ASAP7_75t_L g881 ( .A(n_291), .B(n_326), .Y(n_881) );
OR2x6_ASAP7_75t_L g896 ( .A(n_291), .B(n_574), .Y(n_896) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
NAND2xp33_ASAP7_75t_SL g526 ( .A(n_292), .B(n_294), .Y(n_526) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_294), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_294), .Y(n_900) );
AND3x4_ASAP7_75t_L g947 ( .A(n_294), .B(n_332), .C(n_509), .Y(n_947) );
INVx4_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_297), .A2(n_302), .B1(n_750), .B2(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_297), .A2(n_302), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
AND2x2_ASAP7_75t_L g559 ( .A(n_298), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g940 ( .A(n_298), .B(n_560), .Y(n_940) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_300), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g322 ( .A(n_300), .B(n_304), .Y(n_322) );
BUFx2_ASAP7_75t_L g886 ( .A(n_300), .Y(n_886) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_302), .Y(n_514) );
INVx1_ASAP7_75t_L g564 ( .A(n_303), .Y(n_564) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g310 ( .A(n_306), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_307), .Y(n_515) );
OR2x6_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g970 ( .A(n_308), .Y(n_970) );
INVx1_ASAP7_75t_L g1402 ( .A(n_308), .Y(n_1402) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g354 ( .A(n_309), .Y(n_354) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_309), .Y(n_612) );
BUFx2_ASAP7_75t_L g889 ( .A(n_310), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_313), .Y(n_1152) );
OR2x6_ASAP7_75t_SL g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g321 ( .A(n_315), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_315), .Y(n_533) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
OR2x2_ASAP7_75t_L g556 ( .A(n_316), .B(n_453), .Y(n_556) );
INVx1_ASAP7_75t_L g571 ( .A(n_317), .Y(n_571) );
INVx3_ASAP7_75t_L g702 ( .A(n_317), .Y(n_702) );
BUFx2_ASAP7_75t_L g821 ( .A(n_317), .Y(n_821) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx8_ASAP7_75t_L g329 ( .A(n_318), .Y(n_329) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_318), .Y(n_524) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_321), .B(n_364), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g1151 ( .A1(n_321), .A2(n_1152), .B1(n_1153), .B2(n_1154), .C(n_1155), .Y(n_1151) );
BUFx3_ASAP7_75t_L g352 ( .A(n_322), .Y(n_352) );
BUFx12f_ASAP7_75t_L g520 ( .A(n_322), .Y(n_520) );
INVx5_ASAP7_75t_L g764 ( .A(n_322), .Y(n_764) );
BUFx3_ASAP7_75t_L g951 ( .A(n_322), .Y(n_951) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_342), .C(n_348), .Y(n_323) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g347 ( .A(n_326), .B(n_345), .Y(n_347) );
BUFx2_ASAP7_75t_L g539 ( .A(n_326), .Y(n_539) );
BUFx2_ASAP7_75t_L g592 ( .A(n_326), .Y(n_592) );
BUFx2_ASAP7_75t_L g748 ( .A(n_326), .Y(n_748) );
BUFx2_ASAP7_75t_L g955 ( .A(n_326), .Y(n_955) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g530 ( .A(n_328), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g1450 ( .A1(n_328), .A2(n_331), .B1(n_713), .B2(n_1451), .C(n_1452), .Y(n_1450) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_328), .A2(n_1143), .B1(n_1461), .B2(n_1462), .Y(n_1460) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g554 ( .A(n_329), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g759 ( .A(n_329), .Y(n_759) );
INVx2_ASAP7_75t_SL g774 ( .A(n_329), .Y(n_774) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_329), .Y(n_953) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_329), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_330), .A2(n_429), .B1(n_433), .B2(n_434), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_331), .A2(n_354), .B1(n_1008), .B2(n_1041), .C(n_1042), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1121 ( .A1(n_331), .A2(n_354), .B1(n_720), .B2(n_1094), .C(n_1096), .Y(n_1121) );
INVx3_ASAP7_75t_L g885 ( .A(n_332), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B1(n_337), .B2(n_341), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g356 ( .A(n_335), .Y(n_356) );
INVx2_ASAP7_75t_L g600 ( .A(n_335), .Y(n_600) );
BUFx4f_ASAP7_75t_L g710 ( .A(n_335), .Y(n_710) );
OR2x4_ASAP7_75t_L g894 ( .A(n_335), .B(n_878), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_336), .A2(n_357), .B1(n_436), .B2(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
CKINVDCx8_ASAP7_75t_R g536 ( .A(n_338), .Y(n_536) );
INVx3_ASAP7_75t_L g819 ( .A(n_338), .Y(n_819) );
INVx3_ASAP7_75t_L g1009 ( .A(n_338), .Y(n_1009) );
INVx3_ASAP7_75t_L g1125 ( .A(n_338), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g607 ( .A(n_339), .Y(n_607) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g574 ( .A(n_340), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_341), .A2(n_455), .B1(n_457), .B2(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_344), .A2(n_347), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_350), .A2(n_817), .B1(n_818), .B2(n_819), .Y(n_816) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g535 ( .A(n_351), .Y(n_535) );
AND2x4_ASAP7_75t_L g877 ( .A(n_351), .B(n_878), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_357), .C(n_358), .Y(n_353) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_354), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_354), .A2(n_710), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g768 ( .A(n_354), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g1046 ( .A1(n_354), .A2(n_358), .B1(n_710), .B2(n_1047), .C(n_1048), .Y(n_1046) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_354), .A2(n_356), .B1(n_358), .B2(n_1090), .C(n_1097), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_355), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_443) );
INVx1_ASAP7_75t_L g580 ( .A(n_356), .Y(n_580) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_356), .Y(n_1395) );
OAI221xp5_ASAP7_75t_L g1457 ( .A1(n_356), .A2(n_358), .B1(n_1138), .B2(n_1458), .C(n_1459), .Y(n_1457) );
INVx3_ASAP7_75t_L g528 ( .A(n_358), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_358), .A2(n_767), .B1(n_769), .B2(n_770), .C(n_772), .Y(n_766) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g726 ( .A(n_359), .B(n_365), .Y(n_726) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g1036 ( .A1(n_362), .A2(n_1037), .B(n_1049), .C(n_1053), .Y(n_1036) );
A2O1A1Ixp33_ASAP7_75t_L g1113 ( .A1(n_362), .A2(n_1114), .B(n_1117), .C(n_1126), .Y(n_1113) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g656 ( .A(n_363), .Y(n_656) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI21xp5_ASAP7_75t_SL g664 ( .A1(n_364), .A2(n_665), .B(n_685), .Y(n_664) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g426 ( .A(n_365), .B(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_366), .B(n_387), .Y(n_414) );
INVx2_ASAP7_75t_L g509 ( .A(n_366), .Y(n_509) );
INVx1_ASAP7_75t_L g1158 ( .A(n_368), .Y(n_1158) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_369), .B(n_468), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g734 ( .A1(n_369), .A2(n_403), .B1(n_735), .B2(n_736), .C1(n_739), .C2(n_740), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_369), .B(n_1073), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_369), .B(n_1112), .Y(n_1111) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_374), .Y(n_369) );
AND2x4_ASAP7_75t_L g403 ( .A(n_370), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g614 ( .A(n_371), .Y(n_614) );
INVx1_ASAP7_75t_L g872 ( .A(n_371), .Y(n_872) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_371), .B(n_421), .Y(n_1106) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g453 ( .A(n_372), .Y(n_453) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_374), .Y(n_653) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_375), .B(n_384), .Y(n_391) );
AND2x2_ASAP7_75t_L g404 ( .A(n_375), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_375), .B(n_483), .Y(n_620) );
AND2x4_ASAP7_75t_L g637 ( .A(n_375), .B(n_405), .Y(n_637) );
AND2x4_ASAP7_75t_L g655 ( .A(n_375), .B(n_498), .Y(n_655) );
BUFx2_ASAP7_75t_L g672 ( .A(n_375), .Y(n_672) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_376), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_377), .B(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_377), .Y(n_487) );
INVx3_ASAP7_75t_L g792 ( .A(n_377), .Y(n_792) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g1059 ( .A1(n_381), .A2(n_426), .B1(n_499), .B2(n_1060), .C1(n_1061), .C2(n_1068), .Y(n_1059) );
AOI222xp33_ASAP7_75t_L g1107 ( .A1(n_381), .A2(n_389), .B1(n_396), .B2(n_1108), .C1(n_1109), .C2(n_1110), .Y(n_1107) );
AOI222xp33_ASAP7_75t_L g1177 ( .A1(n_381), .A2(n_389), .B1(n_396), .B2(n_1133), .C1(n_1154), .C2(n_1178), .Y(n_1177) );
AOI332xp33_ASAP7_75t_L g1470 ( .A1(n_381), .A2(n_499), .A3(n_784), .B1(n_1471), .B2(n_1473), .B3(n_1474), .C1(n_1475), .C2(n_1477), .Y(n_1470) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g473 ( .A(n_383), .B(n_386), .Y(n_473) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g597 ( .A(n_384), .Y(n_597) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_387), .B(n_422), .Y(n_421) );
AND2x6_ASAP7_75t_L g633 ( .A(n_387), .B(n_483), .Y(n_633) );
INVx1_ASAP7_75t_L g641 ( .A(n_387), .Y(n_641) );
AND2x2_ASAP7_75t_L g680 ( .A(n_387), .B(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_389), .A2(n_396), .B1(n_475), .B2(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g738 ( .A(n_389), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g1056 ( .A1(n_389), .A2(n_490), .B1(n_492), .B2(n_1050), .C1(n_1057), .C2(n_1058), .Y(n_1056) );
AOI21xp33_ASAP7_75t_L g1467 ( .A1(n_389), .A2(n_1468), .B(n_1469), .Y(n_1467) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g794 ( .A(n_391), .B(n_398), .Y(n_794) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g488 ( .A(n_394), .Y(n_488) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_394), .Y(n_498) );
BUFx3_ASAP7_75t_L g668 ( .A(n_394), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_396), .A2(n_409), .B(n_1075), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1464 ( .A1(n_396), .A2(n_409), .B(n_1448), .Y(n_1464) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g910 ( .A(n_398), .Y(n_910) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_398), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_398), .A2(n_787), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
BUFx2_ASAP7_75t_SL g1385 ( .A(n_398), .Y(n_1385) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_399), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g543 ( .A(n_403), .Y(n_543) );
NAND2xp33_ASAP7_75t_SL g1126 ( .A(n_403), .B(n_1127), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_403), .B(n_1153), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_403), .B(n_1466), .Y(n_1465) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_405), .Y(n_630) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g481 ( .A(n_406), .Y(n_481) );
BUFx3_ASAP7_75t_L g648 ( .A(n_406), .Y(n_648) );
AND2x4_ASAP7_75t_L g869 ( .A(n_406), .B(n_862), .Y(n_869) );
OR3x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_415), .C(n_424), .Y(n_408) );
AOI31xp33_ASAP7_75t_L g478 ( .A1(n_409), .A2(n_426), .A3(n_479), .B(n_485), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g781 ( .A1(n_410), .A2(n_782), .B(n_786), .Y(n_781) );
OR2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_411), .Y(n_433) );
INVx4_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
BUFx4f_ASAP7_75t_L g789 ( .A(n_411), .Y(n_789) );
BUFx4f_ASAP7_75t_L g797 ( .A(n_411), .Y(n_797) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_411), .Y(n_847) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2x2_ASAP7_75t_L g416 ( .A(n_413), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g490 ( .A(n_416), .Y(n_490) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_416), .Y(n_1105) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g640 ( .A(n_419), .Y(n_640) );
BUFx2_ASAP7_75t_L g681 ( .A(n_419), .Y(n_681) );
AND2x4_ASAP7_75t_L g853 ( .A(n_419), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g492 ( .A(n_420), .Y(n_492) );
AND2x4_ASAP7_75t_L g610 ( .A(n_420), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g683 ( .A(n_421), .Y(n_683) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI33xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_428), .A3(n_435), .B1(n_443), .B2(n_450), .B3(n_454), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g828 ( .A1(n_425), .A2(n_829), .A3(n_834), .B1(n_837), .B2(n_841), .B3(n_844), .Y(n_828) );
OAI33xp33_ASAP7_75t_L g1374 ( .A1(n_425), .A2(n_1375), .A3(n_1379), .B1(n_1382), .B2(n_1387), .B3(n_1388), .Y(n_1374) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx4_ASAP7_75t_L g785 ( .A(n_426), .Y(n_785) );
INVx2_ASAP7_75t_L g982 ( .A(n_426), .Y(n_982) );
INVx2_ASAP7_75t_L g1086 ( .A(n_426), .Y(n_1086) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g796 ( .A(n_430), .Y(n_796) );
INVx4_ASAP7_75t_L g1093 ( .A(n_430), .Y(n_1093) );
INVx2_ASAP7_75t_L g1383 ( .A(n_430), .Y(n_1383) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g446 ( .A(n_432), .Y(n_446) );
BUFx3_ASAP7_75t_L g840 ( .A(n_432), .Y(n_840) );
INVx1_ASAP7_75t_L g1170 ( .A(n_432), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1172 ( .A(n_432), .Y(n_1172) );
INVx1_ASAP7_75t_L g1408 ( .A(n_433), .Y(n_1408) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g999 ( .A(n_437), .Y(n_999) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g645 ( .A(n_438), .Y(n_645) );
INVx4_ASAP7_75t_L g1067 ( .A(n_438), .Y(n_1067) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g457 ( .A(n_440), .Y(n_457) );
INVx4_ASAP7_75t_L g626 ( .A(n_440), .Y(n_626) );
INVx2_ASAP7_75t_L g920 ( .A(n_440), .Y(n_920) );
BUFx6f_ASAP7_75t_L g991 ( .A(n_440), .Y(n_991) );
INVx1_ASAP7_75t_L g1002 ( .A(n_440), .Y(n_1002) );
INVx8_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g865 ( .A(n_441), .B(n_854), .Y(n_865) );
BUFx2_ASAP7_75t_L g1166 ( .A(n_441), .Y(n_1166) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_444), .A2(n_1018), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g787 ( .A(n_446), .Y(n_787) );
INVx2_ASAP7_75t_L g912 ( .A(n_446), .Y(n_912) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g836 ( .A(n_449), .Y(n_836) );
OAI33xp33_ASAP7_75t_L g1085 ( .A1(n_450), .A2(n_1086), .A3(n_1087), .B1(n_1091), .B2(n_1095), .B3(n_1098), .Y(n_1085) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g1175 ( .A(n_451), .Y(n_1175) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x4_ASAP7_75t_L g499 ( .A(n_452), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g631 ( .A(n_452), .Y(n_631) );
INVx4_ASAP7_75t_L g691 ( .A(n_452), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_452), .B(n_500), .Y(n_843) );
INVx1_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
OR2x2_ASAP7_75t_L g577 ( .A(n_453), .B(n_526), .Y(n_577) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_453), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1388 ( .A1(n_455), .A2(n_1378), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g623 ( .A(n_456), .Y(n_623) );
BUFx3_ASAP7_75t_L g832 ( .A(n_456), .Y(n_832) );
BUFx6f_ASAP7_75t_L g1164 ( .A(n_456), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_457), .A2(n_987), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_457), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_457), .A2(n_1099), .B1(n_1101), .B2(n_1102), .Y(n_1098) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_546), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI21x1_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B(n_545), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_464), .B(n_467), .C(n_469), .D(n_508), .Y(n_545) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .C(n_508), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_468), .A2(n_493), .B1(n_538), .B2(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g605 ( .A(n_473), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_473), .B(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_475), .A2(n_532), .B1(n_534), .B2(n_540), .Y(n_531) );
NAND3xp33_ASAP7_75t_SL g477 ( .A(n_478), .B(n_489), .C(n_494), .Y(n_477) );
INVx2_ASAP7_75t_L g504 ( .A(n_480), .Y(n_504) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g629 ( .A(n_483), .Y(n_629) );
BUFx3_ASAP7_75t_L g670 ( .A(n_483), .Y(n_670) );
BUFx3_ASAP7_75t_L g688 ( .A(n_483), .Y(n_688) );
AND2x2_ASAP7_75t_L g849 ( .A(n_483), .B(n_850), .Y(n_849) );
BUFx3_ASAP7_75t_L g1472 ( .A(n_483), .Y(n_1472) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g507 ( .A(n_484), .Y(n_507) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g676 ( .A(n_487), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_490), .A2(n_492), .B1(n_747), .B2(n_750), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .C(n_502), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g693 ( .A(n_498), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_499), .Y(n_799) );
INVx2_ASAP7_75t_L g1387 ( .A(n_499), .Y(n_1387) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g687 ( .A(n_504), .Y(n_687) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_510), .B1(n_542), .B2(n_544), .Y(n_508) );
INVx1_ASAP7_75t_L g779 ( .A(n_509), .Y(n_779) );
INVx2_ASAP7_75t_SL g932 ( .A(n_509), .Y(n_932) );
OAI31xp33_ASAP7_75t_SL g1440 ( .A1(n_509), .A2(n_1441), .A3(n_1445), .B(n_1449), .Y(n_1440) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .C(n_531), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g1117 ( .A(n_515), .B(n_1118), .C(n_1122), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_521), .B1(n_527), .B2(n_529), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_518), .A2(n_560), .B(n_669), .C(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_518), .A2(n_739), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx8_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g538 ( .A(n_519), .Y(n_538) );
INVx2_ASAP7_75t_L g591 ( .A(n_519), .Y(n_591) );
INVx2_ASAP7_75t_L g698 ( .A(n_519), .Y(n_698) );
INVx8_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_523), .A2(n_715), .B1(n_716), .B2(n_718), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_523), .A2(n_536), .B1(n_1380), .B2(n_1389), .Y(n_1397) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g588 ( .A(n_524), .Y(n_588) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_524), .Y(n_1008) );
INVx2_ASAP7_75t_SL g1399 ( .A(n_524), .Y(n_1399) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g745 ( .A(n_533), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_536), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
AND2x4_ASAP7_75t_L g566 ( .A(n_539), .B(n_560), .Y(n_566) );
BUFx2_ASAP7_75t_L g949 ( .A(n_539), .Y(n_949) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_542), .B(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_658), .B1(n_659), .B2(n_727), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND3x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_603), .C(n_615), .Y(n_549) );
AOI211xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_552), .B(n_557), .C(n_567), .Y(n_550) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_554), .A2(n_697), .B1(n_929), .B2(n_931), .Y(n_934) );
AND2x4_ASAP7_75t_L g697 ( .A(n_555), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
OR2x2_ASAP7_75t_L g606 ( .A(n_556), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g611 ( .A(n_556), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g562 ( .A(n_560), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_562), .A2(n_939), .B1(n_940), .B2(n_941), .Y(n_938) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND4x1_ASAP7_75t_SL g937 ( .A(n_565), .B(n_938), .C(n_942), .D(n_945), .Y(n_937) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_572), .B2(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_572), .A2(n_589), .B1(n_622), .B2(n_624), .C(n_627), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_573), .A2(n_585), .B1(n_586), .B2(n_589), .C(n_590), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_573), .A2(n_720), .B1(n_994), .B2(n_1003), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_573), .A2(n_1381), .B1(n_1390), .B2(n_1399), .Y(n_1398) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g717 ( .A(n_574), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g1004 ( .A1(n_575), .A2(n_1005), .A3(n_1007), .B1(n_1010), .B2(n_1011), .B3(n_1013), .Y(n_1004) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI33xp33_ASAP7_75t_L g708 ( .A1(n_576), .A2(n_709), .A3(n_714), .B1(n_719), .B2(n_723), .B3(n_726), .Y(n_708) );
BUFx4f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g812 ( .A(n_577), .Y(n_812) );
BUFx4f_ASAP7_75t_L g1392 ( .A(n_577), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_579), .A2(n_984), .B1(n_996), .B2(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_581), .A2(n_624), .B1(n_643), .B2(n_646), .C(n_647), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_582), .A2(n_770), .B1(n_826), .B2(n_827), .Y(n_825) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI33xp33_ASAP7_75t_L g811 ( .A1(n_593), .A2(n_812), .A3(n_813), .B1(n_816), .B2(n_820), .B3(n_825), .Y(n_811) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI33xp33_ASAP7_75t_L g945 ( .A1(n_594), .A2(n_946), .A3(n_948), .B1(n_950), .B2(n_952), .B3(n_954), .Y(n_945) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g1012 ( .A(n_596), .Y(n_1012) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_599), .A2(n_989), .B1(n_997), .B2(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g1455 ( .A(n_600), .Y(n_1455) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g701 ( .A(n_602), .B(n_702), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_609), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_604), .B(n_936), .Y(n_935) );
INVx8_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g823 ( .A(n_607), .Y(n_823) );
INVx1_ASAP7_75t_L g1144 ( .A(n_607), .Y(n_1144) );
INVx2_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_612), .Y(n_713) );
INVx3_ASAP7_75t_L g756 ( .A(n_612), .Y(n_756) );
INVx4_ASAP7_75t_L g1139 ( .A(n_612), .Y(n_1139) );
INVx5_ASAP7_75t_L g944 ( .A(n_613), .Y(n_944) );
OAI31xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_634), .A3(n_651), .B(n_656), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g907 ( .A(n_618), .Y(n_907) );
INVx4_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_622), .A2(n_917), .B1(n_918), .B2(n_921), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_622), .A2(n_1145), .B1(n_1166), .B2(n_1174), .Y(n_1173) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_624), .A2(n_818), .B1(n_824), .B2(n_830), .Y(n_844) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_626), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_626), .A2(n_1048), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g1062 ( .A(n_629), .Y(n_1062) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g923 ( .A1(n_633), .A2(n_924), .B(n_925), .Y(n_923) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_637), .Y(n_930) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_SL g1375 ( .A1(n_645), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1375) );
INVx1_ASAP7_75t_L g1064 ( .A(n_648), .Y(n_1064) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g915 ( .A(n_650), .Y(n_915) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_653), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_694), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_672), .B(n_673), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_667) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_668), .Y(n_927) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_670), .A2(n_675), .B(n_677), .C(n_678), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_679), .Y(n_673) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_684), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_699), .C(n_704), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx2_ASAP7_75t_L g720 ( .A(n_702), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_708), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g771 ( .A(n_710), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g813 ( .A1(n_713), .A2(n_770), .B1(n_814), .B2(n_815), .Y(n_813) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_713), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_716), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_1077), .B1(n_1181), .B2(n_1182), .Y(n_728) );
INVx1_ASAP7_75t_L g1181 ( .A(n_729), .Y(n_1181) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_806), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_741), .C(n_780), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
OAI21xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_765), .B(n_777), .Y(n_741) );
OAI211xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B(n_749), .C(n_752), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_757), .C(n_760), .Y(n_752) );
OAI221xp5_ASAP7_75t_L g795 ( .A1(n_753), .A2(n_769), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_795) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g1014 ( .A(n_756), .Y(n_1014) );
INVx3_ASAP7_75t_L g1148 ( .A(n_756), .Y(n_1148) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_759), .A2(n_1092), .B1(n_1102), .B2(n_1125), .Y(n_1124) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g1120 ( .A(n_762), .Y(n_1120) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g1396 ( .A(n_768), .Y(n_1396) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_775), .A2(n_787), .B1(n_788), .B2(n_789), .C(n_790), .Y(n_786) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
A2O1A1Ixp33_ASAP7_75t_SL g1131 ( .A1(n_778), .A2(n_1132), .B(n_1151), .C(n_1156), .Y(n_1131) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_793), .C(n_801), .Y(n_780) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_787), .A2(n_817), .B1(n_822), .B2(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g926 ( .A(n_792), .Y(n_926) );
INVx2_ASAP7_75t_SL g1476 ( .A(n_792), .Y(n_1476) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_796), .A2(n_847), .B1(n_993), .B2(n_994), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_796), .A2(n_909), .B1(n_996), .B2(n_997), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_797), .A2(n_815), .B1(n_827), .B2(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AO22x2_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_956), .B1(n_957), .B2(n_1076), .Y(n_806) );
INVx1_ASAP7_75t_L g1076 ( .A(n_807), .Y(n_1076) );
XNOR2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_903), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_845), .C(n_873), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_828), .Y(n_810) );
OAI22xp5_ASAP7_75t_SL g829 ( .A1(n_814), .A2(n_826), .B1(n_830), .B2(n_833), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_820) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_836), .A2(n_1092), .B1(n_1093), .B2(n_1094), .Y(n_1091) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI33xp33_ASAP7_75t_L g980 ( .A1(n_841), .A2(n_981), .A3(n_983), .B1(n_992), .B2(n_995), .B3(n_998), .Y(n_980) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OAI31xp33_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_859), .A3(n_866), .B(n_870), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_847), .A2(n_1137), .B1(n_1147), .B2(n_1172), .Y(n_1171) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1413 ( .A(n_849), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_855), .B2(n_856), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_852), .A2(n_883), .B1(n_887), .B2(n_890), .Y(n_882) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_853), .Y(n_1020) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g1411 ( .A(n_857), .Y(n_1411) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g1023 ( .A(n_858), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1026 ( .A(n_861), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_861), .Y(n_1415) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_865), .Y(n_1028) );
INVx3_ASAP7_75t_SL g868 ( .A(n_869), .Y(n_868) );
CKINVDCx16_ASAP7_75t_R g1030 ( .A(n_869), .Y(n_1030) );
INVx4_ASAP7_75t_L g1405 ( .A(n_869), .Y(n_1405) );
OAI31xp33_ASAP7_75t_L g1015 ( .A1(n_870), .A2(n_1016), .A3(n_1024), .B(n_1029), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1403 ( .A1(n_870), .A2(n_1404), .A3(n_1406), .B(n_1414), .Y(n_1403) );
BUFx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OAI31xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_879), .A3(n_891), .B(n_897), .Y(n_873) );
INVx2_ASAP7_75t_SL g966 ( .A(n_875), .Y(n_966) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g967 ( .A(n_877), .Y(n_967) );
INVx1_ASAP7_75t_L g1418 ( .A(n_877), .Y(n_1418) );
CKINVDCx8_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
BUFx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx3_ASAP7_75t_L g972 ( .A(n_884), .Y(n_972) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
AND2x4_ASAP7_75t_L g888 ( .A(n_885), .B(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_887), .A2(n_972), .B1(n_973), .B2(n_974), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_887), .A2(n_972), .B1(n_1410), .B2(n_1422), .Y(n_1421) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
BUFx2_ASAP7_75t_L g976 ( .A(n_894), .Y(n_976) );
BUFx3_ASAP7_75t_L g1424 ( .A(n_894), .Y(n_1424) );
BUFx3_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g978 ( .A(n_896), .Y(n_978) );
INVx1_ASAP7_75t_L g1426 ( .A(n_896), .Y(n_1426) );
OAI31xp33_ASAP7_75t_L g1416 ( .A1(n_897), .A2(n_1417), .A3(n_1419), .B(n_1423), .Y(n_1416) );
BUFx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AND2x2_ASAP7_75t_SL g898 ( .A(n_899), .B(n_901), .Y(n_898) );
AND2x4_ASAP7_75t_L g962 ( .A(n_899), .B(n_901), .Y(n_962) );
INVx1_ASAP7_75t_SL g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND3x1_ASAP7_75t_L g904 ( .A(n_905), .B(n_935), .C(n_937), .Y(n_904) );
O2A1O1Ixp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_922), .B(n_932), .C(n_933), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_911), .B1(n_912), .B2(n_913), .C(n_914), .Y(n_908) );
INVx5_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx6f_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
BUFx3_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .B1(n_1033), .B2(n_1034), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g1031 ( .A(n_960), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_963), .B(n_979), .C(n_1015), .Y(n_960) );
CKINVDCx14_ASAP7_75t_R g961 ( .A(n_962), .Y(n_961) );
NOR3xp33_ASAP7_75t_SL g963 ( .A(n_964), .B(n_968), .C(n_975), .Y(n_963) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_973), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1019) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_1004), .Y(n_979) );
BUFx6f_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_985), .B1(n_989), .B2(n_990), .Y(n_983) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx5_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx6_ASAP7_75t_L g1378 ( .A(n_991), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_993), .A2(n_1000), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1000), .B1(n_1001), .B2(n_1003), .Y(n_998) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
OAI33xp33_ASAP7_75t_L g1391 ( .A1(n_1011), .A2(n_1392), .A3(n_1393), .B1(n_1397), .B2(n_1398), .B3(n_1400), .Y(n_1391) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_1018), .A2(n_1142), .B1(n_1168), .B2(n_1169), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_1020), .A2(n_1410), .B1(n_1411), .B2(n_1412), .Y(n_1409) );
INVx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1055), .Y(n_1035) );
NOR3xp33_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .C(n_1043), .Y(n_1037) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_1045), .A2(n_1142), .B1(n_1143), .B2(n_1145), .Y(n_1141) );
NAND4xp25_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1059), .C(n_1072), .D(n_1074), .Y(n_1055) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1077), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1079), .B1(n_1128), .B2(n_1180), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
XNOR2x1_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
NOR2x1_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1113), .Y(n_1082) );
NAND3xp33_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1107), .C(n_1111), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1103), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1161 ( .A1(n_1086), .A2(n_1162), .A3(n_1167), .B1(n_1171), .B2(n_1173), .B3(n_1175), .Y(n_1161) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_1125), .A2(n_1454), .B1(n_1455), .B2(n_1456), .Y(n_1453) );
BUFx2_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1129), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1159), .Y(n_1130) );
OAI21xp33_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1141), .B(n_1146), .Y(n_1135) );
OAI21xp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1138), .B(n_1140), .Y(n_1136) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx2_ASAP7_75t_L g1420 ( .A(n_1139), .Y(n_1420) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI211xp5_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1148), .B(n_1149), .C(n_1150), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1158), .Y(n_1156) );
NAND3xp33_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1177), .C(n_1179), .Y(n_1159) );
NOR2xp33_ASAP7_75t_SL g1160 ( .A(n_1161), .B(n_1176), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1162 ( .A1(n_1163), .A2(n_1164), .B1(n_1165), .B2(n_1166), .Y(n_1162) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1368), .B1(n_1370), .B2(n_1427), .C(n_1430), .Y(n_1183) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1307), .C(n_1344), .Y(n_1184) );
AOI32xp33_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1273), .A3(n_1292), .B1(n_1296), .B2(n_1306), .Y(n_1185) );
AOI211xp5_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1202), .B(n_1237), .C(n_1261), .Y(n_1186) );
OAI311xp33_ASAP7_75t_L g1237 ( .A1(n_1187), .A2(n_1238), .A3(n_1243), .B1(n_1244), .C1(n_1256), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1187), .B(n_1208), .Y(n_1305) );
AOI21xp33_ASAP7_75t_L g1340 ( .A1(n_1187), .A2(n_1341), .B(n_1343), .Y(n_1340) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1187), .B(n_1204), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1187), .B(n_1231), .Y(n_1366) );
INVx3_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_1188), .B(n_1246), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1188), .B(n_1208), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1188), .B(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1188), .B(n_1242), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1188), .B(n_1257), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1188), .B(n_1272), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1188), .B(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1188), .B(n_1306), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1188), .B(n_1208), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1188), .B(n_1228), .Y(n_1357) );
AND2x4_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1196), .Y(n_1188) );
AND2x6_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1191), .B(n_1195), .Y(n_1194) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_1191), .B(n_1198), .Y(n_1197) );
AND2x6_ASAP7_75t_L g1200 ( .A(n_1191), .B(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1191), .B(n_1195), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1191), .B(n_1195), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1191), .B(n_1198), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1193), .B(n_1199), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1482 ( .A(n_1198), .Y(n_1482) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_1203), .A2(n_1212), .B1(n_1228), .B2(n_1230), .Y(n_1202) );
A2O1A1Ixp33_ASAP7_75t_L g1288 ( .A1(n_1203), .A2(n_1231), .B(n_1289), .C(n_1290), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1203), .B(n_1263), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1203), .B(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1208), .Y(n_1204) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1205), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1205), .B(n_1208), .Y(n_1242) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1205), .Y(n_1247) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1205), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1208), .B(n_1247), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1208), .B(n_1300), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1211), .Y(n_1208) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1209), .B(n_1211), .Y(n_1264) );
AOI31xp33_ASAP7_75t_L g1314 ( .A1(n_1212), .A2(n_1310), .A3(n_1312), .B(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
OAI21xp5_ASAP7_75t_L g1321 ( .A1(n_1213), .A2(n_1322), .B(n_1324), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1219), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1214), .B(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1214), .B(n_1236), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1214), .B(n_1283), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1214), .B(n_1291), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1214), .B(n_1313), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_1215), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1215), .B(n_1236), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1248 ( .A(n_1215), .B(n_1221), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1215), .B(n_1220), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1215), .B(n_1231), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1215), .B(n_1291), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1215), .B(n_1231), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1218), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1216), .B(n_1218), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1219), .B(n_1240), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1219), .B(n_1277), .Y(n_1302) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1219), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1224), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1221), .B(n_1224), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1221), .B(n_1224), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1221), .B(n_1225), .Y(n_1291) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1221), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1224), .Y(n_1236) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1225), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1228), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1228), .B(n_1332), .Y(n_1342) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1234), .Y(n_1230) );
INVx3_ASAP7_75t_L g1241 ( .A(n_1231), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1231), .B(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1231), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1233), .Y(n_1231) );
OAI332xp33_ASAP7_75t_L g1359 ( .A1(n_1234), .A2(n_1275), .A3(n_1338), .B1(n_1360), .B2(n_1363), .B3(n_1364), .C1(n_1365), .C2(n_1367), .Y(n_1359) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1235), .B(n_1240), .Y(n_1323) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1242), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1240), .B(n_1270), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1240), .B(n_1248), .Y(n_1346) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1241), .B(n_1260), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1241), .B(n_1271), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1241), .B(n_1302), .Y(n_1358) );
CKINVDCx14_ASAP7_75t_R g1267 ( .A(n_1242), .Y(n_1267) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1243), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1248), .B1(n_1249), .B2(n_1251), .C(n_1252), .Y(n_1244) );
CKINVDCx14_ASAP7_75t_R g1326 ( .A(n_1246), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1247), .B(n_1264), .Y(n_1336) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1334 ( .A1(n_1250), .A2(n_1262), .B1(n_1335), .B2(n_1338), .C(n_1339), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1251), .B(n_1263), .Y(n_1262) );
CKINVDCx14_ASAP7_75t_R g1367 ( .A(n_1251), .Y(n_1367) );
OAI31xp33_ASAP7_75t_L g1308 ( .A1(n_1252), .A2(n_1309), .A3(n_1314), .B(n_1317), .Y(n_1308) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1253), .Y(n_1306) );
AOI21xp33_ASAP7_75t_SL g1354 ( .A1(n_1253), .A2(n_1355), .B(n_1356), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1255), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1257), .Y(n_1270) );
A2O1A1Ixp33_ASAP7_75t_SL g1296 ( .A1(n_1257), .A2(n_1297), .B(n_1299), .C(n_1305), .Y(n_1296) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1258), .Y(n_1343) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1260), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1264), .B1(n_1265), .B2(n_1267), .C(n_1268), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1263), .B(n_1295), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_1263), .A2(n_1300), .B1(n_1301), .B2(n_1303), .Y(n_1299) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1263), .Y(n_1300) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1264), .Y(n_1272) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
AOI21xp33_ASAP7_75t_L g1309 ( .A1(n_1267), .A2(n_1310), .B(n_1312), .Y(n_1309) );
A2O1A1Ixp33_ASAP7_75t_L g1330 ( .A1(n_1267), .A2(n_1319), .B(n_1331), .C(n_1333), .Y(n_1330) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1271), .C(n_1272), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1270), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1271), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1271), .B(n_1298), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1271), .B(n_1311), .Y(n_1332) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1277), .B1(n_1278), .B2(n_1279), .C(n_1280), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx2_ASAP7_75t_SL g1328 ( .A(n_1276), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1277), .B(n_1285), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1278), .B(n_1282), .Y(n_1333) );
AOI321xp33_ASAP7_75t_L g1353 ( .A1(n_1279), .A2(n_1300), .A3(n_1349), .B1(n_1354), .B2(n_1358), .C(n_1359), .Y(n_1353) );
A2O1A1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1284), .B(n_1286), .C(n_1288), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1283), .B(n_1298), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1283), .B(n_1311), .Y(n_1310) );
A2O1A1Ixp33_ASAP7_75t_L g1344 ( .A1(n_1284), .A2(n_1345), .B(n_1347), .C(n_1353), .Y(n_1344) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1290), .Y(n_1295) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1291), .Y(n_1362) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
NAND3xp33_ASAP7_75t_L g1335 ( .A(n_1300), .B(n_1336), .C(n_1337), .Y(n_1335) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OAI21xp5_ASAP7_75t_L g1339 ( .A1(n_1302), .A2(n_1322), .B(n_1328), .Y(n_1339) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
OAI21xp33_ASAP7_75t_L g1325 ( .A1(n_1304), .A2(n_1326), .B(n_1327), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1329), .Y(n_1307) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
OAI211xp5_ASAP7_75t_L g1317 ( .A1(n_1318), .A2(n_1319), .B(n_1321), .C(n_1325), .Y(n_1317) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
NOR3xp33_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1334), .C(n_1340), .Y(n_1329) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1336), .Y(n_1355) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1337), .Y(n_1364) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
CKINVDCx14_ASAP7_75t_R g1345 ( .A(n_1346), .Y(n_1345) );
AOI21xp5_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B(n_1351), .Y(n_1347) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1362), .Y(n_1360) );
BUFx2_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_1371), .Y(n_1370) );
NAND3xp33_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1403), .C(n_1416), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1391), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_1376), .A2(n_1384), .B1(n_1394), .B2(n_1396), .Y(n_1393) );
OAI22xp33_ASAP7_75t_L g1400 ( .A1(n_1377), .A2(n_1386), .B1(n_1394), .B2(n_1401), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1384), .B1(n_1385), .B2(n_1386), .Y(n_1382) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
HB1xp67_ASAP7_75t_SL g1431 ( .A(n_1432), .Y(n_1431) );
BUFx3_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVxp33_ASAP7_75t_SL g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1437), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1463), .Y(n_1438) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_1450), .A2(n_1453), .B1(n_1457), .B2(n_1460), .Y(n_1449) );
NAND4xp25_ASAP7_75t_SL g1463 ( .A(n_1464), .B(n_1465), .C(n_1467), .D(n_1470), .Y(n_1463) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
OAI21xp5_ASAP7_75t_L g1480 ( .A1(n_1481), .A2(n_1482), .B(n_1483), .Y(n_1480) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
endmodule