module fake_jpeg_3419_n_20 (n_3, n_2, n_1, n_0, n_4, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_20;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_4),
.Y(n_5)
);

INVx2_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_SL g7 ( 
.A(n_1),
.Y(n_7)
);

AND2x2_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

AOI32xp33_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NAND2x1p5_ASAP7_75t_R g13 ( 
.A(n_10),
.B(n_8),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_11),
.B1(n_7),
.B2(n_12),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_17),
.C(n_14),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_6),
.C(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_17),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_15),
.C(n_6),
.Y(n_20)
);


endmodule