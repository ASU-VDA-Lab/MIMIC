module fake_netlist_6_3411_n_1775 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1775);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1775;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_91),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_11),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_49),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_22),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_18),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_63),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_74),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_80),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_17),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_73),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

BUFx8_ASAP7_75t_SL g177 ( 
.A(n_62),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_66),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_11),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_28),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_24),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_9),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_37),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_48),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_103),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_69),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_53),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_143),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_132),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_96),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_31),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_3),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_12),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_136),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_39),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_51),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_112),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_50),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_105),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_98),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_19),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_119),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_52),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_20),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_126),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_72),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_67),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_13),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_32),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_60),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_76),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_28),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_118),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_83),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_139),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_38),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_100),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_10),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_141),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_95),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_92),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_57),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_46),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_55),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_99),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_117),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_20),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_19),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_148),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_133),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_36),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_22),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_45),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_27),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_109),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_104),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_31),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_12),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_18),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_35),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_33),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_61),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_122),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_121),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_154),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_229),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_187),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_240),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_201),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_187),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_177),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_191),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_203),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_179),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_242),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_207),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_204),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_180),
.Y(n_334)
);

BUFx2_ASAP7_75t_SL g335 ( 
.A(n_289),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_201),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_208),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_201),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_274),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_185),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_244),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_155),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_198),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_181),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_182),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_189),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_218),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_222),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_156),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_235),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_245),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_268),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_223),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_205),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_159),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_252),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_201),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_279),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_295),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_254),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_211),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_254),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_164),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_215),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_216),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_166),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_174),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_224),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_284),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_307),
.B(n_289),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_153),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_309),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_377),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

NAND2x1p5_ASAP7_75t_L g394 ( 
.A(n_316),
.B(n_174),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_336),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_153),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_347),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_174),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_306),
.Y(n_402)
);

AND3x2_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_246),
.C(n_184),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_311),
.B(n_184),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_316),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_167),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

CKINVDCx11_ASAP7_75t_R g411 ( 
.A(n_334),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_308),
.B(n_324),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_318),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_308),
.B(n_168),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_324),
.B(n_172),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_335),
.B(n_160),
.Y(n_422)
);

AND3x2_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_195),
.C(n_288),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_312),
.A2(n_200),
.B1(n_300),
.B2(n_262),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_312),
.B(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_358),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_333),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_337),
.A2(n_238),
.B1(n_275),
.B2(n_301),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_364),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_360),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_339),
.B(n_160),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_314),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_339),
.B(n_176),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_337),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_415),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_415),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_415),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_409),
.A2(n_330),
.B1(n_332),
.B2(n_315),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_365),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_409),
.A2(n_327),
.B1(n_296),
.B2(n_297),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

INVx8_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_416),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_375),
.C(n_369),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_374),
.B1(n_378),
.B2(n_367),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_433),
.B(n_367),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_219),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_442),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_442),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_448),
.A2(n_174),
.B1(n_303),
.B2(n_341),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_422),
.B(n_319),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_422),
.B(n_370),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_431),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_395),
.B(n_221),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_431),
.B(n_249),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_438),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_380),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_417),
.B(n_341),
.Y(n_497)
);

BUFx6f_ASAP7_75t_SL g498 ( 
.A(n_432),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_427),
.B(n_344),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_427),
.A2(n_342),
.B1(n_343),
.B2(n_183),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_385),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_423),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_417),
.B(n_344),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_387),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_384),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_225),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_392),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_384),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_384),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_383),
.B(n_161),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_419),
.B(n_232),
.Y(n_520)
);

NOR2x1p5_ASAP7_75t_L g521 ( 
.A(n_399),
.B(n_157),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_410),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_396),
.B(n_349),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_445),
.B(n_349),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_435),
.B(n_221),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_234),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_401),
.Y(n_533)
);

NAND3xp33_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_396),
.C(n_437),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_404),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_401),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_413),
.B(n_350),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_391),
.B(n_161),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_404),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_401),
.Y(n_541)
);

NOR2x1p5_ASAP7_75t_L g542 ( 
.A(n_432),
.B(n_157),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_401),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_411),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_393),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_391),
.B(n_302),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_393),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_393),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_419),
.B(n_241),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_423),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_381),
.B(n_448),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_391),
.B(n_162),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_390),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_437),
.A2(n_188),
.B1(n_183),
.B2(n_304),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_436),
.A2(n_210),
.B1(n_305),
.B2(n_194),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_R g558 ( 
.A(n_390),
.B(n_162),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_406),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_448),
.B(n_302),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_404),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_412),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_381),
.B(n_243),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_394),
.B(n_174),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_394),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_393),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_412),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_394),
.B(n_303),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_414),
.Y(n_573)
);

INVx8_ASAP7_75t_L g574 ( 
.A(n_381),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_406),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_314),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_414),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_436),
.B(n_163),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_428),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_381),
.B(n_248),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_381),
.A2(n_444),
.B1(n_441),
.B2(n_439),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_403),
.B(n_197),
.C(n_193),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_428),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_406),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_403),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_394),
.B(n_303),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_406),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_420),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_439),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_441),
.B(n_302),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_393),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_420),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_458),
.B(n_303),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_510),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_527),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_450),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_449),
.B(n_528),
.Y(n_604)
);

AOI22x1_ASAP7_75t_L g605 ( 
.A1(n_542),
.A2(n_231),
.B1(n_178),
.B2(n_299),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_450),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_458),
.B(n_303),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_458),
.A2(n_280),
.B1(n_271),
.B2(n_250),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_449),
.B(n_163),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_458),
.B(n_440),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_528),
.B(n_165),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_460),
.B(n_464),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_519),
.B(n_440),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_451),
.B(n_440),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_534),
.B(n_165),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_482),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_451),
.B(n_440),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_568),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_542),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_452),
.B(n_440),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_452),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_538),
.B(n_418),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_553),
.B(n_565),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_565),
.B(n_440),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_571),
.B(n_440),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_571),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_573),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_574),
.A2(n_421),
.B(n_420),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_529),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_420),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_465),
.B(n_190),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_529),
.A2(n_265),
.B1(n_171),
.B2(n_304),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_561),
.A2(n_402),
.B1(n_407),
.B2(n_418),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_579),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_486),
.B(n_169),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_579),
.B(n_420),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_522),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_529),
.B(n_169),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_585),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_535),
.B(n_421),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_554),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_592),
.B(n_421),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_466),
.B(n_411),
.C(n_351),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_592),
.A2(n_352),
.B(n_379),
.C(n_371),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_522),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_487),
.B(n_421),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_487),
.B(n_421),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_525),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_497),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_192),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_540),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_497),
.B(n_199),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_508),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_578),
.B(n_421),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_525),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_538),
.B(n_350),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_469),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_545),
.B(n_421),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_529),
.B(n_424),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_560),
.B(n_424),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_239),
.B1(n_290),
.B2(n_292),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_538),
.B(n_254),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_500),
.B(n_447),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_564),
.B(n_424),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_469),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_564),
.B(n_424),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_492),
.B(n_424),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_492),
.B(n_424),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_499),
.A2(n_171),
.B1(n_173),
.B2(n_188),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_576),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_576),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_493),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_581),
.B(n_424),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_471),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_498),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_461),
.B(n_425),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_498),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_493),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_508),
.A2(n_226),
.B1(n_228),
.B2(n_201),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_494),
.B(n_425),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_494),
.B(n_425),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_501),
.B(n_425),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_501),
.B(n_425),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_476),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_506),
.B(n_425),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_547),
.B(n_173),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_538),
.B(n_255),
.Y(n_699)
);

O2A1O1Ixp5_ASAP7_75t_L g700 ( 
.A1(n_566),
.A2(n_388),
.B(n_382),
.C(n_447),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_506),
.B(n_425),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_574),
.B(n_201),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_498),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_461),
.B(n_429),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_429),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_511),
.B(n_429),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_512),
.B(n_429),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_512),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_476),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_478),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_515),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_507),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_515),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_574),
.B(n_400),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_488),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_523),
.B(n_429),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_461),
.B(n_429),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_453),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_478),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_523),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_524),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_482),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_507),
.B(n_261),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_559),
.A2(n_362),
.B(n_351),
.C(n_352),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_454),
.A2(n_276),
.B1(n_261),
.B2(n_298),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_481),
.B(n_461),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_479),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_456),
.B(n_255),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_499),
.A2(n_278),
.B1(n_263),
.B2(n_298),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_524),
.B(n_429),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_479),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_461),
.B(n_263),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_582),
.B(n_447),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_457),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_482),
.B(n_531),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_457),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_480),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_552),
.B(n_265),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_558),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_488),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_552),
.B(n_266),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_499),
.A2(n_400),
.B1(n_170),
.B2(n_285),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_499),
.A2(n_291),
.B1(n_278),
.B2(n_276),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_459),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_467),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_480),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_584),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_584),
.B(n_266),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_514),
.B(n_382),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_520),
.B(n_382),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_584),
.B(n_533),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_580),
.A2(n_291),
.B1(n_269),
.B2(n_400),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_532),
.B(n_382),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_531),
.B(n_402),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_490),
.B(n_269),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_550),
.B(n_382),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_531),
.B(n_556),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_455),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_SL g759 ( 
.A(n_544),
.B(n_407),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_L g760 ( 
.A(n_557),
.B(n_237),
.C(n_206),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_584),
.B(n_393),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_584),
.B(n_397),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_459),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_533),
.B(n_397),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_536),
.B(n_400),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_587),
.B(n_362),
.C(n_371),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_617),
.B(n_587),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_604),
.B(n_611),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_648),
.B(n_489),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_603),
.B(n_521),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_616),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_619),
.B(n_596),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_626),
.B(n_470),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_604),
.B(n_485),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_658),
.B(n_536),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_599),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_658),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_621),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_661),
.Y(n_779)
);

OR2x2_ASAP7_75t_SL g780 ( 
.A(n_668),
.B(n_530),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_662),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_739),
.B(n_521),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_663),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_R g784 ( 
.A(n_754),
.B(n_544),
.Y(n_784)
);

NOR2x2_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_563),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_722),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_SL g787 ( 
.A(n_725),
.B(n_170),
.C(n_158),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_659),
.B(n_594),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_599),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_722),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_745),
.B(n_505),
.Y(n_791)
);

BUFx8_ASAP7_75t_L g792 ( 
.A(n_735),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_SL g793 ( 
.A(n_698),
.B(n_186),
.C(n_158),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_755),
.B(n_758),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_755),
.B(n_537),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_612),
.B(n_537),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_601),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_758),
.B(n_541),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_615),
.A2(n_596),
.B1(n_543),
.B2(n_593),
.Y(n_800)
);

AND2x4_ASAP7_75t_SL g801 ( 
.A(n_712),
.B(n_625),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_665),
.B(n_541),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_634),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_687),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_723),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_601),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_602),
.B(n_354),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_611),
.B(n_505),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_620),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_682),
.B(n_470),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_620),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_641),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_687),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_675),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_643),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_600),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_606),
.B(n_354),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_747),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_615),
.A2(n_475),
.B1(n_472),
.B2(n_473),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_683),
.B(n_472),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_473),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_664),
.A2(n_483),
.B1(n_477),
.B2(n_475),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_747),
.Y(n_823)
);

OAI221xp5_ASAP7_75t_L g824 ( 
.A1(n_681),
.A2(n_258),
.B1(n_253),
.B2(n_251),
.C(n_247),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_624),
.B(n_355),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_SL g826 ( 
.A1(n_698),
.A2(n_267),
.B1(n_264),
.B2(n_273),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_630),
.B(n_474),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_643),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_653),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_723),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_689),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_738),
.A2(n_267),
.B(n_186),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_635),
.B(n_474),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_609),
.B(n_255),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_609),
.B(n_509),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_747),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_658),
.B(n_543),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_636),
.B(n_562),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_640),
.A2(n_562),
.B(n_593),
.C(n_591),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_738),
.B(n_509),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_653),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_639),
.B(n_569),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_741),
.B(n_355),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_657),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_634),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_657),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_741),
.B(n_551),
.Y(n_848)
);

AOI21xp33_ASAP7_75t_L g849 ( 
.A1(n_671),
.A2(n_567),
.B(n_572),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_667),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_658),
.B(n_569),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_634),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_699),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_667),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_645),
.B(n_551),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_622),
.B(n_356),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_610),
.A2(n_551),
.B(n_586),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_645),
.B(n_586),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_644),
.B(n_477),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_733),
.A2(n_575),
.B1(n_591),
.B2(n_590),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_757),
.B(n_379),
.C(n_356),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_600),
.B(n_575),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_724),
.A2(n_567),
.B(n_588),
.C(n_572),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_646),
.B(n_583),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_652),
.B(n_583),
.Y(n_865)
);

NOR2x2_ASAP7_75t_L g866 ( 
.A(n_728),
.B(n_264),
.Y(n_866)
);

AO22x1_ASAP7_75t_L g867 ( 
.A1(n_640),
.A2(n_273),
.B1(n_282),
.B2(n_285),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_689),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_654),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_684),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_690),
.B(n_590),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_689),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_660),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_669),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_660),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_632),
.B(n_488),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_703),
.Y(n_877)
);

AND2x6_ASAP7_75t_SL g878 ( 
.A(n_759),
.B(n_357),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_708),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_660),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_664),
.A2(n_483),
.B1(n_495),
.B2(n_496),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_711),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_713),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_720),
.B(n_491),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_637),
.B(n_488),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_721),
.B(n_491),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_664),
.B(n_357),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_677),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_766),
.B(n_366),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_605),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_742),
.A2(n_608),
.B1(n_673),
.B2(n_685),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_729),
.B(n_586),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_760),
.B(n_488),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_703),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_743),
.B(n_589),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_685),
.A2(n_651),
.B1(n_691),
.B2(n_598),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_734),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_677),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_740),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_703),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_686),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_SL g902 ( 
.A(n_650),
.B(n_294),
.C(n_293),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_613),
.B(n_495),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_715),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_740),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_740),
.B(n_504),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_614),
.B(n_366),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_651),
.B(n_317),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_598),
.B(n_607),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_700),
.A2(n_588),
.B(n_502),
.C(n_503),
.Y(n_910)
);

BUFx6f_ASAP7_75t_SL g911 ( 
.A(n_736),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_744),
.B(n_496),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_718),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_607),
.B(n_317),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_SL g915 ( 
.A1(n_752),
.A2(n_301),
.B1(n_294),
.B2(n_293),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_749),
.B(n_589),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_763),
.B(n_321),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_618),
.B(n_504),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_686),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_750),
.B(n_589),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_666),
.B(n_696),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_623),
.B(n_504),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_696),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_709),
.B(n_502),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_709),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_710),
.Y(n_926)
);

NOR2x1_ASAP7_75t_R g927 ( 
.A(n_732),
.B(n_282),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_751),
.B(n_321),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_719),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_751),
.B(n_322),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_726),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_726),
.A2(n_287),
.B1(n_286),
.B2(n_213),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_647),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_719),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_753),
.B(n_212),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_727),
.Y(n_936)
);

BUFx8_ASAP7_75t_SL g937 ( 
.A(n_727),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_756),
.Y(n_938)
);

AOI22x1_ASAP7_75t_L g939 ( 
.A1(n_731),
.A2(n_526),
.B1(n_570),
.B2(n_462),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_627),
.A2(n_287),
.B1(n_286),
.B2(n_230),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_731),
.B(n_503),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_748),
.B(n_655),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_702),
.A2(n_546),
.B1(n_570),
.B2(n_526),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_672),
.B(n_504),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_737),
.B(n_484),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_768),
.A2(n_748),
.B1(n_702),
.B2(n_670),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_805),
.B(n_656),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_899),
.A2(n_714),
.B(n_631),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_931),
.A2(n_679),
.B1(n_692),
.B2(n_633),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_794),
.B(n_647),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_779),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_891),
.A2(n_706),
.B1(n_642),
.B2(n_649),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_899),
.A2(n_714),
.B(n_676),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_891),
.A2(n_678),
.B1(n_670),
.B2(n_628),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_774),
.A2(n_678),
.B1(n_765),
.B2(n_705),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_746),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_813),
.Y(n_957)
);

AOI21x1_ASAP7_75t_SL g958 ( 
.A1(n_890),
.A2(n_701),
.B(n_680),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_830),
.A2(n_694),
.B(n_693),
.C(n_695),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_777),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_769),
.B(n_794),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_773),
.A2(n_909),
.B1(n_843),
.B2(n_896),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_834),
.A2(n_697),
.B(n_707),
.C(n_730),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_824),
.B(n_214),
.C(n_217),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_773),
.A2(n_716),
.B1(n_746),
.B2(n_236),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_794),
.B(n_513),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_899),
.A2(n_688),
.B(n_704),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_818),
.A2(n_688),
.B(n_704),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_938),
.B(n_764),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_781),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_818),
.A2(n_717),
.B(n_765),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_783),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_813),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_777),
.B(n_761),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_808),
.A2(n_764),
.B(n_717),
.C(n_484),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_935),
.A2(n_526),
.B(n_570),
.C(n_546),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_814),
.A2(n_453),
.B(n_463),
.C(n_468),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_840),
.B(n_546),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_909),
.A2(n_233),
.B1(n_322),
.B2(n_323),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_853),
.B(n_548),
.Y(n_981)
);

AND2x2_ASAP7_75t_SL g982 ( 
.A(n_813),
.B(n_323),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_869),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_SL g984 ( 
.A(n_784),
.B(n_331),
.C(n_329),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_870),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_872),
.B(n_894),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_770),
.B(n_845),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_888),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_848),
.B(n_548),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_818),
.A2(n_836),
.B(n_823),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_778),
.B(n_328),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_861),
.A2(n_468),
.B(n_463),
.C(n_328),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_896),
.A2(n_762),
.B(n_548),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_803),
.B(n_513),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_853),
.B(n_331),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_942),
.A2(n_762),
.B(n_329),
.C(n_388),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_823),
.A2(n_595),
.B(n_549),
.Y(n_997)
);

OAI21xp33_ASAP7_75t_L g998 ( 
.A1(n_832),
.A2(n_595),
.B(n_549),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_770),
.B(n_852),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_782),
.B(n_595),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_909),
.A2(n_595),
.B1(n_549),
.B2(n_518),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_787),
.B(n_595),
.C(n_549),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_823),
.A2(n_549),
.B(n_518),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_SL g1004 ( 
.A(n_902),
.B(n_4),
.C(n_5),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_907),
.B(n_518),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_873),
.B(n_518),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_900),
.B(n_145),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_771),
.B(n_90),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_767),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_823),
.A2(n_518),
.B(n_516),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_831),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_879),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_875),
.B(n_516),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_839),
.A2(n_400),
.B(n_516),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_937),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_855),
.A2(n_513),
.B(n_516),
.C(n_397),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_831),
.Y(n_1017)
);

OA22x2_ASAP7_75t_L g1018 ( 
.A1(n_826),
.A2(n_801),
.B1(n_915),
.B2(n_847),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_907),
.B(n_516),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_788),
.B(n_513),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_835),
.A2(n_88),
.B(n_138),
.C(n_127),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_898),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_858),
.A2(n_513),
.B(n_397),
.C(n_10),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_892),
.A2(n_397),
.B(n_8),
.C(n_13),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_880),
.B(n_123),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_895),
.A2(n_400),
.B(n_115),
.C(n_107),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_887),
.B(n_397),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_867),
.A2(n_6),
.B1(n_14),
.B2(n_15),
.C(n_21),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_831),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_940),
.B(n_23),
.C(n_25),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_836),
.A2(n_397),
.B(n_400),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_887),
.B(n_94),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_877),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_856),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_882),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_807),
.B(n_93),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_780),
.B(n_29),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_807),
.B(n_89),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_877),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_816),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_817),
.B(n_86),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_901),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_836),
.B(n_79),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_883),
.A2(n_30),
.B(n_33),
.C(n_34),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_897),
.A2(n_30),
.B(n_35),
.C(n_36),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_791),
.B(n_38),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_817),
.B(n_39),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_940),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_856),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_825),
.B(n_75),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_919),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_789),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_878),
.B(n_43),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_816),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_810),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_798),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_877),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_797),
.A2(n_44),
.B(n_48),
.C(n_50),
.Y(n_1058)
);

INVx6_ASAP7_75t_L g1059 ( 
.A(n_792),
.Y(n_1059)
);

CKINVDCx10_ASAP7_75t_R g1060 ( 
.A(n_911),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_925),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_825),
.B(n_51),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_916),
.A2(n_56),
.B(n_58),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_810),
.B(n_820),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_920),
.A2(n_64),
.B(n_54),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_939),
.A2(n_857),
.B(n_924),
.Y(n_1066)
);

CKINVDCx8_ASAP7_75t_R g1067 ( 
.A(n_790),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_927),
.B(n_889),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_806),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_L g1070 ( 
.A(n_932),
.B(n_889),
.C(n_868),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_786),
.B(n_933),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_804),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_904),
.B(n_917),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_921),
.A2(n_918),
.B(n_903),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_793),
.B(n_928),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_893),
.A2(n_796),
.B(n_921),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_809),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_903),
.A2(n_772),
.B(n_876),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_933),
.B(n_913),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_849),
.A2(n_863),
.B(n_819),
.C(n_822),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_928),
.A2(n_930),
.B1(n_933),
.B2(n_923),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_849),
.A2(n_913),
.B(n_885),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_792),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_820),
.B(n_859),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_930),
.A2(n_802),
.B1(n_799),
.B2(n_914),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_821),
.A2(n_833),
.B(n_827),
.C(n_859),
.Y(n_1087)
);

O2A1O1Ixp5_ASAP7_75t_L g1088 ( 
.A1(n_837),
.A2(n_851),
.B(n_922),
.C(n_944),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_811),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_929),
.B(n_827),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1049),
.B(n_884),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1039),
.B(n_833),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1079),
.A2(n_913),
.B(n_821),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_SL g1094 ( 
.A(n_1085),
.B(n_914),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_962),
.A2(n_910),
.B(n_800),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_SL g1096 ( 
.A1(n_1064),
.A2(n_884),
.B(n_886),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1064),
.B(n_886),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1085),
.B(n_947),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_995),
.B(n_908),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1066),
.A2(n_941),
.B(n_924),
.Y(n_1100)
);

AO32x2_ASAP7_75t_L g1101 ( 
.A1(n_962),
.A2(n_1055),
.A3(n_952),
.B1(n_980),
.B2(n_965),
.Y(n_1101)
);

CKINVDCx6p67_ASAP7_75t_R g1102 ( 
.A(n_1060),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1034),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_987),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_982),
.B(n_913),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1075),
.A2(n_905),
.B(n_941),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1016),
.A2(n_865),
.A3(n_871),
.B(n_864),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1083),
.A2(n_842),
.B(n_838),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1030),
.B(n_881),
.C(n_908),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_951),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_948),
.A2(n_912),
.B(n_945),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_R g1112 ( 
.A(n_986),
.B(n_914),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_952),
.A2(n_860),
.B(n_943),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_993),
.A2(n_963),
.B(n_1081),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_987),
.B(n_908),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_973),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1087),
.A2(n_854),
.B(n_844),
.C(n_841),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_991),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_846),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_999),
.B(n_776),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1077),
.A2(n_862),
.B(n_829),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_1067),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1090),
.B(n_815),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_SL g1124 ( 
.A1(n_1046),
.A2(n_785),
.B(n_866),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_970),
.Y(n_1125)
);

AND2x6_ASAP7_75t_L g1126 ( 
.A(n_960),
.B(n_936),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_1084),
.B(n_775),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1023),
.A2(n_929),
.A3(n_934),
.B(n_926),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1014),
.A2(n_812),
.B(n_828),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_979),
.A2(n_905),
.B(n_906),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_989),
.A2(n_905),
.B(n_850),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_972),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1068),
.B(n_775),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_949),
.A2(n_775),
.B(n_1074),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_993),
.A2(n_775),
.B(n_946),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_949),
.A2(n_953),
.B(n_956),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_1073),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1001),
.A2(n_971),
.B(n_998),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1001),
.A2(n_975),
.B(n_976),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1014),
.A2(n_990),
.B(n_1088),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_961),
.B(n_983),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_985),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_1047),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1059),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_997),
.A2(n_1003),
.B(n_1010),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_959),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1070),
.A2(n_964),
.B1(n_1076),
.B2(n_1037),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1059),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1072),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_954),
.A2(n_955),
.B(n_1021),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1012),
.B(n_1082),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1048),
.A2(n_1024),
.B1(n_1028),
.B2(n_1035),
.C(n_1044),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_960),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_968),
.A2(n_1019),
.B(n_1005),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1053),
.B(n_1004),
.C(n_1009),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_977),
.Y(n_1156)
);

O2A1O1Ixp5_ASAP7_75t_L g1157 ( 
.A1(n_1065),
.A2(n_980),
.B(n_965),
.C(n_1080),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_978),
.A2(n_967),
.B(n_1031),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1020),
.A2(n_969),
.B(n_966),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_1086),
.B(n_1062),
.C(n_981),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_950),
.B(n_1089),
.Y(n_1161)
);

NAND3x1_ASAP7_75t_L g1162 ( 
.A(n_1000),
.B(n_1008),
.C(n_1018),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1072),
.B(n_1022),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_950),
.B(n_1078),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1027),
.A2(n_1013),
.B(n_1006),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_994),
.A2(n_1043),
.B(n_1069),
.Y(n_1166)
);

CKINVDCx11_ASAP7_75t_R g1167 ( 
.A(n_1015),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1045),
.B(n_1035),
.C(n_1038),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_L g1169 ( 
.A(n_957),
.B(n_1011),
.Y(n_1169)
);

O2A1O1Ixp5_ASAP7_75t_SL g1170 ( 
.A1(n_1052),
.A2(n_1056),
.B(n_1041),
.C(n_1036),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_1071),
.B(n_984),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_996),
.A2(n_992),
.B(n_1002),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1029),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_957),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_988),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1072),
.B(n_1033),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_957),
.Y(n_1177)
);

INVx3_ASAP7_75t_SL g1178 ( 
.A(n_1011),
.Y(n_1178)
);

AO22x2_ASAP7_75t_L g1179 ( 
.A1(n_1050),
.A2(n_1032),
.B1(n_1018),
.B2(n_1025),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1040),
.B(n_1054),
.Y(n_1180)
);

AOI221x1_ASAP7_75t_L g1181 ( 
.A1(n_1025),
.A2(n_1026),
.B1(n_1040),
.B2(n_1061),
.C(n_1042),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_974),
.A2(n_1051),
.B(n_1007),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1017),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1017),
.B(n_1057),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1057),
.A2(n_1066),
.B(n_958),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1057),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_957),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1079),
.A2(n_1075),
.B(n_1085),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1064),
.B(n_768),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1016),
.A2(n_1079),
.B(n_1066),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_617),
.B(n_648),
.C(n_805),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1079),
.A2(n_1075),
.B(n_1085),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_SL g1194 ( 
.A1(n_962),
.A2(n_931),
.B(n_658),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_957),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_999),
.B(n_987),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_951),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_951),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_995),
.B(n_604),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1066),
.A2(n_958),
.B(n_948),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1049),
.B(n_604),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1064),
.B(n_768),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_951),
.Y(n_1205)
);

AO32x2_ASAP7_75t_L g1206 ( 
.A1(n_962),
.A2(n_1055),
.A3(n_952),
.B1(n_980),
.B2(n_965),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_951),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1064),
.B(n_768),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1064),
.B(n_768),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1087),
.A2(n_769),
.B(n_615),
.C(n_612),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_SL g1211 ( 
.A(n_973),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_951),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_957),
.Y(n_1213)
);

AOI221x1_ASAP7_75t_L g1214 ( 
.A1(n_1024),
.A2(n_962),
.B1(n_1023),
.B2(n_1065),
.C(n_1016),
.Y(n_1214)
);

AOI21xp33_ASAP7_75t_L g1215 ( 
.A1(n_962),
.A2(n_768),
.B(n_615),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1049),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1079),
.A2(n_1075),
.B(n_1085),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_SL g1218 ( 
.A(n_1067),
.B(n_722),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1064),
.B(n_768),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_SL g1220 ( 
.A(n_1085),
.B(n_777),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1064),
.A2(n_1085),
.B1(n_962),
.B2(n_931),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_951),
.Y(n_1222)
);

AOI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_962),
.A2(n_768),
.B(n_615),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1064),
.A2(n_1085),
.B1(n_962),
.B2(n_931),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1090),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1087),
.A2(n_769),
.B(n_615),
.C(n_612),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1083),
.A2(n_1077),
.B(n_1079),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_951),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1039),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1066),
.A2(n_958),
.B(n_948),
.Y(n_1232)
);

AND3x4_ASAP7_75t_L g1233 ( 
.A(n_987),
.B(n_650),
.C(n_1070),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1079),
.Y(n_1234)
);

INVx8_ASAP7_75t_L g1235 ( 
.A(n_1144),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1204),
.B(n_1190),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1214),
.A2(n_1136),
.A3(n_1139),
.B(n_1193),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1100),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1229),
.A2(n_1145),
.B(n_1111),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1147),
.A2(n_1209),
.B1(n_1219),
.B2(n_1208),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1233),
.A2(n_1155),
.B1(n_1200),
.B2(n_1099),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1210),
.B(n_1228),
.C(n_1223),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1207),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1230),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1110),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1188),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1227),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1125),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1204),
.B(n_1098),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1217),
.A2(n_1194),
.B(n_1226),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1118),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1167),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1215),
.A2(n_1223),
.B(n_1192),
.C(n_1168),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1103),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1189),
.A2(n_1234),
.B(n_1226),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1189),
.A2(n_1234),
.B(n_1196),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1216),
.B(n_1163),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1097),
.A2(n_1215),
.B(n_1170),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1157),
.A2(n_1160),
.B(n_1134),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1202),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_1180),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1106),
.A2(n_1154),
.B(n_1093),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1132),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1137),
.B(n_1122),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1094),
.A2(n_1096),
.B(n_1220),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1138),
.A2(n_1225),
.A3(n_1221),
.B(n_1181),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1142),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1221),
.A2(n_1225),
.B(n_1159),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1149),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1102),
.B(n_1148),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_L g1272 ( 
.A(n_1203),
.B(n_1092),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1198),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1179),
.A2(n_1109),
.B1(n_1143),
.B2(n_1171),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1150),
.A2(n_1196),
.B(n_1224),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1114),
.A2(n_1202),
.B(n_1224),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1199),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1118),
.B(n_1123),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1143),
.B(n_1091),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1095),
.A2(n_1135),
.B(n_1113),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1129),
.A2(n_1121),
.B(n_1095),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1135),
.A2(n_1113),
.B(n_1108),
.Y(n_1282)
);

OAI221xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1109),
.B2(n_1151),
.C(n_1124),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1108),
.A2(n_1166),
.B(n_1191),
.Y(n_1284)
);

AO21x2_ASAP7_75t_L g1285 ( 
.A1(n_1172),
.A2(n_1117),
.B(n_1131),
.Y(n_1285)
);

AOI221xp5_ASAP7_75t_L g1286 ( 
.A1(n_1152),
.A2(n_1212),
.B1(n_1222),
.B2(n_1141),
.C(n_1172),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1174),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1165),
.A2(n_1130),
.B(n_1182),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1174),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1191),
.A2(n_1105),
.B(n_1161),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1153),
.A2(n_1164),
.B(n_1175),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1101),
.A2(n_1206),
.B(n_1107),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1101),
.A2(n_1206),
.B(n_1107),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1156),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1153),
.A2(n_1162),
.B(n_1133),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1197),
.B(n_1104),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1107),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1126),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1197),
.B(n_1119),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1169),
.A2(n_1127),
.B(n_1092),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1092),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1187),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1206),
.A2(n_1128),
.B(n_1120),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1184),
.A2(n_1186),
.B(n_1128),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1218),
.B(n_1176),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1126),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1177),
.A2(n_1195),
.A3(n_1183),
.B(n_1126),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1176),
.B(n_1187),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1187),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1213),
.B(n_1177),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1116),
.Y(n_1311)
);

INVx3_ASAP7_75t_SL g1312 ( 
.A(n_1178),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1213),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1213),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1183),
.B(n_1195),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1211),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1173),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1127),
.A2(n_1112),
.B(n_1211),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1231),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1210),
.A2(n_1228),
.B(n_648),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1322)
);

INVxp33_ASAP7_75t_L g1323 ( 
.A(n_1200),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1214),
.A2(n_1136),
.A3(n_1139),
.B(n_1188),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1205),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1234),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1200),
.B(n_306),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1234),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1204),
.B(n_1190),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1174),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1103),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1166),
.B(n_1140),
.Y(n_1336)
);

CKINVDCx16_ASAP7_75t_R g1337 ( 
.A(n_1122),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1094),
.A2(n_1096),
.B(n_1220),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1205),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1205),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1155),
.A2(n_1168),
.B1(n_964),
.B2(n_615),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1098),
.A2(n_1227),
.B1(n_648),
.B2(n_617),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1210),
.A2(n_1228),
.B(n_648),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1205),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1205),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1118),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1234),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1115),
.B(n_1180),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1118),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1174),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1174),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1227),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1200),
.B(n_1098),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1200),
.B(n_1098),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1098),
.A2(n_1227),
.B1(n_648),
.B2(n_617),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1234),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_SL g1361 ( 
.A1(n_1210),
.A2(n_1228),
.B(n_1024),
.C(n_1081),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1200),
.B(n_1098),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1122),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1147),
.A2(n_754),
.B1(n_499),
.B2(n_561),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1205),
.Y(n_1365)
);

BUFx2_ASAP7_75t_SL g1366 ( 
.A(n_1211),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1201),
.A2(n_1232),
.B(n_1185),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1234),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1253),
.A2(n_1364),
.B(n_1320),
.C(n_1345),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_L g1370 ( 
.A1(n_1255),
.A2(n_1256),
.B(n_1259),
.C(n_1250),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1323),
.B(n_1241),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1249),
.B(n_1236),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1323),
.B(n_1236),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1344),
.A2(n_1358),
.B(n_1300),
.Y(n_1375)
);

O2A1O1Ixp5_ASAP7_75t_L g1376 ( 
.A1(n_1268),
.A2(n_1283),
.B(n_1242),
.C(n_1297),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1343),
.A2(n_1274),
.B1(n_1356),
.B2(n_1357),
.Y(n_1377)
);

AND2x4_ASAP7_75t_SL g1378 ( 
.A(n_1311),
.B(n_1349),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1332),
.B(n_1362),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1308),
.B(n_1261),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1278),
.A2(n_1352),
.B1(n_1251),
.B2(n_1257),
.Y(n_1381)
);

OA22x2_ASAP7_75t_L g1382 ( 
.A1(n_1301),
.A2(n_1247),
.B1(n_1355),
.B2(n_1270),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1240),
.B(n_1247),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1269),
.A2(n_1275),
.B(n_1289),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1355),
.B(n_1270),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1308),
.B(n_1261),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1361),
.A2(n_1258),
.B(n_1335),
.C(n_1254),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1312),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1319),
.B(n_1261),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1305),
.A2(n_1329),
.B1(n_1272),
.B2(n_1318),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1351),
.B(n_1299),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1286),
.A2(n_1295),
.B(n_1290),
.C(n_1351),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1273),
.B(n_1296),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1351),
.B(n_1243),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1361),
.A2(n_1280),
.B(n_1267),
.C(n_1277),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1305),
.A2(n_1312),
.B1(n_1317),
.B2(n_1319),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1347),
.B(n_1294),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1305),
.A2(n_1317),
.B1(n_1316),
.B2(n_1366),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1244),
.B(n_1327),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1366),
.A2(n_1353),
.B1(n_1354),
.B2(n_1289),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1331),
.B(n_1339),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1248),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1346),
.B(n_1365),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1310),
.B(n_1263),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1304),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1295),
.B(n_1306),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1306),
.B(n_1354),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1280),
.A2(n_1275),
.B(n_1338),
.C(n_1265),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_SL g1410 ( 
.A1(n_1260),
.A2(n_1328),
.B(n_1330),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1269),
.A2(n_1334),
.B(n_1353),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1298),
.B(n_1269),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1260),
.A2(n_1368),
.B(n_1359),
.C(n_1350),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1309),
.B(n_1313),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1298),
.B(n_1269),
.Y(n_1415)
);

AOI211xp5_ASAP7_75t_L g1416 ( 
.A1(n_1271),
.A2(n_1363),
.B(n_1334),
.C(n_1314),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1291),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1260),
.A2(n_1368),
.B(n_1359),
.C(n_1350),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1302),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1337),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1276),
.B(n_1368),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1284),
.A2(n_1281),
.B(n_1246),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1276),
.B(n_1328),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1315),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1330),
.B(n_1282),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1287),
.A2(n_1363),
.B1(n_1282),
.B2(n_1235),
.Y(n_1426)
);

OAI211xp5_ASAP7_75t_L g1427 ( 
.A1(n_1282),
.A2(n_1293),
.B(n_1292),
.C(n_1235),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1237),
.B(n_1324),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1287),
.A2(n_1235),
.B1(n_1252),
.B2(n_1303),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1252),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1284),
.A2(n_1281),
.B(n_1246),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1235),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1237),
.B(n_1324),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1307),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1336),
.A2(n_1293),
.B1(n_1292),
.B2(n_1266),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1237),
.B(n_1324),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1307),
.B(n_1285),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1307),
.B(n_1288),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1266),
.B(n_1293),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1266),
.B(n_1292),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1336),
.A2(n_1288),
.B(n_1262),
.C(n_1239),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1288),
.B(n_1336),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1262),
.B(n_1239),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1321),
.A2(n_1333),
.B(n_1360),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1238),
.B(n_1321),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1322),
.A2(n_1341),
.B(n_1325),
.C(n_1326),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1333),
.A2(n_1341),
.B(n_1348),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1367),
.A2(n_1343),
.B1(n_1147),
.B2(n_1241),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1367),
.A2(n_1343),
.B1(n_1147),
.B2(n_1241),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1245),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1343),
.A2(n_1147),
.B1(n_1241),
.B2(n_1162),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1259),
.A2(n_1284),
.B(n_1114),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1247),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1453),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1373),
.B(n_1383),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1417),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1425),
.B(n_1421),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1379),
.B(n_1402),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1407),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1423),
.B(n_1433),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1409),
.B(n_1441),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1407),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1428),
.B(n_1436),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1444),
.A2(n_1447),
.B(n_1441),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1437),
.B(n_1452),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1452),
.B(n_1370),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_1395),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1450),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1424),
.B(n_1371),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1451),
.A2(n_1377),
.B1(n_1448),
.B2(n_1449),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1395),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1375),
.B(n_1390),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1409),
.B(n_1384),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1439),
.A2(n_1376),
.B(n_1427),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1438),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1369),
.A2(n_1416),
.B1(n_1385),
.B2(n_1389),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1442),
.B(n_1440),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1427),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1422),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1422),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1435),
.B(n_1445),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1369),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1413),
.B(n_1418),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1434),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1382),
.Y(n_1486)
);

NOR2x1_ASAP7_75t_L g1487 ( 
.A(n_1426),
.B(n_1387),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1431),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1382),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1412),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1431),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1374),
.B(n_1405),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1446),
.A2(n_1392),
.B(n_1410),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1393),
.B(n_1397),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1420),
.Y(n_1495)
);

INVxp67_ASAP7_75t_R g1496 ( 
.A(n_1396),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1476),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1476),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1458),
.B(n_1387),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1468),
.A2(n_1376),
.B(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1458),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1460),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1466),
.B(n_1394),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1458),
.B(n_1399),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1466),
.B(n_1372),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1454),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1470),
.B(n_1381),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1454),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1466),
.B(n_1380),
.Y(n_1509)
);

NOR2x1_ASAP7_75t_SL g1510 ( 
.A(n_1474),
.B(n_1398),
.Y(n_1510)
);

CKINVDCx14_ASAP7_75t_R g1511 ( 
.A(n_1495),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1386),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1480),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1478),
.B(n_1410),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1414),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1471),
.A2(n_1429),
.B1(n_1388),
.B2(n_1391),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1480),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1461),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1470),
.B(n_1401),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1488),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1457),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1467),
.B(n_1484),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1465),
.B(n_1415),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1471),
.A2(n_1400),
.B1(n_1419),
.B2(n_1408),
.Y(n_1525)
);

OAI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1500),
.A2(n_1473),
.B1(n_1487),
.B2(n_1477),
.C(n_1456),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1500),
.A2(n_1487),
.B(n_1468),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1497),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1501),
.Y(n_1530)
);

AOI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1499),
.A2(n_1489),
.B1(n_1486),
.B2(n_1479),
.C(n_1477),
.Y(n_1531)
);

OAI211xp5_ASAP7_75t_L g1532 ( 
.A1(n_1499),
.A2(n_1489),
.B(n_1479),
.C(n_1456),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1513),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1507),
.B(n_1430),
.Y(n_1534)
);

OA222x2_ASAP7_75t_L g1535 ( 
.A1(n_1507),
.A2(n_1474),
.B1(n_1483),
.B2(n_1462),
.C1(n_1472),
.C2(n_1482),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_R g1536 ( 
.A(n_1511),
.B(n_1432),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1523),
.B(n_1485),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1463),
.Y(n_1538)
);

NAND2x1_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_R g1541 ( 
.A(n_1511),
.B(n_1490),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1506),
.Y(n_1542)
);

NOR2x1_ASAP7_75t_SL g1543 ( 
.A(n_1502),
.B(n_1474),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1506),
.Y(n_1544)
);

AOI221x1_ASAP7_75t_L g1545 ( 
.A1(n_1522),
.A2(n_1411),
.B1(n_1472),
.B2(n_1408),
.C(n_1469),
.Y(n_1545)
);

OAI33xp33_ASAP7_75t_L g1546 ( 
.A1(n_1522),
.A2(n_1455),
.A3(n_1459),
.B1(n_1464),
.B2(n_1482),
.B3(n_1461),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1516),
.A2(n_1485),
.B1(n_1496),
.B2(n_1474),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1492),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

AOI222xp33_ASAP7_75t_L g1551 ( 
.A1(n_1516),
.A2(n_1485),
.B1(n_1484),
.B2(n_1467),
.C1(n_1455),
.C2(n_1378),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1492),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1525),
.A2(n_1496),
.B1(n_1483),
.B2(n_1474),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1501),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1523),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1508),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1517),
.A2(n_1465),
.B(n_1481),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1504),
.B(n_1492),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1510),
.A2(n_1474),
.B(n_1483),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1515),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1498),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1504),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1505),
.B(n_1494),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1508),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1515),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1557),
.A2(n_1528),
.B(n_1559),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1555),
.B(n_1519),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1540),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1555),
.B(n_1530),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1533),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1554),
.B(n_1505),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1557),
.A2(n_1465),
.B(n_1488),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1542),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1561),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1562),
.B(n_1505),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1514),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1544),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1556),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1556),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1549),
.B(n_1552),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1527),
.B(n_1498),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1545),
.A2(n_1491),
.B(n_1517),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1545),
.A2(n_1491),
.B(n_1517),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1529),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1531),
.A2(n_1491),
.B(n_1521),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1564),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1526),
.B(n_1525),
.C(n_1467),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_SL g1592 ( 
.A(n_1534),
.B(n_1524),
.C(n_1484),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1564),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1553),
.A2(n_1483),
.B(n_1459),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1550),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1597)
);

INVx4_ASAP7_75t_SL g1598 ( 
.A(n_1529),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1532),
.B(n_1483),
.C(n_1475),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1599),
.B(n_1539),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1599),
.A2(n_1518),
.B(n_1521),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1598),
.B(n_1535),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1598),
.B(n_1535),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1567),
.Y(n_1606)
);

INVx3_ASAP7_75t_SL g1607 ( 
.A(n_1598),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1567),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1598),
.B(n_1543),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1611)
);

AOI211xp5_ASAP7_75t_L g1612 ( 
.A1(n_1591),
.A2(n_1548),
.B(n_1553),
.C(n_1546),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1570),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1614)
);

OAI211xp5_ASAP7_75t_L g1615 ( 
.A1(n_1591),
.A2(n_1551),
.B(n_1536),
.C(n_1539),
.Y(n_1615)
);

NAND4xp25_ASAP7_75t_L g1616 ( 
.A(n_1592),
.B(n_1482),
.C(n_1403),
.D(n_1404),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1570),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1578),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1575),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1580),
.B(n_1543),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1594),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1537),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1547),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1566),
.B(n_1510),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1589),
.B(n_1550),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1589),
.A2(n_1483),
.B(n_1493),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1566),
.B(n_1510),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1566),
.B(n_1560),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1568),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1589),
.B(n_1514),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1584),
.B(n_1563),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1589),
.B(n_1538),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1586),
.B(n_1538),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1576),
.B(n_1515),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1568),
.B(n_1572),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1576),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1607),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1588),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1622),
.A2(n_1483),
.B1(n_1496),
.B2(n_1573),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1603),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1606),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1616),
.A2(n_1586),
.B1(n_1587),
.B2(n_1462),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.Y(n_1647)
);

NOR2x1p5_ASAP7_75t_SL g1648 ( 
.A(n_1628),
.B(n_1572),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1616),
.A2(n_1587),
.B1(n_1462),
.B2(n_1571),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1612),
.B(n_1541),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1609),
.Y(n_1652)
);

OR4x1_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1588),
.C(n_1581),
.D(n_1582),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1579),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1613),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1608),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1608),
.B(n_1577),
.Y(n_1657)
);

AOI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1615),
.A2(n_1587),
.B(n_1571),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1509),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1607),
.B(n_1509),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1615),
.B(n_1596),
.C(n_1572),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1603),
.A2(n_1585),
.B(n_1569),
.C(n_1573),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1611),
.B(n_1634),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1619),
.B(n_1512),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1607),
.Y(n_1665)
);

AOI322xp5_ASAP7_75t_L g1666 ( 
.A1(n_1622),
.A2(n_1509),
.A3(n_1503),
.B1(n_1512),
.B2(n_1498),
.C1(n_1582),
.C2(n_1593),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1624),
.B(n_1585),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1617),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1629),
.A2(n_1569),
.B(n_1462),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1610),
.B(n_1577),
.Y(n_1672)
);

NAND4xp25_ASAP7_75t_L g1673 ( 
.A(n_1603),
.B(n_1581),
.C(n_1590),
.D(n_1583),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1624),
.B(n_1623),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1512),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1601),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1642),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1674),
.B(n_1644),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1651),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1665),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1670),
.B(n_1611),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1614),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1656),
.B(n_1623),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1661),
.A2(n_1604),
.B1(n_1600),
.B2(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1652),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1658),
.A2(n_1604),
.B1(n_1600),
.B2(n_1601),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1663),
.B(n_1638),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1667),
.B(n_1604),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1659),
.B(n_1610),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1657),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1646),
.B(n_1605),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1657),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1657),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1655),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1677),
.A2(n_1646),
.B(n_1650),
.C(n_1662),
.Y(n_1701)
);

AOI22x1_ASAP7_75t_L g1702 ( 
.A1(n_1699),
.A2(n_1605),
.B1(n_1618),
.B2(n_1668),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1699),
.A2(n_1647),
.B(n_1626),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1680),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1680),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1681),
.A2(n_1648),
.B(n_1671),
.C(n_1662),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1693),
.B(n_1660),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1682),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1686),
.A2(n_1650),
.B1(n_1600),
.B2(n_1643),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1696),
.A2(n_1600),
.B(n_1601),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1682),
.Y(n_1712)
);

OAI32xp33_ASAP7_75t_L g1713 ( 
.A1(n_1684),
.A2(n_1618),
.A3(n_1605),
.B1(n_1653),
.B2(n_1633),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1696),
.A2(n_1600),
.B(n_1666),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1684),
.A2(n_1688),
.B1(n_1685),
.B2(n_1683),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

OAI32xp33_ASAP7_75t_L g1717 ( 
.A1(n_1691),
.A2(n_1676),
.A3(n_1697),
.B1(n_1695),
.B2(n_1618),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1675),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1678),
.A2(n_1600),
.B(n_1601),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1704),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1705),
.B(n_1679),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1707),
.B(n_1679),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1708),
.B(n_1679),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1702),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1709),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1715),
.B(n_1687),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1712),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1718),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1716),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1727),
.A2(n_1701),
.B1(n_1713),
.B2(n_1717),
.C(n_1715),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1725),
.A2(n_1714),
.B(n_1706),
.C(n_1711),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1725),
.A2(n_1706),
.B1(n_1719),
.B2(n_1710),
.C(n_1689),
.Y(n_1733)
);

OAI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1729),
.A2(n_1600),
.B1(n_1692),
.B2(n_1690),
.C(n_1700),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_SL g1735 ( 
.A(n_1724),
.B(n_1694),
.C(n_1692),
.D(n_1700),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1721),
.A2(n_1694),
.B1(n_1601),
.B2(n_1690),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1723),
.A2(n_1676),
.B1(n_1601),
.B2(n_1618),
.C(n_1605),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1722),
.B(n_1724),
.Y(n_1738)
);

AOI31xp33_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_1676),
.A3(n_1669),
.B(n_1664),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1721),
.A2(n_1720),
.B(n_1728),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1740),
.Y(n_1741)
);

OAI31xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1731),
.A2(n_1730),
.A3(n_1726),
.B(n_1630),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1738),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1735),
.B(n_1739),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1732),
.Y(n_1745)
);

AOI21xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1734),
.A2(n_1703),
.B(n_1647),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1742),
.B(n_1733),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1743),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1741),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1744),
.B(n_1737),
.C(n_1736),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1745),
.B(n_1621),
.Y(n_1751)
);

OAI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1746),
.A2(n_1672),
.B(n_1618),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1743),
.Y(n_1753)
);

XNOR2xp5_ASAP7_75t_L g1754 ( 
.A(n_1751),
.B(n_1703),
.Y(n_1754)
);

OAI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1747),
.A2(n_1703),
.B(n_1630),
.C(n_1627),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_R g1756 ( 
.A(n_1750),
.B(n_1672),
.Y(n_1756)
);

OA22x2_ASAP7_75t_L g1757 ( 
.A1(n_1752),
.A2(n_1672),
.B1(n_1625),
.B2(n_1630),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1749),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1753),
.C(n_1748),
.Y(n_1759)
);

AND3x2_ASAP7_75t_L g1760 ( 
.A(n_1756),
.B(n_1750),
.C(n_1625),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1754),
.B(n_1624),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1761),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1759),
.B1(n_1755),
.B2(n_1757),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1760),
.B1(n_1625),
.B2(n_1627),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1763),
.B(n_1675),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1632),
.B1(n_1635),
.B2(n_1602),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1765),
.A2(n_1632),
.B1(n_1635),
.B2(n_1602),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1767),
.A2(n_1635),
.B1(n_1632),
.B2(n_1602),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_L g1769 ( 
.A(n_1766),
.B(n_1627),
.C(n_1631),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1769),
.B(n_1631),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1626),
.B(n_1639),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1626),
.B1(n_1631),
.B2(n_1637),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1636),
.B1(n_1626),
.B2(n_1633),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1640),
.B(n_1617),
.C(n_1620),
.Y(n_1775)
);


endmodule