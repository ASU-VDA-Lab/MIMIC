module fake_jpeg_8147_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_26),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_16),
.C(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_35),
.C(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_58),
.B1(n_41),
.B2(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_43),
.B1(n_18),
.B2(n_20),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_66),
.B(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_33),
.B(n_21),
.C(n_28),
.Y(n_66)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_74),
.B1(n_56),
.B2(n_63),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_76),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_41),
.B1(n_43),
.B2(n_28),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_27),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_27),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_23),
.C(n_26),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_37),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_0),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_62),
.B1(n_20),
.B2(n_29),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_103),
.B1(n_110),
.B2(n_67),
.Y(n_120)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_51),
.B1(n_62),
.B2(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_17),
.B(n_25),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_114),
.C(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_17),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_90),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_67),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_25),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_119),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_123),
.B1(n_98),
.B2(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_87),
.B1(n_68),
.B2(n_70),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_68),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_98),
.B(n_113),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_149),
.B(n_152),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_84),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_146),
.B(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_154),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_153),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_84),
.B(n_109),
.Y(n_146)
);

AO21x1_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_117),
.B(n_118),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_94),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_156),
.C(n_160),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_70),
.B(n_77),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_128),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_101),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_2),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_146),
.B1(n_142),
.B2(n_152),
.Y(n_192)
);

NOR4xp25_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_132),
.C(n_126),
.D(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_179),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_126),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_172),
.C(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_160),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_129),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_119),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_181),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_124),
.B1(n_135),
.B2(n_78),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_182),
.A2(n_159),
.B1(n_174),
.B2(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_195),
.C(n_197),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_166),
.B(n_183),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_146),
.B1(n_141),
.B2(n_157),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_183),
.B1(n_178),
.B2(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_156),
.C(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_157),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_162),
.C(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_106),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_106),
.C(n_97),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.C(n_25),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_95),
.C(n_82),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_203),
.B(n_204),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_170),
.B1(n_163),
.B2(n_181),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_215),
.B(n_69),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_163),
.B1(n_171),
.B2(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_78),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_176),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_210),
.C(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_77),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_95),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_78),
.B(n_69),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_200),
.C(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_218),
.C(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_201),
.C(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_31),
.Y(n_232)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_211),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_15),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_15),
.C(n_14),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_13),
.C(n_69),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_226),
.Y(n_231)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_214),
.A3(n_202),
.B1(n_210),
.B2(n_215),
.C1(n_31),
.C2(n_8),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_2),
.Y(n_238)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_241),
.B1(n_233),
.B2(n_229),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_231),
.B1(n_230),
.B2(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.C(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_4),
.C(n_5),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_4),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_245),
.A3(n_246),
.B1(n_240),
.B2(n_238),
.C1(n_8),
.C2(n_9),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_5),
.B(n_6),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_6),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_245),
.B(n_7),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_251),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_9),
.Y(n_254)
);


endmodule