module fake_jpeg_25346_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_35),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_17),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_37),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_24),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_58),
.B(n_40),
.C(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_62),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_32),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_91),
.B1(n_37),
.B2(n_40),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_22),
.A3(n_45),
.B1(n_20),
.B2(n_44),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_81),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_35),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_36),
.A3(n_19),
.B1(n_33),
.B2(n_41),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_80),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_41),
.B(n_29),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_95),
.B1(n_46),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_21),
.B1(n_16),
.B2(n_36),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_36),
.B1(n_46),
.B2(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_44),
.A3(n_42),
.B1(n_39),
.B2(n_27),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_33),
.B1(n_29),
.B2(n_46),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_102),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_44),
.C(n_51),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_44),
.C(n_40),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_59),
.B1(n_39),
.B2(n_63),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_122),
.B1(n_84),
.B2(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_118),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_59),
.B1(n_15),
.B2(n_11),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_92),
.B1(n_74),
.B2(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_35),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_38),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_136),
.B1(n_149),
.B2(n_126),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_134),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_155),
.B1(n_100),
.B2(n_114),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_117),
.B(n_114),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_124),
.B1(n_119),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_141),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_75),
.B1(n_72),
.B2(n_76),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_142),
.B1(n_153),
.B2(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_75),
.B1(n_82),
.B2(n_42),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_142),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_44),
.B1(n_80),
.B2(n_42),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_121),
.B(n_37),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_44),
.C(n_40),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_125),
.C(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_189),
.C(n_34),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_169),
.B1(n_151),
.B2(n_144),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_125),
.B1(n_126),
.B2(n_99),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_191),
.B1(n_167),
.B2(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_104),
.B1(n_116),
.B2(n_117),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_147),
.B(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_175),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_187),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_176),
.B(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_181),
.B1(n_148),
.B2(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_188),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_17),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_23),
.B(n_17),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_38),
.A3(n_27),
.B1(n_23),
.B2(n_32),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_38),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_101),
.C(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_101),
.B1(n_26),
.B2(n_25),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_204),
.B1(n_206),
.B2(n_216),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_141),
.B(n_138),
.C(n_32),
.D(n_23),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_185),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_160),
.CI(n_163),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_222),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_152),
.B1(n_26),
.B2(n_34),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_32),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_209),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_34),
.B1(n_38),
.B2(n_23),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_212),
.C(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_14),
.C(n_13),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_14),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_169),
.B1(n_166),
.B2(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_160),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_185),
.B1(n_186),
.B2(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_0),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_12),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_213),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_168),
.B(n_183),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_226),
.B(n_238),
.Y(n_250)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_225),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_176),
.B(n_188),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_228),
.A2(n_216),
.B1(n_214),
.B2(n_210),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_12),
.C(n_11),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_236),
.C(n_212),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_234),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_11),
.C(n_10),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_0),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_9),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_9),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_0),
.B(n_1),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_206),
.B(n_202),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_8),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_195),
.C(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_246),
.B1(n_238),
.B2(n_231),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_1),
.Y(n_285)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_208),
.C(n_221),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_198),
.CI(n_214),
.CON(n_264),
.SN(n_264)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_266),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_204),
.C(n_10),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_8),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_278),
.B1(n_250),
.B2(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_2),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_226),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_281),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_246),
.B1(n_238),
.B2(n_229),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_230),
.B(n_243),
.C(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_227),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_233),
.C(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_263),
.C(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_241),
.B1(n_225),
.B2(n_240),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_2),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_252),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_250),
.B(n_264),
.C(n_269),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_285),
.B(n_282),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_297),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_298),
.Y(n_311)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_256),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_275),
.B(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_310),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

INVx11_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_281),
.C(n_276),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_286),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_4),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_290),
.B(n_289),
.Y(n_315)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_294),
.C(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_310),
.C(n_305),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_5),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_7),
.B(n_5),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_5),
.B(n_6),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_304),
.Y(n_328)
);

NOR2x1_ASAP7_75t_R g325 ( 
.A(n_316),
.B(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_309),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_329),
.C(n_331),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_326),
.C(n_323),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_323),
.B1(n_312),
.B2(n_304),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_320),
.C(n_303),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule