module fake_jpeg_8064_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_22),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_16),
.C(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_17),
.C(n_19),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_21),
.B1(n_32),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_67),
.B1(n_19),
.B2(n_20),
.Y(n_110)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_64),
.B1(n_68),
.B2(n_72),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_17),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_32),
.B1(n_21),
.B2(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_31),
.B1(n_16),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_30),
.B1(n_25),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_30),
.B1(n_25),
.B2(n_26),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_29),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_29),
.CI(n_38),
.CON(n_104),
.SN(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_77),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_71),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_41),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_106),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_102),
.B(n_104),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_33),
.B(n_22),
.C(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_109),
.B1(n_27),
.B2(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_48),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_20),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_47),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_37),
.B1(n_17),
.B2(n_19),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_23),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_0),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_27),
.B(n_23),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_29),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

OAI22x1_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_38),
.B1(n_36),
.B2(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_118),
.A2(n_119),
.B1(n_135),
.B2(n_136),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_145),
.B1(n_107),
.B2(n_90),
.Y(n_171)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_82),
.A2(n_65),
.B1(n_59),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_75),
.B1(n_58),
.B2(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_24),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_143),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_91),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_38),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_58),
.B1(n_56),
.B2(n_51),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_97),
.B1(n_104),
.B2(n_106),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_171),
.B1(n_119),
.B2(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_152),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_86),
.B1(n_102),
.B2(n_92),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_133),
.B1(n_138),
.B2(n_90),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_98),
.B(n_104),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_165),
.B(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_106),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_161),
.B(n_124),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_97),
.B(n_103),
.C(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_177),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_166),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_170),
.C(n_124),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_113),
.B(n_97),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_113),
.B(n_83),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_112),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_36),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_117),
.B(n_84),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_80),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_94),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_R g180 ( 
.A(n_129),
.B(n_38),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_144),
.B(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_165),
.B1(n_161),
.B2(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_156),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_195),
.B1(n_202),
.B2(n_197),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_189),
.B1(n_211),
.B2(n_151),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_201),
.B(n_205),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_134),
.B1(n_124),
.B2(n_143),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_194),
.C(n_208),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_147),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_146),
.B1(n_133),
.B2(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

FAx1_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_24),
.CI(n_16),
.CON(n_201),
.SN(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_101),
.B1(n_99),
.B2(n_127),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_212),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_127),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_24),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_156),
.B(n_144),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_101),
.B1(n_99),
.B2(n_86),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_11),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_51),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_161),
.B1(n_167),
.B2(n_160),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_220),
.B(n_200),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_214),
.A2(n_160),
.B1(n_169),
.B2(n_156),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_222),
.B(n_226),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_14),
.C(n_13),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_227),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_235),
.B1(n_188),
.B2(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_0),
.B(n_1),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_158),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_240),
.C(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_238),
.B1(n_200),
.B2(n_182),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_184),
.A2(n_151),
.B1(n_132),
.B2(n_111),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_189),
.B1(n_183),
.B2(n_204),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_237),
.B1(n_199),
.B2(n_207),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_1),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_183),
.B1(n_201),
.B2(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_248),
.B1(n_249),
.B2(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_233),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_250),
.C(n_259),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_235),
.B1(n_239),
.B2(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_254),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_182),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_263),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_201),
.B1(n_188),
.B2(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_216),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_194),
.C(n_208),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_232),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_226),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_205),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_215),
.A2(n_205),
.B1(n_203),
.B2(n_4),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_234),
.B1(n_244),
.B2(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_274),
.B1(n_278),
.B2(n_281),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_257),
.B1(n_243),
.B2(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_221),
.C(n_218),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_276),
.C(n_264),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_218),
.C(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_227),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_220),
.B1(n_219),
.B2(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_240),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_2),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_2),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

AO21x2_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_246),
.B(n_242),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_287),
.B(n_269),
.Y(n_301)
);

FAx1_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_242),
.CI(n_263),
.CON(n_287),
.SN(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_247),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_293),
.C(n_273),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_250),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_7),
.B(n_8),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_297),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_253),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_271),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

BUFx12_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_265),
.A2(n_262),
.B1(n_4),
.B2(n_6),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_281),
.B1(n_279),
.B2(n_271),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_275),
.B(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_304),
.B1(n_284),
.B2(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_285),
.B1(n_286),
.B2(n_299),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_273),
.C(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_267),
.C(n_269),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_3),
.C(n_6),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_7),
.C(n_8),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_311),
.C(n_9),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_7),
.C(n_8),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_292),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_295),
.B1(n_290),
.B2(n_284),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_320),
.C(n_319),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_305),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_324),
.C(n_325),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_313),
.C(n_310),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_297),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_9),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_320),
.B1(n_10),
.B2(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_330),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_323),
.B(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_321),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_9),
.Y(n_337)
);


endmodule