module fake_jpeg_27165_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_16),
.C(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_15),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_66),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_22),
.B1(n_23),
.B2(n_14),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_17),
.B1(n_43),
.B2(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_45),
.B1(n_52),
.B2(n_13),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_33),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_17),
.B1(n_36),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_51),
.B1(n_49),
.B2(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_33),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_76),
.Y(n_79)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_25),
.C(n_14),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_91),
.B1(n_76),
.B2(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_51),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_0),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_70),
.B(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_61),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_104),
.Y(n_107)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_74),
.C(n_60),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_65),
.A3(n_90),
.B1(n_81),
.B2(n_9),
.C1(n_8),
.C2(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_90),
.C(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_85),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_108),
.B(n_86),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_104),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_119),
.C(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_90),
.C(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_98),
.B1(n_57),
.B2(n_60),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_114),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_126),
.C(n_118),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_83),
.B(n_67),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_93),
.B(n_71),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_116),
.C(n_117),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_71),
.C(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_2),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_130),
.A3(n_75),
.B1(n_121),
.B2(n_72),
.C1(n_78),
.C2(n_57),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_77),
.C(n_78),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_2),
.Y(n_137)
);


endmodule