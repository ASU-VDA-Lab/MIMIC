module fake_aes_8089_n_1012 (n_120, n_136, n_155, n_107, n_103, n_157, n_52, n_162, n_114, n_156, n_154, n_50, n_7, n_3, n_34, n_142, n_25, n_9, n_163, n_96, n_72, n_77, n_90, n_169, n_178, n_180, n_99, n_43, n_73, n_62, n_167, n_97, n_133, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_153, n_187, n_66, n_88, n_46, n_121, n_174, n_188, n_108, n_161, n_37, n_122, n_165, n_18, n_65, n_87, n_5, n_81, n_85, n_112, n_102, n_172, n_47, n_109, n_1, n_16, n_78, n_95, n_40, n_68, n_105, n_36, n_11, n_115, n_179, n_15, n_168, n_139, n_152, n_151, n_71, n_117, n_176, n_70, n_94, n_2, n_17, n_58, n_113, n_20, n_84, n_130, n_12, n_56, n_80, n_67, n_116, n_22, n_118, n_19, n_26, n_39, n_101, n_98, n_150, n_38, n_104, n_100, n_159, n_24, n_141, n_35, n_91, n_146, n_160, n_32, n_148, n_149, n_93, n_143, n_134, n_48, n_63, n_54, n_125, n_41, n_147, n_55, n_145, n_185, n_29, n_166, n_173, n_181, n_123, n_171, n_60, n_135, n_138, n_140, n_111, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_183, n_64, n_132, n_69, n_175, n_127, n_128, n_170, n_83, n_158, n_23, n_0, n_126, n_110, n_184, n_182, n_119, n_57, n_51, n_144, n_106, n_186, n_45, n_42, n_21, n_137, n_131, n_86, n_27, n_124, n_89, n_177, n_28, n_79, n_129, n_164, n_49, n_14, n_31, n_1012, n_981);
input n_120;
input n_136;
input n_155;
input n_107;
input n_103;
input n_157;
input n_52;
input n_162;
input n_114;
input n_156;
input n_154;
input n_50;
input n_7;
input n_3;
input n_34;
input n_142;
input n_25;
input n_9;
input n_163;
input n_96;
input n_72;
input n_77;
input n_90;
input n_169;
input n_178;
input n_180;
input n_99;
input n_43;
input n_73;
input n_62;
input n_167;
input n_97;
input n_133;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_153;
input n_187;
input n_66;
input n_88;
input n_46;
input n_121;
input n_174;
input n_188;
input n_108;
input n_161;
input n_37;
input n_122;
input n_165;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_112;
input n_102;
input n_172;
input n_47;
input n_109;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_105;
input n_36;
input n_11;
input n_115;
input n_179;
input n_15;
input n_168;
input n_139;
input n_152;
input n_151;
input n_71;
input n_117;
input n_176;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_113;
input n_20;
input n_84;
input n_130;
input n_12;
input n_56;
input n_80;
input n_67;
input n_116;
input n_22;
input n_118;
input n_19;
input n_26;
input n_39;
input n_101;
input n_98;
input n_150;
input n_38;
input n_104;
input n_100;
input n_159;
input n_24;
input n_141;
input n_35;
input n_91;
input n_146;
input n_160;
input n_32;
input n_148;
input n_149;
input n_93;
input n_143;
input n_134;
input n_48;
input n_63;
input n_54;
input n_125;
input n_41;
input n_147;
input n_55;
input n_145;
input n_185;
input n_29;
input n_166;
input n_173;
input n_181;
input n_123;
input n_171;
input n_60;
input n_135;
input n_138;
input n_140;
input n_111;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_183;
input n_64;
input n_132;
input n_69;
input n_175;
input n_127;
input n_128;
input n_170;
input n_83;
input n_158;
input n_23;
input n_0;
input n_126;
input n_110;
input n_184;
input n_182;
input n_119;
input n_57;
input n_51;
input n_144;
input n_106;
input n_186;
input n_45;
input n_42;
input n_21;
input n_137;
input n_131;
input n_86;
input n_27;
input n_124;
input n_89;
input n_177;
input n_28;
input n_79;
input n_129;
input n_164;
input n_49;
input n_14;
input n_31;
output n_1012;
output n_981;
wire n_890;
wire n_107;
wire n_646;
wire n_759;
wire n_987;
wire n_658;
wire n_673;
wire n_156;
wire n_239;
wire n_154;
wire n_7;
wire n_309;
wire n_944;
wire n_356;
wire n_895;
wire n_327;
wire n_25;
wire n_994;
wire n_204;
wire n_592;
wire n_769;
wire n_929;
wire n_169;
wire n_384;
wire n_370;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_44;
wire n_394;
wire n_189;
wire n_681;
wire n_352;
wire n_226;
wire n_447;
wire n_66;
wire n_379;
wire n_903;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_952;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_949;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_942;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_753;
wire n_859;
wire n_436;
wire n_438;
wire n_900;
wire n_869;
wire n_931;
wire n_935;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_971;
wire n_482;
wire n_838;
wire n_967;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_963;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_961;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_553;
wire n_494;
wire n_555;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_981;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_990;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_993;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_977;
wire n_772;
wire n_50;
wire n_789;
wire n_816;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_999;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_991;
wire n_133;
wire n_324;
wire n_442;
wire n_982;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_998;
wire n_578;
wire n_928;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_801;
wire n_682;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_920;
wire n_912;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_905;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_934;
wire n_653;
wire n_351;
wire n_1;
wire n_979;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_989;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_984;
wire n_404;
wire n_289;
wire n_179;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_980;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_911;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_711;
wire n_491;
wire n_800;
wire n_973;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_906;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_879;
wire n_888;
wire n_576;
wire n_992;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_909;
wire n_493;
wire n_274;
wire n_910;
wire n_972;
wire n_235;
wire n_150;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_965;
wire n_100;
wire n_299;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_344;
wire n_232;
wire n_878;
wire n_783;
wire n_812;
wire n_147;
wire n_185;
wire n_367;
wire n_955;
wire n_795;
wire n_267;
wire n_1007;
wire n_687;
wire n_950;
wire n_171;
wire n_638;
wire n_873;
wire n_899;
wire n_450;
wire n_644;
wire n_140;
wire n_585;
wire n_111;
wire n_746;
wire n_212;
wire n_779;
wire n_978;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_728;
wire n_435;
wire n_704;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_970;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_986;
wire n_262;
wire n_921;
wire n_119;
wire n_667;
wire n_503;
wire n_969;
wire n_856;
wire n_927;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_904;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_325;
wire n_273;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_951;
wire n_163;
wire n_348;
wire n_96;
wire n_669;
wire n_685;
wire n_90;
wire n_77;
wire n_72;
wire n_594;
wire n_762;
wire n_214;
wire n_787;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_908;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_355;
wire n_153;
wire n_216;
wire n_609;
wire n_946;
wire n_121;
wire n_286;
wire n_408;
wire n_1003;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_65;
wire n_537;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_932;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_297;
wire n_276;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_854;
wire n_523;
wire n_815;
wire n_901;
wire n_528;
wire n_419;
wire n_985;
wire n_252;
wire n_922;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_966;
wire n_693;
wire n_1011;
wire n_785;
wire n_896;
wire n_739;
wire n_94;
wire n_997;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_741;
wire n_698;
wire n_257;
wire n_705;
wire n_828;
wire n_722;
wire n_988;
wire n_203;
wire n_26;
wire n_477;
wire n_996;
wire n_460;
wire n_318;
wire n_243;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_337;
wire n_146;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_872;
wire n_957;
wire n_93;
wire n_539;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_923;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_918;
wire n_1009;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_948;
wire n_732;
wire n_926;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_1001;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_1006;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_925;
wire n_205;
wire n_158;
wire n_915;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_975;
wire n_89;
wire n_480;
wire n_939;
wire n_940;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_260;
wire n_136;
wire n_891;
wire n_1004;
wire n_1002;
wire n_580;
wire n_976;
wire n_610;
wire n_938;
wire n_1008;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_964;
wire n_34;
wire n_142;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_943;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_956;
wire n_781;
wire n_954;
wire n_914;
wire n_945;
wire n_852;
wire n_376;
wire n_902;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_87;
wire n_466;
wire n_207;
wire n_197;
wire n_81;
wire n_541;
wire n_572;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_983;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_919;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_36;
wire n_416;
wire n_962;
wire n_916;
wire n_870;
wire n_889;
wire n_432;
wire n_913;
wire n_917;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_960;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_796;
wire n_804;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_907;
wire n_591;
wire n_391;
wire n_209;
wire n_241;
wire n_874;
wire n_84;
wire n_20;
wire n_782;
wire n_449;
wire n_832;
wire n_56;
wire n_12;
wire n_412;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_862;
wire n_930;
wire n_819;
wire n_39;
wire n_101;
wire n_953;
wire n_941;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_933;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_947;
wire n_840;
wire n_1010;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_968;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_138;
wire n_60;
wire n_936;
wire n_937;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_924;
wire n_745;
wire n_305;
wire n_495;
wire n_430;
wire n_505;
wire n_418;
wire n_313;
wire n_358;
wire n_333;
wire n_92;
wire n_627;
wire n_740;
wire n_706;
wire n_589;
wire n_750;
wire n_175;
wire n_897;
wire n_128;
wire n_306;
wire n_415;
wire n_31;
wire n_697;
wire n_958;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_974;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_1000;
wire n_1005;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_995;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_349;
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_101), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_184), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_9), .Y(n_191) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_71), .Y(n_192) );
NOR2xp67_ASAP7_75t_L g193 ( .A(n_163), .B(n_16), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_6), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_22), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_161), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_24), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_36), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_50), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_79), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_46), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_120), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_160), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_129), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_186), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_148), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_169), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_126), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_110), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_111), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_17), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_47), .Y(n_217) );
NOR2xp67_ASAP7_75t_L g218 ( .A(n_49), .B(n_84), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_127), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_119), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_78), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_0), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_39), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_135), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_34), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_174), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_167), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_112), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_105), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_85), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_17), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_142), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_18), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_20), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_93), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_90), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_183), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_37), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_54), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_13), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_29), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_104), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_70), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_32), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_14), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_89), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_10), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_155), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_178), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_86), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_176), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_9), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_115), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_171), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_96), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_138), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_50), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_37), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_166), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_168), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_151), .Y(n_266) );
XNOR2xp5_ASAP7_75t_L g267 ( .A(n_125), .B(n_47), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_177), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_175), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_131), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_68), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_25), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_83), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_29), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_39), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_121), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_36), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_23), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_173), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_109), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_130), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_10), .Y(n_282) );
XNOR2x1_ASAP7_75t_L g283 ( .A(n_80), .B(n_95), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_56), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_42), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_49), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_64), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_100), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_19), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_25), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_76), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_164), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_117), .Y(n_293) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_91), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_132), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_159), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_128), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_133), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_0), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_180), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_67), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_106), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_137), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_165), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_6), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_38), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_7), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_69), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_122), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_252), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_217), .Y(n_311) );
AOI22x1_ASAP7_75t_SL g312 ( .A1(n_195), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
OAI22xp5_ASAP7_75t_SL g314 ( .A1(n_195), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_217), .Y(n_316) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_190), .A2(n_75), .B(n_74), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_242), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
BUFx2_ASAP7_75t_SL g320 ( .A(n_283), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_238), .B(n_4), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_242), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_254), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_252), .Y(n_324) );
AOI22x1_ASAP7_75t_SL g325 ( .A1(n_246), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_290), .Y(n_326) );
AND2x6_ASAP7_75t_L g327 ( .A(n_239), .B(n_77), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_201), .B(n_5), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_194), .B(n_8), .Y(n_331) );
BUFx8_ASAP7_75t_L g332 ( .A(n_254), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_301), .B(n_8), .Y(n_333) );
CKINVDCx6p67_ASAP7_75t_R g334 ( .A(n_240), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_190), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_254), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_234), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_268), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_263), .B(n_11), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_197), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_202), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_239), .B(n_14), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_340), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_313), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_341), .B(n_229), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_337), .A2(n_299), .B1(n_284), .B2(n_246), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_336), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_315), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_341), .B(n_189), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_343), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_343), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_336), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_313), .Y(n_358) );
AND3x1_ASAP7_75t_L g359 ( .A(n_337), .B(n_205), .C(n_191), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_342), .B(n_245), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_342), .B(n_204), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_343), .B(n_204), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_343), .B(n_206), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_332), .B(n_206), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_334), .B(n_294), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_334), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_332), .B(n_207), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_324), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_319), .B(n_208), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_200), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_319), .B(n_212), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_324), .B(n_207), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_324), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_313), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_321), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_333), .Y(n_380) );
OAI21xp33_ASAP7_75t_SL g381 ( .A1(n_311), .A2(n_283), .B(n_222), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_339), .A2(n_305), .B1(n_284), .B2(n_198), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_335), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_335), .Y(n_385) );
AND3x4_ASAP7_75t_L g386 ( .A(n_320), .B(n_218), .C(n_193), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_316), .B(n_211), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_336), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_331), .A2(n_215), .B(n_214), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_384), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_378), .B(n_320), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_347), .A2(n_360), .B(n_361), .Y(n_393) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_365), .B(n_317), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_378), .B(n_316), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_373), .A2(n_196), .B1(n_220), .B2(n_210), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_384), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_352), .B(n_298), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_373), .B(n_298), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_381), .A2(n_196), .B1(n_220), .B2(n_210), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_375), .B(n_303), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_362), .A2(n_317), .B(n_209), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_317), .B(n_209), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_345), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_385), .Y(n_408) );
AO22x1_ASAP7_75t_L g409 ( .A1(n_366), .A2(n_327), .B1(n_192), .B2(n_325), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_354), .B(n_294), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_344), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_389), .A2(n_354), .B1(n_355), .B2(n_367), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_355), .B(n_318), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_355), .B(n_322), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_353), .B(n_322), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_383), .A2(n_314), .B1(n_328), .B2(n_329), .C(n_326), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_371), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_387), .B(n_328), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_380), .B(n_329), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_382), .B(n_199), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_381), .A2(n_233), .B1(n_253), .B2(n_221), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_345), .B(n_216), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_389), .A2(n_327), .B1(n_223), .B2(n_237), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_367), .B(n_213), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_350), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_350), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_389), .A2(n_327), .B1(n_226), .B2(n_243), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_369), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_369), .B(n_219), .Y(n_433) );
XOR2xp5_ASAP7_75t_L g434 ( .A(n_349), .B(n_312), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_356), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_369), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_369), .B(n_224), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_359), .A2(n_221), .B1(n_253), .B2(n_233), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_364), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_359), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_386), .A2(n_327), .B1(n_241), .B2(n_247), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_372), .Y(n_442) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_374), .B(n_317), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_368), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_386), .B(n_225), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_388), .B(n_230), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_386), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_388), .B(n_236), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_346), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_357), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_379), .B(n_244), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_379), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_377), .A2(n_251), .B(n_256), .C(n_249), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_346), .A2(n_282), .B(n_285), .C(n_278), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_346), .B(n_227), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_358), .B(n_228), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_358), .B(n_266), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_377), .B(n_279), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_377), .B(n_280), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_377), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_377), .A2(n_293), .B1(n_295), .B2(n_292), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_348), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_461), .Y(n_463) );
BUFx2_ASAP7_75t_SL g464 ( .A(n_411), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_395), .B(n_292), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_395), .B(n_261), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_391), .A2(n_295), .B1(n_293), .B2(n_271), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_396), .B(n_305), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_392), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_442), .B(n_312), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_399), .A2(n_272), .B1(n_275), .B2(n_274), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_438), .B(n_286), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_448), .B(n_287), .Y(n_473) );
AO21x1_ASAP7_75t_L g474 ( .A1(n_404), .A2(n_232), .B(n_231), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_454), .A2(n_307), .B(n_308), .C(n_306), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_406), .A2(n_250), .B(n_248), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_448), .B(n_267), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_436), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_413), .Y(n_479) );
BUFx8_ASAP7_75t_L g480 ( .A(n_440), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_441), .A2(n_258), .B1(n_260), .B2(n_259), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_400), .B(n_203), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_423), .A2(n_262), .B1(n_269), .B2(n_265), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_426), .B(n_281), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_398), .B(n_15), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_412), .A2(n_288), .B1(n_297), .B2(n_291), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_443), .A2(n_302), .B(n_300), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_426), .B(n_203), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_401), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_421), .A2(n_304), .B1(n_289), .B2(n_203), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_427), .A2(n_289), .B1(n_257), .B2(n_276), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_409), .B(n_289), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_443), .A2(n_257), .B(n_235), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_407), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_431), .A2(n_289), .B1(n_255), .B2(n_273), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_415), .A2(n_264), .B(n_273), .C(n_16), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_445), .B(n_309), .C(n_296), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_403), .A2(n_270), .B1(n_268), .B2(n_323), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_436), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_432), .A2(n_270), .B(n_268), .C(n_338), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_403), .B(n_327), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_439), .B(n_15), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_407), .B(n_313), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_439), .B(n_18), .Y(n_505) );
INVx4_ASAP7_75t_L g506 ( .A(n_416), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_434), .B(n_19), .Y(n_507) );
AO21x1_ASAP7_75t_L g508 ( .A1(n_455), .A2(n_338), .B(n_323), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_390), .A2(n_338), .B(n_323), .C(n_23), .Y(n_509) );
BUFx12f_ASAP7_75t_L g510 ( .A(n_451), .Y(n_510) );
AO32x2_ASAP7_75t_L g511 ( .A1(n_460), .A2(n_338), .A3(n_323), .B1(n_24), .B2(n_26), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_424), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_402), .B(n_21), .Y(n_513) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_462), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_397), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_515) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_417), .B(n_28), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_444), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_422), .B(n_30), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_405), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_410), .A2(n_82), .B(n_81), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_420), .B(n_31), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_408), .B(n_33), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_428), .B(n_34), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_433), .B(n_35), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_437), .B(n_35), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_414), .B(n_38), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_419), .B(n_40), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_425), .B(n_40), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_451), .B(n_41), .Y(n_529) );
INVx3_ASAP7_75t_SL g530 ( .A(n_449), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_446), .B(n_41), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_429), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_430), .Y(n_533) );
NOR2xp33_ASAP7_75t_SL g534 ( .A(n_453), .B(n_87), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_457), .B(n_43), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_435), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_458), .A2(n_124), .B(n_182), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_435), .B(n_43), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_456), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_459), .A2(n_123), .B(n_179), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_450), .A2(n_44), .B(n_45), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_452), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_411), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_441), .A2(n_48), .B1(n_51), .B2(n_52), .Y(n_544) );
CKINVDCx11_ASAP7_75t_R g545 ( .A(n_411), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_447), .A2(n_48), .B1(n_51), .B2(n_52), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_395), .B(n_53), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_407), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_391), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_395), .B(n_55), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_391), .B(n_56), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_393), .A2(n_57), .B(n_58), .C(n_59), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_411), .B(n_57), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_477), .B(n_58), .Y(n_554) );
BUFx2_ASAP7_75t_R g555 ( .A(n_464), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_543), .B(n_59), .Y(n_556) );
AO31x2_ASAP7_75t_L g557 ( .A1(n_474), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_557) );
OAI22x1_ASAP7_75t_L g558 ( .A1(n_468), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_543), .B(n_63), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_465), .B(n_63), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_476), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_488), .A2(n_134), .B(n_157), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_465), .B(n_66), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_479), .B(n_67), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_530), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_467), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_514), .A2(n_136), .B(n_154), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_72), .B(n_73), .C(n_88), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g572 ( .A(n_470), .B(n_72), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_545), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_527), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_547), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_523), .A2(n_73), .B(n_92), .C(n_94), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_525), .A2(n_97), .B(n_98), .C(n_99), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_480), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_469), .B(n_187), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_504), .A2(n_102), .B(n_103), .Y(n_581) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_496), .A2(n_107), .A3(n_108), .B(n_113), .Y(n_582) );
BUFx10_ASAP7_75t_L g583 ( .A(n_503), .Y(n_583) );
CKINVDCx9p33_ASAP7_75t_R g584 ( .A(n_505), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_518), .A2(n_114), .B(n_116), .C(n_118), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_550), .Y(n_586) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_492), .A2(n_139), .A3(n_140), .B(n_141), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_542), .A2(n_143), .B(n_144), .Y(n_588) );
INVx3_ASAP7_75t_SL g589 ( .A(n_507), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_553), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_519), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_484), .A2(n_145), .B1(n_146), .B2(n_147), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_472), .B(n_149), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_480), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_484), .B(n_150), .Y(n_596) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_466), .A2(n_551), .B(n_473), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_532), .A2(n_536), .B(n_533), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_487), .A2(n_535), .B(n_538), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_489), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_521), .A2(n_481), .B1(n_471), .B2(n_483), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_490), .B(n_485), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_529), .Y(n_603) );
AO31x2_ASAP7_75t_L g604 ( .A1(n_552), .A2(n_508), .A3(n_509), .B(n_491), .Y(n_604) );
INVx6_ASAP7_75t_SL g605 ( .A(n_493), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_528), .A2(n_531), .B(n_497), .C(n_475), .Y(n_606) );
AOI221x1_ASAP7_75t_L g607 ( .A1(n_541), .A2(n_544), .B1(n_491), .B2(n_520), .C(n_499), .Y(n_607) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_501), .A2(n_499), .A3(n_540), .B(n_537), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_534), .B(n_539), .C(n_524), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_486), .B(n_481), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_500), .A2(n_478), .B(n_482), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_516), .B(n_549), .Y(n_612) );
BUFx8_ASAP7_75t_L g613 ( .A(n_511), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_517), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_495), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_512), .B(n_544), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_548), .B(n_493), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_498), .B(n_548), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_546), .B(n_515), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_511), .B(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_543), .B(n_395), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_543), .B(n_396), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_463), .A2(n_490), .B1(n_514), .B2(n_465), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_484), .A2(n_381), .B(n_383), .C(n_487), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_463), .A2(n_490), .B1(n_514), .B2(n_465), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_526), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_543), .B(n_411), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_543), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_543), .B(n_506), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_477), .B(n_320), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_506), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_543), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_543), .B(n_396), .Y(n_640) );
AO31x2_ASAP7_75t_L g641 ( .A1(n_474), .A2(n_494), .A3(n_476), .B(n_496), .Y(n_641) );
NOR2xp33_ASAP7_75t_R g642 ( .A(n_545), .B(n_543), .Y(n_642) );
AO21x1_ASAP7_75t_L g643 ( .A1(n_494), .A2(n_496), .B(n_476), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_644) );
AOI21xp5_ASAP7_75t_SL g645 ( .A1(n_527), .A2(n_514), .B(n_506), .Y(n_645) );
OAI22x1_ASAP7_75t_L g646 ( .A1(n_468), .A2(n_423), .B1(n_400), .B2(n_434), .Y(n_646) );
AO32x2_ASAP7_75t_L g647 ( .A1(n_487), .A2(n_496), .A3(n_492), .B1(n_491), .B2(n_544), .Y(n_647) );
BUFx4f_ASAP7_75t_L g648 ( .A(n_510), .Y(n_648) );
CKINVDCx11_ASAP7_75t_R g649 ( .A(n_545), .Y(n_649) );
AOI21xp5_ASAP7_75t_SL g650 ( .A1(n_527), .A2(n_514), .B(n_506), .Y(n_650) );
NOR2xp33_ASAP7_75t_SL g651 ( .A(n_543), .B(n_461), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_502), .A2(n_476), .B(n_394), .Y(n_652) );
INVx5_ASAP7_75t_L g653 ( .A(n_510), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_484), .A2(n_381), .B(n_383), .C(n_487), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_506), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_484), .A2(n_381), .B1(n_349), .B2(n_383), .C(n_418), .Y(n_656) );
BUFx10_ASAP7_75t_L g657 ( .A(n_527), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_543), .B(n_465), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_545), .Y(n_659) );
AND2x6_ASAP7_75t_L g660 ( .A(n_527), .B(n_479), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_526), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_495), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_543), .B(n_366), .C(n_386), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_635), .B(n_623), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_567), .B(n_574), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_634), .B(n_653), .Y(n_666) );
INVx4_ASAP7_75t_L g667 ( .A(n_653), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_642), .B(n_580), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_634), .B(n_653), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_658), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_622), .A2(n_627), .B(n_625), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_629), .B(n_661), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_565), .Y(n_674) );
NOR2xp33_ASAP7_75t_R g675 ( .A(n_649), .B(n_573), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_631), .A2(n_636), .B(n_633), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_565), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_626), .A2(n_654), .B(n_597), .C(n_596), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_606), .A2(n_599), .B(n_560), .C(n_554), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_656), .A2(n_646), .B1(n_614), .B2(n_660), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_660), .B(n_580), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_648), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_640), .B(n_663), .Y(n_683) );
AO31x2_ASAP7_75t_L g684 ( .A1(n_643), .A2(n_644), .A3(n_652), .B(n_637), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_632), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_594), .A2(n_586), .B(n_576), .C(n_601), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_621), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_660), .B(n_612), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_660), .B(n_610), .Y(n_689) );
AO31x2_ASAP7_75t_L g690 ( .A1(n_616), .A2(n_628), .A3(n_624), .B(n_578), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_575), .B(n_603), .Y(n_691) );
CKINVDCx11_ASAP7_75t_R g692 ( .A(n_579), .Y(n_692) );
OAI221xp5_ASAP7_75t_SL g693 ( .A1(n_569), .A2(n_639), .B1(n_593), .B2(n_619), .C(n_556), .Y(n_693) );
BUFx2_ASAP7_75t_L g694 ( .A(n_561), .Y(n_694) );
AO21x2_ASAP7_75t_L g695 ( .A1(n_620), .A2(n_563), .B(n_609), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_568), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_566), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_564), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_555), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_602), .B(n_600), .Y(n_700) );
INVx8_ASAP7_75t_L g701 ( .A(n_659), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_595), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_651), .B(n_590), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_558), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_630), .B(n_657), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_657), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_562), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_641), .B(n_598), .Y(n_708) );
HB1xp67_ASAP7_75t_SL g709 ( .A(n_613), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_559), .B(n_589), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_605), .A2(n_617), .B1(n_592), .B2(n_647), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_572), .B(n_615), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_583), .B(n_638), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_584), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_641), .B(n_655), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_583), .A2(n_613), .B1(n_605), .B2(n_618), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_662), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_641), .B(n_611), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_604), .B(n_571), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_557), .B(n_604), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_557), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_557), .Y(n_722) );
AO31x2_ASAP7_75t_L g723 ( .A1(n_585), .A2(n_577), .A3(n_570), .B(n_588), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_581), .A2(n_608), .B(n_582), .Y(n_724) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_608), .A2(n_582), .B(n_587), .Y(n_725) );
AO31x2_ASAP7_75t_L g726 ( .A1(n_647), .A2(n_474), .A3(n_643), .B(n_607), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_591), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_635), .B(n_320), .Y(n_728) );
INVxp67_ASAP7_75t_L g729 ( .A(n_632), .Y(n_729) );
AOI21xp33_ASAP7_75t_SL g730 ( .A1(n_573), .A2(n_659), .B(n_396), .Y(n_730) );
OR2x6_ASAP7_75t_L g731 ( .A(n_645), .B(n_650), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_642), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_632), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_635), .B(n_320), .Y(n_734) );
BUFx2_ASAP7_75t_L g735 ( .A(n_642), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_632), .Y(n_736) );
BUFx8_ASAP7_75t_L g737 ( .A(n_561), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_591), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_567), .B(n_574), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g740 ( .A1(n_656), .A2(n_381), .B(n_654), .C(n_626), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_621), .B(n_543), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_649), .Y(n_742) );
INVx4_ASAP7_75t_L g743 ( .A(n_653), .Y(n_743) );
BUFx3_ASAP7_75t_L g744 ( .A(n_653), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_567), .B(n_574), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_567), .B(n_574), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_621), .B(n_543), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_740), .B(n_687), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_741), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_666), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_731), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_715), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_715), .Y(n_753) );
OR2x6_ASAP7_75t_L g754 ( .A(n_681), .B(n_731), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_721), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_671), .B(n_664), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_680), .B(n_700), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_722), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_731), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_707), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_747), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_665), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_666), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_672), .A2(n_676), .B(n_725), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_673), .Y(n_765) );
BUFx12f_ASAP7_75t_L g766 ( .A(n_692), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_673), .Y(n_767) );
BUFx3_ASAP7_75t_L g768 ( .A(n_670), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_739), .Y(n_769) );
OA21x2_ASAP7_75t_L g770 ( .A1(n_672), .A2(n_676), .B(n_724), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_739), .Y(n_771) );
BUFx3_ASAP7_75t_L g772 ( .A(n_670), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_745), .B(n_746), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_717), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_746), .B(n_686), .Y(n_775) );
AO21x2_ASAP7_75t_L g776 ( .A1(n_719), .A2(n_708), .B(n_718), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_718), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_668), .B(n_727), .Y(n_778) );
AND2x4_ASAP7_75t_L g779 ( .A(n_689), .B(n_674), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_744), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_733), .B(n_688), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_738), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_698), .B(n_678), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_728), .A2(n_734), .B1(n_683), .B2(n_688), .Y(n_784) );
BUFx3_ASAP7_75t_L g785 ( .A(n_737), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_689), .B(n_677), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_720), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_726), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_704), .A2(n_703), .B1(n_669), .B2(n_711), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_697), .B(n_679), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_726), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_733), .B(n_703), .Y(n_792) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_685), .Y(n_793) );
INVx2_ASAP7_75t_SL g794 ( .A(n_667), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_684), .Y(n_795) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_667), .B(n_743), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_736), .B(n_729), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g798 ( .A(n_693), .B(n_710), .C(n_691), .D(n_730), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_696), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_694), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_743), .Y(n_801) );
INVx4_ASAP7_75t_L g802 ( .A(n_705), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_768), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_759), .B(n_695), .Y(n_804) );
OR2x2_ASAP7_75t_L g805 ( .A(n_792), .B(n_690), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_762), .B(n_695), .Y(n_806) );
INVxp67_ASAP7_75t_R g807 ( .A(n_801), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_773), .B(n_716), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_762), .B(n_712), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_760), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_751), .Y(n_811) );
INVx2_ASAP7_75t_SL g812 ( .A(n_754), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_787), .B(n_713), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_749), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_759), .B(n_723), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_765), .B(n_723), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_787), .B(n_723), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_783), .B(n_699), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_792), .B(n_699), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_765), .B(n_706), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_768), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_761), .Y(n_822) );
BUFx3_ASAP7_75t_L g823 ( .A(n_772), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_783), .B(n_735), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_790), .B(n_752), .Y(n_825) );
BUFx3_ASAP7_75t_L g826 ( .A(n_772), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_799), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_757), .A2(n_714), .B1(n_709), .B2(n_732), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_793), .Y(n_829) );
NOR2x1p5_ASAP7_75t_L g830 ( .A(n_785), .B(n_742), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_790), .B(n_682), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_767), .B(n_737), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_752), .B(n_702), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_781), .B(n_701), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_777), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_753), .B(n_675), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_767), .B(n_701), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_755), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_758), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_769), .B(n_701), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_798), .B(n_756), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_758), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_775), .A2(n_789), .B1(n_784), .B2(n_748), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_778), .B(n_782), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_778), .B(n_782), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_779), .B(n_786), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_779), .B(n_786), .Y(n_847) );
AND2x4_ASAP7_75t_L g848 ( .A(n_754), .B(n_779), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_794), .Y(n_849) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_797), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_750), .Y(n_851) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_769), .Y(n_852) );
HB1xp67_ASAP7_75t_SL g853 ( .A(n_750), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_849), .Y(n_854) );
BUFx2_ASAP7_75t_L g855 ( .A(n_852), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_825), .B(n_788), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_825), .B(n_788), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_846), .B(n_791), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_846), .B(n_791), .Y(n_859) );
INVx1_ASAP7_75t_SL g860 ( .A(n_853), .Y(n_860) );
AND2x2_ASAP7_75t_SL g861 ( .A(n_848), .B(n_811), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_810), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_849), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_810), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_847), .B(n_764), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_827), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_805), .B(n_781), .Y(n_867) );
NAND2x1p5_ASAP7_75t_L g868 ( .A(n_803), .B(n_796), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_844), .B(n_771), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_829), .Y(n_870) );
INVx2_ASAP7_75t_SL g871 ( .A(n_848), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_814), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_844), .B(n_776), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_845), .B(n_776), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_845), .B(n_776), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_817), .B(n_764), .Y(n_876) );
AND2x4_ASAP7_75t_SL g877 ( .A(n_848), .B(n_802), .Y(n_877) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_853), .Y(n_878) );
BUFx8_ASAP7_75t_SL g879 ( .A(n_832), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_817), .B(n_795), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g881 ( .A(n_803), .B(n_794), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_803), .Y(n_882) );
INVx2_ASAP7_75t_SL g883 ( .A(n_848), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_822), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_804), .Y(n_885) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_854), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_873), .B(n_838), .Y(n_887) );
NAND2x1p5_ASAP7_75t_L g888 ( .A(n_855), .B(n_821), .Y(n_888) );
XNOR2x1_ASAP7_75t_L g889 ( .A(n_860), .B(n_830), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_865), .B(n_815), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_862), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_856), .B(n_850), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_865), .B(n_815), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_873), .B(n_816), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_863), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_874), .B(n_875), .Y(n_896) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_855), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_879), .B(n_785), .Y(n_898) );
INVx3_ASAP7_75t_L g899 ( .A(n_885), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_874), .B(n_816), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_856), .B(n_808), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_857), .B(n_808), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_862), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_858), .B(n_839), .Y(n_904) );
INVxp67_ASAP7_75t_L g905 ( .A(n_866), .Y(n_905) );
OR2x2_ASAP7_75t_L g906 ( .A(n_875), .B(n_806), .Y(n_906) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_870), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_864), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_859), .B(n_839), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_857), .B(n_813), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_859), .B(n_842), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_867), .B(n_806), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_872), .B(n_813), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_864), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_876), .B(n_842), .Y(n_915) );
INVx3_ASAP7_75t_SL g916 ( .A(n_860), .Y(n_916) );
INVx1_ASAP7_75t_SL g917 ( .A(n_882), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_885), .B(n_812), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_884), .B(n_841), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_869), .B(n_835), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_880), .B(n_770), .Y(n_921) );
INVx1_ASAP7_75t_SL g922 ( .A(n_889), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_897), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_915), .B(n_869), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_886), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_898), .B(n_766), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_921), .B(n_871), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_891), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_921), .B(n_871), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_919), .A2(n_818), .B1(n_824), .B2(n_831), .Y(n_930) );
NOR2xp67_ASAP7_75t_L g931 ( .A(n_899), .B(n_766), .Y(n_931) );
OAI222xp33_ASAP7_75t_L g932 ( .A1(n_888), .A2(n_878), .B1(n_882), .B2(n_871), .C1(n_883), .C2(n_828), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g933 ( .A1(n_907), .A2(n_828), .B(n_878), .C(n_843), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_891), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_903), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_889), .A2(n_861), .B1(n_807), .B2(n_877), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_905), .B(n_836), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_903), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_908), .Y(n_939) );
AOI32xp33_ASAP7_75t_L g940 ( .A1(n_904), .A2(n_836), .A3(n_877), .B1(n_800), .B2(n_833), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_913), .B(n_774), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_908), .Y(n_942) );
NAND2x1p5_ASAP7_75t_L g943 ( .A(n_917), .B(n_881), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_890), .B(n_883), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_892), .B(n_774), .Y(n_945) );
A2O1A1Ixp33_ASAP7_75t_L g946 ( .A1(n_918), .A2(n_877), .B(n_861), .C(n_826), .Y(n_946) );
AND2x4_ASAP7_75t_L g947 ( .A(n_899), .B(n_883), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_914), .Y(n_948) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_936), .A2(n_916), .B1(n_807), .B2(n_888), .Y(n_949) );
O2A1O1Ixp5_ASAP7_75t_L g950 ( .A1(n_932), .A2(n_887), .B(n_899), .C(n_920), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_923), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_928), .B(n_896), .Y(n_952) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_925), .Y(n_953) );
NOR2x1_ASAP7_75t_L g954 ( .A(n_946), .B(n_830), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_924), .B(n_896), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_927), .B(n_910), .Y(n_956) );
AO22x1_ASAP7_75t_L g957 ( .A1(n_922), .A2(n_916), .B1(n_895), .B2(n_917), .Y(n_957) );
NOR3xp33_ASAP7_75t_L g958 ( .A(n_933), .B(n_832), .C(n_837), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_937), .A2(n_818), .B1(n_824), .B2(n_831), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_930), .A2(n_915), .B1(n_893), .B2(n_890), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_927), .B(n_906), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_928), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_934), .B(n_904), .Y(n_963) );
INVxp33_ASAP7_75t_L g964 ( .A(n_926), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_940), .B(n_895), .C(n_887), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_929), .B(n_909), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_941), .B(n_916), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_929), .B(n_909), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_953), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_954), .A2(n_946), .B1(n_931), .B2(n_861), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g971 ( .A1(n_950), .A2(n_945), .B1(n_833), .B2(n_942), .C(n_939), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_958), .A2(n_948), .B1(n_938), .B2(n_935), .C(n_901), .Y(n_972) );
NAND2xp5_ASAP7_75t_SL g973 ( .A(n_949), .B(n_943), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_952), .Y(n_974) );
OAI322xp33_ASAP7_75t_L g975 ( .A1(n_960), .A2(n_894), .A3(n_900), .B1(n_902), .B2(n_906), .C1(n_819), .C2(n_912), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_961), .B(n_944), .Y(n_976) );
INVxp67_ASAP7_75t_L g977 ( .A(n_951), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g978 ( .A1(n_965), .A2(n_943), .B1(n_888), .B2(n_899), .C(n_900), .Y(n_978) );
AOI21xp33_ASAP7_75t_L g979 ( .A1(n_964), .A2(n_819), .B(n_809), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_962), .Y(n_980) );
UNKNOWN g981 ( );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_967), .B(n_944), .Y(n_982) );
AOI21xp5_ASAP7_75t_L g983 ( .A1(n_957), .A2(n_947), .B(n_943), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_963), .B(n_911), .Y(n_984) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_963), .Y(n_985) );
NOR2xp33_ASAP7_75t_SL g986 ( .A(n_956), .B(n_780), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_955), .B(n_911), .Y(n_987) );
NAND3xp33_ASAP7_75t_SL g988 ( .A(n_966), .B(n_868), .C(n_834), .Y(n_988) );
NAND3xp33_ASAP7_75t_L g989 ( .A(n_968), .B(n_809), .C(n_837), .Y(n_989) );
OAI211xp5_ASAP7_75t_SL g990 ( .A1(n_971), .A2(n_973), .B(n_978), .C(n_970), .Y(n_990) );
AOI211xp5_ASAP7_75t_L g991 ( .A1(n_971), .A2(n_983), .B(n_988), .C(n_975), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_972), .B(n_977), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_977), .B(n_985), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g994 ( .A(n_985), .B(n_969), .Y(n_994) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_986), .A2(n_972), .B1(n_989), .B2(n_974), .Y(n_995) );
NOR2x1_ASAP7_75t_L g996 ( .A(n_990), .B(n_780), .Y(n_996) );
NOR2x1_ASAP7_75t_L g997 ( .A(n_992), .B(n_796), .Y(n_997) );
NAND4xp25_ASAP7_75t_L g998 ( .A(n_991), .B(n_840), .C(n_981), .D(n_979), .Y(n_998) );
NOR3xp33_ASAP7_75t_L g999 ( .A(n_993), .B(n_840), .C(n_982), .Y(n_999) );
AND3x1_ASAP7_75t_L g1000 ( .A(n_996), .B(n_994), .C(n_995), .Y(n_1000) );
OR4x2_ASAP7_75t_L g1001 ( .A(n_998), .B(n_976), .C(n_987), .D(n_984), .Y(n_1001) );
NOR3xp33_ASAP7_75t_L g1002 ( .A(n_997), .B(n_820), .C(n_763), .Y(n_1002) );
NAND4xp75_ASAP7_75t_L g1003 ( .A(n_1000), .B(n_999), .C(n_763), .D(n_820), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_1001), .Y(n_1004) );
XNOR2xp5_ASAP7_75t_L g1005 ( .A(n_1004), .B(n_1002), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_1003), .Y(n_1006) );
OAI22x1_ASAP7_75t_SL g1007 ( .A1(n_1005), .A2(n_1003), .B1(n_980), .B2(n_802), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1006), .Y(n_1008) );
INVxp67_ASAP7_75t_L g1009 ( .A(n_1008), .Y(n_1009) );
OR2x6_ASAP7_75t_L g1010 ( .A(n_1009), .B(n_1007), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_1010), .A2(n_826), .B1(n_823), .B2(n_821), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_1011), .A2(n_947), .B(n_851), .Y(n_1012) );
endmodule