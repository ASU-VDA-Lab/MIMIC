module fake_ariane_1337_n_194 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_194);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_194;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_30;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVxp33_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_R g52 ( 
.A(n_31),
.B(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_4),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_4),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_R g61 ( 
.A(n_49),
.B(n_5),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx11_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2x1p5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_45),
.B1(n_28),
.B2(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_46),
.Y(n_80)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_33),
.B1(n_43),
.B2(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_34),
.C(n_28),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_34),
.Y(n_84)
);

OAI221xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_33),
.B1(n_43),
.B2(n_41),
.C(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_36),
.B(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_72),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_36),
.B(n_51),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_74),
.B(n_86),
.C(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_56),
.C(n_64),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_65),
.Y(n_97)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_59),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_61),
.C(n_85),
.D(n_60),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_94),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_83),
.B(n_54),
.C(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2x1_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_99),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_100),
.B1(n_97),
.B2(n_90),
.C(n_96),
.Y(n_110)
);

OAI222xp33_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_70),
.B1(n_67),
.B2(n_54),
.C1(n_104),
.C2(n_102),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_91),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OR2x6_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_81),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_81),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_98),
.B(n_108),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_103),
.B1(n_73),
.B2(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

OAI211xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_107),
.B(n_101),
.C(n_37),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_107),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_115),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_115),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_114),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_114),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_81),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_32),
.Y(n_134)
);

AOI33xp33_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_32),
.A3(n_44),
.B1(n_41),
.B2(n_38),
.B3(n_37),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_29),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_87),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_29),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_127),
.B(n_125),
.C(n_30),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_127),
.B(n_73),
.C(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_130),
.B1(n_131),
.B2(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_125),
.C(n_30),
.Y(n_147)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_144),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_148),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_44),
.B(n_131),
.C(n_122),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_122),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_126),
.C(n_92),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_122),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_126),
.Y(n_157)
);

OAI211xp5_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_139),
.B(n_86),
.C(n_11),
.Y(n_158)
);

OAI211xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_139),
.B(n_10),
.C(n_12),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_9),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_10),
.B(n_13),
.Y(n_162)
);

AOI221x1_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_126),
.B1(n_133),
.B2(n_108),
.C(n_82),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_52),
.B1(n_73),
.B2(n_17),
.C(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_165),
.B(n_161),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_154),
.A3(n_157),
.B1(n_150),
.B2(n_129),
.C(n_124),
.Y(n_168)
);

AND3x4_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_154),
.C(n_15),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_52),
.B1(n_123),
.B2(n_82),
.C(n_87),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_158),
.B1(n_123),
.B2(n_129),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_14),
.Y(n_173)
);

OAI321xp33_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_124),
.A3(n_88),
.B1(n_87),
.B2(n_17),
.C(n_99),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_SL g175 ( 
.A(n_172),
.B(n_124),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_171),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_105),
.B(n_88),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_170),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_18),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_176),
.B1(n_181),
.B2(n_177),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_175),
.B1(n_180),
.B2(n_75),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

OAI211xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_182),
.B(n_184),
.C(n_180),
.Y(n_191)
);

OAI211xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_182),
.B(n_175),
.C(n_95),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_105),
.B1(n_98),
.B2(n_20),
.Y(n_193)
);

AOI221xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_190),
.B1(n_192),
.B2(n_98),
.C(n_23),
.Y(n_194)
);


endmodule