module fake_jpeg_1317_n_421 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_55),
.Y(n_121)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_58),
.B(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_66),
.Y(n_120)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_70),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_71),
.B(n_89),
.Y(n_177)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_81),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_83),
.B(n_84),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_8),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_25),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_102),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_10),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_107),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_26),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_101),
.B(n_103),
.Y(n_153)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_26),
.B(n_6),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_106),
.B(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_111),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_28),
.B(n_11),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_16),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_28),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_16),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_112),
.A2(n_118),
.B1(n_162),
.B2(n_174),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_33),
.B1(n_40),
.B2(n_48),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_36),
.B1(n_44),
.B2(n_22),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_22),
.B1(n_46),
.B2(n_45),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_68),
.A2(n_22),
.B1(n_46),
.B2(n_43),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_31),
.B1(n_43),
.B2(n_39),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_159),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_30),
.B1(n_39),
.B2(n_38),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_40),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_140),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_48),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_77),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_142),
.A2(n_149),
.B1(n_151),
.B2(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_155),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_37),
.B(n_42),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_145),
.B(n_120),
.C(n_123),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_63),
.B(n_1),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_2),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_156),
.B(n_158),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_11),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_80),
.A2(n_13),
.B(n_15),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_87),
.A2(n_3),
.B1(n_16),
.B2(n_96),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_171),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_54),
.A2(n_3),
.B1(n_72),
.B2(n_92),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_82),
.A2(n_105),
.B1(n_107),
.B2(n_73),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_166),
.A2(n_173),
.B1(n_178),
.B2(n_182),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_69),
.A2(n_111),
.B1(n_109),
.B2(n_106),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_169),
.A2(n_132),
.B1(n_134),
.B2(n_167),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_109),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_80),
.A2(n_23),
.B1(n_47),
.B2(n_20),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_58),
.A2(n_55),
.B1(n_53),
.B2(n_81),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_161),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_58),
.A2(n_55),
.B1(n_53),
.B2(n_81),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_140),
.B1(n_144),
.B2(n_128),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_76),
.A2(n_23),
.B1(n_47),
.B2(n_20),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_76),
.A2(n_23),
.B1(n_47),
.B2(n_20),
.Y(n_182)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_205),
.Y(n_244)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_197),
.B(n_208),
.Y(n_245)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_146),
.B(n_148),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_198),
.B(n_230),
.Y(n_271)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_202),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_204),
.B(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_114),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_153),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_114),
.B(n_127),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_233),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_138),
.B(n_145),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_215),
.B(n_217),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_143),
.A2(n_147),
.B1(n_183),
.B2(n_130),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_237),
.B1(n_214),
.B2(n_199),
.Y(n_261)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_169),
.A2(n_154),
.B1(n_172),
.B2(n_117),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_234),
.B1(n_116),
.B2(n_165),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_158),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_167),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_223),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_227),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_225),
.Y(n_282)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_120),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_232),
.Y(n_278)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_135),
.A2(n_180),
.B1(n_139),
.B2(n_116),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_123),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_150),
.B(n_168),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_132),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_168),
.A2(n_141),
.B1(n_117),
.B2(n_179),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_243),
.B1(n_209),
.B2(n_240),
.Y(n_280)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_219),
.B1(n_185),
.B2(n_235),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_205),
.B(n_165),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_261),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_152),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_259),
.C(n_212),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_186),
.B(n_215),
.C(n_193),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_252),
.B(n_264),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_190),
.A2(n_179),
.B1(n_135),
.B2(n_139),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_257),
.A2(n_277),
.B1(n_279),
.B2(n_246),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_184),
.B(n_152),
.CI(n_180),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_216),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_195),
.B(n_211),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_186),
.A2(n_198),
.B(n_201),
.C(n_207),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_203),
.A2(n_201),
.B(n_241),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_271),
.B(n_264),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_192),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_232),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_243),
.B1(n_228),
.B2(n_191),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_229),
.A2(n_196),
.B1(n_187),
.B2(n_188),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_225),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_285),
.B(n_299),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_288),
.C(n_268),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_302),
.B1(n_308),
.B2(n_276),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_194),
.C(n_200),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_291),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_235),
.B1(n_236),
.B2(n_224),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_297),
.B1(n_262),
.B2(n_308),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_244),
.B(n_236),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_224),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_295),
.B(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_216),
.B1(n_259),
.B2(n_266),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_216),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_301),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_247),
.A2(n_250),
.B1(n_277),
.B2(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_271),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_248),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_306),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_272),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_314),
.B(n_316),
.Y(n_329)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_249),
.B(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_322),
.A2(n_327),
.B1(n_333),
.B2(n_298),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_267),
.B(n_276),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_338),
.B(n_341),
.C(n_305),
.Y(n_350)
);

AO22x1_ASAP7_75t_L g330 ( 
.A1(n_302),
.A2(n_258),
.B1(n_247),
.B2(n_254),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_305),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_279),
.B(n_265),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_331),
.B(n_315),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_298),
.A2(n_265),
.B1(n_282),
.B2(n_253),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_268),
.B(n_254),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_292),
.C(n_284),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_297),
.B(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_347),
.B1(n_349),
.B2(n_352),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_305),
.C(n_286),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_344),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_332),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_346),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_336),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_336),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_283),
.B1(n_284),
.B2(n_293),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_325),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_359),
.B1(n_340),
.B2(n_324),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_316),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_355),
.B1(n_360),
.B2(n_326),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_326),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_357),
.C(n_338),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_291),
.C(n_300),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_323),
.B(n_331),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_358),
.B(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_263),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_304),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_333),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_368),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_341),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_369),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_328),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_373),
.C(n_361),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_328),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_358),
.B(n_330),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_348),
.C(n_289),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_355),
.A2(n_320),
.B1(n_322),
.B2(n_337),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_347),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_320),
.B1(n_337),
.B2(n_334),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_376),
.B(n_334),
.Y(n_382)
);

FAx1_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_335),
.CI(n_329),
.CON(n_377),
.SN(n_377)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_329),
.B(n_342),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_346),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_379),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_380),
.A2(n_382),
.B1(n_386),
.B2(n_371),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_377),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_384),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_367),
.B(n_325),
.Y(n_384)
);

NOR3xp33_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_350),
.C(n_348),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_365),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_381),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_391),
.B(n_396),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_393),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_370),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_395),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_373),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_364),
.C(n_372),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_385),
.C(n_389),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_399),
.B(n_404),
.Y(n_410)
);

AOI321xp33_ASAP7_75t_L g400 ( 
.A1(n_390),
.A2(n_377),
.A3(n_386),
.B1(n_362),
.B2(n_359),
.C(n_379),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_401),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_374),
.C(n_368),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_319),
.C(n_318),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_405),
.A2(n_398),
.B1(n_312),
.B2(n_324),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_406),
.A2(n_409),
.B1(n_312),
.B2(n_318),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_393),
.B(n_397),
.Y(n_407)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_407),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_SL g409 ( 
.A(n_403),
.B(n_395),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_410),
.B(n_408),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_413),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_406),
.B(n_402),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_354),
.B1(n_290),
.B2(n_287),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_411),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_417),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_416),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_419),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_418),
.Y(n_421)
);


endmodule