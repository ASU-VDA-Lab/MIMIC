module fake_ariane_2815_n_1199 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1199);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1199;

wire n_556;
wire n_356;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_1187;
wire n_985;
wire n_421;
wire n_1167;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_1180;
wire n_969;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_1184;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_336;
wire n_665;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_402;
wire n_1068;
wire n_1052;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_1185;
wire n_485;
wire n_401;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_721;
wire n_433;
wire n_481;
wire n_426;
wire n_600;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_1153;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_369;
wire n_1192;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_1172;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_1160;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_654;
wire n_429;
wire n_455;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_1188;
wire n_539;
wire n_1150;
wire n_728;
wire n_388;
wire n_333;
wire n_612;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_459;
wire n_321;
wire n_911;
wire n_1136;
wire n_458;
wire n_361;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_1194;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_1135;
wire n_888;
wire n_918;
wire n_639;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_551;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_571;
wire n_414;
wire n_680;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_666;
wire n_1000;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_746;
wire n_456;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_615;
wire n_1070;
wire n_1027;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g314 ( 
.A(n_91),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_0),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_310),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_104),
.B(n_99),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_112),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_229),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_6),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_115),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_202),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_136),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_135),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_5),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_199),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_59),
.B(n_89),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_81),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_114),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_76),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_149),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_46),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_79),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_133),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_52),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_95),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_176),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_13),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_254),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_282),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_289),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_248),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_145),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_131),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_73),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_204),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_34),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_34),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_118),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_64),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_252),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_235),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_158),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_236),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_228),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_62),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_18),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_103),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_170),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_243),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_166),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_172),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_301),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_85),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_223),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_65),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_261),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_192),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_302),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_124),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_222),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_77),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_183),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_196),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_290),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_187),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_299),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_116),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_249),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_181),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_210),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_120),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_185),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_123),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_241),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_127),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_110),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_201),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_107),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_258),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_264),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_182),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_68),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_72),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_303),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_60),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_96),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_178),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_93),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_209),
.B(n_286),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_43),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_105),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_230),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_6),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_1),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_70),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_188),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_263),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_22),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_100),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_4),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_13),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_82),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_280),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_208),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_50),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_300),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_140),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_279),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_27),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_67),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_4),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_285),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_311),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_71),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_92),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_220),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_142),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_10),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_179),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_224),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_233),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_306),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_106),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_259),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_152),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_205),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_74),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_270),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_9),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_238),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_217),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_281),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_295),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_195),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_277),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_121),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_49),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_117),
.Y(n_466)
);

BUFx8_ASAP7_75t_SL g467 ( 
.A(n_168),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_113),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_273),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_206),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_90),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_274),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_255),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_22),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_276),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_130),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_66),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_251),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_21),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_3),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_54),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_153),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_422),
.B(n_0),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_355),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_323),
.B(n_1),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_355),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_434),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_387),
.B(n_2),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_315),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_341),
.A2(n_42),
.B(n_41),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_445),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_7),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_8),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_370),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_320),
.A2(n_352),
.B1(n_364),
.B2(n_362),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_355),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_316),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_329),
.B(n_11),
.Y(n_503)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_314),
.A2(n_11),
.B(n_12),
.Y(n_504)
);

OAI22x1_ASAP7_75t_SL g505 ( 
.A1(n_424),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_14),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_405),
.B(n_44),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_383),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_365),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_315),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_348),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_332),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_321),
.B(n_16),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_358),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

OAI22x1_ASAP7_75t_R g516 ( 
.A1(n_357),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_443),
.B(n_19),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_326),
.B(n_20),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_436),
.B(n_21),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_348),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_444),
.B(n_23),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_454),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_391),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_384),
.A2(n_478),
.B1(n_433),
.B2(n_368),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_405),
.B(n_45),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_467),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_328),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_418),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_405),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_334),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_23),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_427),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_385),
.B(n_24),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_442),
.B(n_24),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_350),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_335),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_350),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_336),
.Y(n_546)
);

AOI22x1_ASAP7_75t_SL g547 ( 
.A1(n_338),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

NOR2x1_ASAP7_75t_L g549 ( 
.A(n_340),
.B(n_47),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_318),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_337),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_337),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_342),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_458),
.B(n_32),
.Y(n_556)
);

INVxp33_ASAP7_75t_SL g557 ( 
.A(n_317),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_343),
.B(n_33),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_344),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_346),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_354),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_360),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_319),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_324),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_446),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_369),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_378),
.B(n_35),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_469),
.B(n_36),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_379),
.B(n_37),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_381),
.A2(n_173),
.B(n_312),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_388),
.B(n_38),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

INVx8_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_489),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_541),
.B(n_322),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_485),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g583 ( 
.A1(n_483),
.A2(n_392),
.B(n_390),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_461),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_571),
.B(n_325),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_488),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_488),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_511),
.B(n_396),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_518),
.B(n_399),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_400),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_533),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_518),
.B(n_563),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_517),
.B(n_331),
.Y(n_605)
);

BUFx6f_ASAP7_75t_SL g606 ( 
.A(n_510),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_529),
.B(n_438),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_571),
.Y(n_608)
);

INVxp33_ASAP7_75t_L g609 ( 
.A(n_536),
.Y(n_609)
);

NOR2x1p5_ASAP7_75t_L g610 ( 
.A(n_530),
.B(n_401),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_538),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_538),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_574),
.B(n_482),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_542),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_487),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_574),
.B(n_327),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_540),
.B(n_375),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_491),
.B(n_481),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_527),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_508),
.B(n_402),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_557),
.B(n_407),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_565),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_565),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_526),
.B(n_414),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_531),
.B(n_415),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_508),
.B(n_419),
.Y(n_638)
);

INVx8_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

BUFx6f_ASAP7_75t_SL g641 ( 
.A(n_484),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_567),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_570),
.Y(n_644)
);

BUFx6f_ASAP7_75t_SL g645 ( 
.A(n_484),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_555),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_506),
.B(n_477),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_556),
.B(n_569),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_570),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_545),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_543),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_631),
.B(n_496),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_561),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_585),
.B(n_513),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_631),
.B(n_499),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_619),
.A2(n_551),
.B1(n_544),
.B2(n_509),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_622),
.B(n_534),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_608),
.B(n_537),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_578),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_605),
.A2(n_521),
.B1(n_523),
.B2(n_503),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_654),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_585),
.B(n_546),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_592),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_644),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_646),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_649),
.A2(n_521),
.B1(n_523),
.B2(n_503),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_648),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_585),
.B(n_562),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_585),
.B(n_566),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_650),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_585),
.B(n_573),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_586),
.B(n_560),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_593),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_579),
.A2(n_558),
.B1(n_495),
.B2(n_564),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_584),
.B(n_535),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_587),
.B(n_535),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_608),
.B(n_497),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_630),
.B(n_497),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_652),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_627),
.B(n_647),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_649),
.B(n_539),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_618),
.B(n_627),
.Y(n_691)
);

INVxp67_ASAP7_75t_SL g692 ( 
.A(n_618),
.Y(n_692)
);

AOI221xp5_ASAP7_75t_L g693 ( 
.A1(n_614),
.A2(n_552),
.B1(n_554),
.B2(n_505),
.C(n_575),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_576),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_638),
.B(n_520),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_636),
.B(n_545),
.Y(n_696)
);

BUFx5_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_636),
.B(n_553),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_635),
.B(n_553),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_609),
.B(n_568),
.Y(n_700)
);

AND2x2_ASAP7_75t_SL g701 ( 
.A(n_619),
.B(n_500),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_590),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_602),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_647),
.B(n_579),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_652),
.Y(n_705)
);

OAI22x1_ASAP7_75t_R g706 ( 
.A1(n_629),
.A2(n_516),
.B1(n_547),
.B2(n_432),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_625),
.B(n_504),
.C(n_549),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_597),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_603),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_635),
.B(n_421),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_601),
.B(n_539),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_613),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_588),
.B(n_539),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_588),
.B(n_550),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_614),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_623),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_617),
.B(n_550),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_617),
.B(n_550),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_609),
.B(n_504),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_606),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_576),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_621),
.B(n_435),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_621),
.B(n_437),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_639),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_653),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_596),
.B(n_330),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_639),
.B(n_507),
.Y(n_729)
);

XNOR2xp5_ASAP7_75t_L g730 ( 
.A(n_607),
.B(n_547),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_610),
.A2(n_572),
.B(n_470),
.C(n_439),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_R g732 ( 
.A(n_598),
.B(n_493),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_641),
.B(n_440),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_581),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_582),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_682),
.B(n_639),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_660),
.A2(n_645),
.B1(n_641),
.B2(n_453),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_695),
.A2(n_463),
.B(n_460),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_657),
.A2(n_466),
.B(n_472),
.C(n_464),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_715),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_675),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_694),
.B(n_637),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_707),
.A2(n_583),
.B(n_475),
.Y(n_744)
);

AOI221x1_ASAP7_75t_SL g745 ( 
.A1(n_663),
.A2(n_703),
.B1(n_702),
.B2(n_674),
.C(n_678),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_724),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_659),
.A2(n_476),
.B(n_473),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_667),
.A2(n_645),
.B1(n_456),
.B2(n_451),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_704),
.A2(n_339),
.B(n_333),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_731),
.A2(n_347),
.B(n_345),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_711),
.A2(n_351),
.B(n_349),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_690),
.A2(n_356),
.B(n_353),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_660),
.B(n_637),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_673),
.A2(n_431),
.B1(n_361),
.B2(n_363),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_725),
.B(n_359),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_664),
.B(n_366),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_675),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_727),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_655),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_721),
.B(n_367),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_656),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_691),
.A2(n_372),
.B(n_371),
.Y(n_763)
);

AOI21xp33_ASAP7_75t_L g764 ( 
.A1(n_692),
.A2(n_374),
.B(n_373),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_683),
.B(n_376),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_665),
.A2(n_380),
.B(n_377),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_709),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_700),
.A2(n_393),
.B(n_382),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_658),
.A2(n_397),
.B(n_395),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_696),
.B(n_398),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_403),
.Y(n_771)
);

OAI21xp33_ASAP7_75t_L g772 ( 
.A1(n_710),
.A2(n_408),
.B(n_406),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_710),
.A2(n_413),
.B(n_616),
.C(n_611),
.Y(n_773)
);

AO21x2_ASAP7_75t_L g774 ( 
.A1(n_707),
.A2(n_651),
.B(n_591),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_732),
.A2(n_658),
.B(n_714),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_668),
.B(n_606),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_686),
.A2(n_465),
.B1(n_410),
.B2(n_411),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_729),
.B(n_409),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_684),
.A2(n_416),
.B(n_412),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_675),
.B(n_612),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_698),
.A2(n_528),
.B(n_507),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_698),
.B(n_420),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_723),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_685),
.A2(n_426),
.B(n_423),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_699),
.B(n_428),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_680),
.A2(n_634),
.B(n_643),
.C(n_642),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_680),
.A2(n_651),
.B(n_643),
.C(n_642),
.Y(n_787)
);

AOI21xp33_ASAP7_75t_L g788 ( 
.A1(n_669),
.A2(n_430),
.B(n_429),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_729),
.A2(n_441),
.B1(n_448),
.B2(n_449),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_687),
.B(n_450),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_713),
.A2(n_452),
.B1(n_455),
.B2(n_459),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_662),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_733),
.A2(n_640),
.B(n_633),
.C(n_628),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_726),
.B(n_462),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_718),
.A2(n_468),
.B(n_589),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_722),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_712),
.B(n_717),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_719),
.B(n_38),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_728),
.A2(n_666),
.B(n_661),
.Y(n_800)
);

BUFx8_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_661),
.A2(n_591),
.B(n_589),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_676),
.A2(n_677),
.B1(n_699),
.B2(n_679),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_670),
.A2(n_595),
.B(n_594),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_671),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_681),
.A2(n_595),
.B(n_594),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_697),
.B(n_39),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_697),
.B(n_599),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_688),
.A2(n_528),
.B(n_507),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_705),
.A2(n_600),
.B(n_599),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_697),
.A2(n_528),
.B1(n_507),
.B2(n_628),
.Y(n_812)
);

BUFx8_ASAP7_75t_L g813 ( 
.A(n_697),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_693),
.A2(n_640),
.B1(n_633),
.B2(n_626),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_734),
.A2(n_626),
.B(n_624),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_720),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_735),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_746),
.A2(n_736),
.B(n_735),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_807),
.B(n_735),
.C(n_708),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_744),
.A2(n_620),
.B(n_600),
.Y(n_820)
);

AOI21xp33_ASAP7_75t_L g821 ( 
.A1(n_748),
.A2(n_706),
.B(n_624),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_787),
.A2(n_528),
.B(n_708),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_SL g823 ( 
.A(n_756),
.B(n_620),
.C(n_40),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_738),
.B(n_697),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_745),
.A2(n_708),
.B(n_604),
.C(n_597),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_776),
.B(n_789),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_763),
.B(n_708),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_808),
.A2(n_604),
.B(n_597),
.Y(n_828)
);

OA22x2_ASAP7_75t_L g829 ( 
.A1(n_810),
.A2(n_39),
.B1(n_40),
.B2(n_375),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_809),
.A2(n_375),
.B(n_51),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_760),
.B(n_604),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_747),
.A2(n_375),
.B(n_53),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_800),
.A2(n_604),
.B(n_375),
.Y(n_833)
);

AO21x2_ASAP7_75t_L g834 ( 
.A1(n_775),
.A2(n_375),
.B(n_55),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_802),
.A2(n_48),
.B(n_56),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_803),
.A2(n_57),
.B(n_58),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_815),
.A2(n_61),
.B(n_63),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_761),
.A2(n_69),
.B(n_75),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_770),
.B(n_78),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_785),
.A2(n_782),
.B(n_771),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_817),
.B(n_80),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_750),
.A2(n_83),
.B(n_84),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_739),
.A2(n_86),
.B(n_87),
.Y(n_843)
);

AO31x2_ASAP7_75t_L g844 ( 
.A1(n_773),
.A2(n_88),
.A3(n_94),
.B(n_97),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_798),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_755),
.B(n_98),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_758),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_799),
.A2(n_101),
.B(n_102),
.C(n_108),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_737),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_741),
.A2(n_109),
.B1(n_111),
.B2(n_119),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_790),
.B(n_122),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_749),
.A2(n_781),
.B(n_769),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_793),
.A2(n_786),
.B(n_795),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_753),
.A2(n_125),
.B(n_126),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_783),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_804),
.A2(n_806),
.B(n_811),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_752),
.A2(n_128),
.B(n_129),
.Y(n_857)
);

CKINVDCx8_ASAP7_75t_R g858 ( 
.A(n_780),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_765),
.A2(n_772),
.B(n_740),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_812),
.A2(n_132),
.B(n_134),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_797),
.B(n_780),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_751),
.A2(n_137),
.B(n_138),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_817),
.A2(n_139),
.B(n_141),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_742),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_794),
.A2(n_143),
.B(n_144),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_774),
.A2(n_146),
.B(n_147),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_813),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_780),
.B(n_148),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_757),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_779),
.A2(n_150),
.B(n_151),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_774),
.A2(n_154),
.B(n_155),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_L g872 ( 
.A1(n_754),
.A2(n_156),
.B(n_157),
.Y(n_872)
);

BUFx2_ASAP7_75t_SL g873 ( 
.A(n_858),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_855),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_830),
.A2(n_814),
.B(n_778),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_836),
.A2(n_767),
.B(n_759),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_847),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_845),
.B(n_798),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_864),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_861),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_852),
.A2(n_762),
.B(n_792),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_868),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_831),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_868),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_866),
.A2(n_816),
.B(n_784),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_834),
.A2(n_788),
.B(n_764),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_867),
.B(n_805),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_871),
.A2(n_768),
.B(n_766),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_860),
.A2(n_791),
.B(n_743),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_840),
.A2(n_777),
.B(n_796),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_856),
.A2(n_813),
.B(n_161),
.Y(n_891)
);

OAI21x1_ASAP7_75t_SL g892 ( 
.A1(n_859),
.A2(n_801),
.B(n_162),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_820),
.A2(n_160),
.B(n_163),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_826),
.B(n_801),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_869),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_861),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_820),
.A2(n_164),
.B(n_165),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_867),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_861),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_834),
.A2(n_832),
.B(n_819),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_849),
.B(n_167),
.Y(n_901)
);

BUFx12f_ASAP7_75t_L g902 ( 
.A(n_829),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_863),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_851),
.B(n_171),
.Y(n_904)
);

AO21x2_ASAP7_75t_L g905 ( 
.A1(n_819),
.A2(n_853),
.B(n_838),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_825),
.B(n_872),
.C(n_843),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_833),
.A2(n_174),
.B(n_175),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_L g908 ( 
.A1(n_846),
.A2(n_177),
.B(n_180),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_835),
.A2(n_184),
.B(n_186),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_837),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_824),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_839),
.A2(n_189),
.B(n_190),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_844),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_881),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_877),
.Y(n_915)
);

CKINVDCx6p67_ASAP7_75t_R g916 ( 
.A(n_880),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_882),
.B(n_841),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_881),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_876),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_913),
.A2(n_842),
.B(n_828),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_879),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_876),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_896),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_878),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_911),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_882),
.B(n_821),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_883),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_882),
.B(n_844),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_913),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_884),
.B(n_827),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_895),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_887),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_887),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_887),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_911),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_884),
.B(n_841),
.Y(n_936)
);

OAI21x1_ASAP7_75t_SL g937 ( 
.A1(n_892),
.A2(n_870),
.B(n_865),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_884),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_901),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_901),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_901),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_902),
.B(n_844),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_901),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_874),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_911),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_893),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_902),
.A2(n_823),
.B1(n_850),
.B2(n_854),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_898),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_891),
.A2(n_818),
.B(n_862),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_927),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_925),
.B(n_905),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_925),
.B(n_942),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_935),
.B(n_899),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_929),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_928),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_942),
.B(n_905),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_929),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_928),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_926),
.B(n_900),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_915),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_927),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_914),
.Y(n_963)
);

INVxp67_ASAP7_75t_R g964 ( 
.A(n_931),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_SL g965 ( 
.A1(n_923),
.A2(n_894),
.B1(n_896),
.B2(n_895),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_939),
.B(n_899),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_919),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_926),
.B(n_900),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_935),
.B(n_911),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_924),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_919),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_922),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_914),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_918),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_922),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_918),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_944),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_935),
.B(n_898),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_940),
.B(n_873),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_945),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_945),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_945),
.B(n_891),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_946),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_945),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_945),
.B(n_886),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_930),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_941),
.B(n_886),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_947),
.A2(n_890),
.B1(n_906),
.B2(n_904),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_962),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_962),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_955),
.B(n_959),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_988),
.A2(n_943),
.B1(n_923),
.B2(n_930),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_954),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_955),
.B(n_959),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_954),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_982),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_SL g997 ( 
.A1(n_956),
.A2(n_937),
.B1(n_880),
.B2(n_933),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_958),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_958),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_987),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_960),
.B(n_938),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_957),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_987),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_982),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_983),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_983),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_967),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_965),
.A2(n_948),
.B1(n_916),
.B2(n_848),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_961),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_960),
.B(n_946),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_981),
.B(n_903),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_967),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_952),
.B(n_932),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_963),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_950),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_952),
.A2(n_934),
.B1(n_937),
.B2(n_916),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_971),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_963),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_970),
.B(n_917),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_968),
.A2(n_912),
.B(n_908),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_977),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_951),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_951),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_986),
.B(n_917),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_978),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_986),
.B(n_917),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_956),
.A2(n_936),
.B1(n_920),
.B2(n_885),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_981),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_968),
.B(n_920),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_953),
.B(n_936),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_973),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1016),
.A2(n_964),
.B1(n_979),
.B2(n_978),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1020),
.A2(n_992),
.B(n_1008),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_989),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_989),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1021),
.B(n_969),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_991),
.B(n_971),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_991),
.B(n_966),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_990),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_990),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_998),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1002),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1009),
.B(n_969),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_994),
.B(n_985),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_998),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_996),
.B(n_985),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_996),
.B(n_972),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1004),
.B(n_972),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_1022),
.B(n_966),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1004),
.B(n_982),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1001),
.B(n_980),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1013),
.B(n_953),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1023),
.B(n_1010),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_999),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1010),
.B(n_975),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1001),
.Y(n_1057)
);

NOR2x1p5_ASAP7_75t_L g1058 ( 
.A(n_1025),
.B(n_979),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_999),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_993),
.Y(n_1060)
);

INVx3_ASAP7_75t_SL g1061 ( 
.A(n_1028),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1013),
.B(n_953),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_1029),
.B(n_975),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1029),
.B(n_976),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_1025),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1028),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1007),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1057),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1064),
.B(n_1000),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1039),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1033),
.B(n_1053),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1039),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1040),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1032),
.A2(n_997),
.B1(n_1013),
.B2(n_1030),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1054),
.B(n_1000),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_1042),
.B(n_1028),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1041),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1044),
.B(n_964),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1045),
.B(n_1003),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1040),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1041),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1034),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1054),
.B(n_1003),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1035),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1060),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1067),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1046),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1055),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1064),
.B(n_1007),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1059),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1037),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1036),
.B(n_978),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1037),
.Y(n_1093)
);

AOI222xp33_ASAP7_75t_L g1094 ( 
.A1(n_1071),
.A2(n_1020),
.B1(n_1015),
.B2(n_1058),
.C1(n_1019),
.C2(n_1017),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1071),
.A2(n_1043),
.B(n_1024),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1082),
.Y(n_1096)
);

AOI32xp33_ASAP7_75t_L g1097 ( 
.A1(n_1092),
.A2(n_1045),
.A3(n_1048),
.B1(n_1049),
.B2(n_1047),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1084),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1078),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1086),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1087),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1081),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1089),
.B(n_1038),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1088),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1079),
.B(n_1068),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1090),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1074),
.A2(n_1056),
.B1(n_1053),
.B2(n_1062),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1070),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1072),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1073),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1094),
.A2(n_1092),
.B1(n_1093),
.B2(n_1091),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1101),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1097),
.A2(n_1065),
.B(n_1061),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1095),
.A2(n_1069),
.B1(n_1089),
.B2(n_1080),
.C(n_1083),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1094),
.A2(n_1051),
.B1(n_1056),
.B2(n_1081),
.Y(n_1115)
);

AOI31xp33_ASAP7_75t_L g1116 ( 
.A1(n_1095),
.A2(n_1065),
.A3(n_1076),
.B(n_1069),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1102),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_SL g1118 ( 
.A(n_1105),
.B(n_1075),
.Y(n_1118)
);

OAI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1107),
.A2(n_1052),
.B(n_1063),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_1104),
.A2(n_1063),
.B(n_1050),
.Y(n_1120)
);

OAI31xp33_ASAP7_75t_L g1121 ( 
.A1(n_1108),
.A2(n_1051),
.A3(n_1062),
.B(n_1053),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1109),
.A2(n_1051),
.B1(n_1062),
.B2(n_1047),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1099),
.B(n_1061),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1103),
.B(n_1048),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_1106),
.A2(n_1049),
.B(n_1026),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1096),
.B(n_1066),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1098),
.A2(n_1077),
.B(n_1012),
.C(n_1017),
.Y(n_1127)
);

AOI222xp33_ASAP7_75t_L g1128 ( 
.A1(n_1111),
.A2(n_1110),
.B1(n_1100),
.B2(n_1012),
.C1(n_1027),
.C2(n_1085),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_SL g1129 ( 
.A(n_1113),
.B(n_936),
.C(n_1060),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1123),
.Y(n_1130)
);

NOR4xp25_ASAP7_75t_L g1131 ( 
.A(n_1115),
.B(n_981),
.C(n_984),
.D(n_976),
.Y(n_1131)
);

OAI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1121),
.A2(n_1011),
.B1(n_857),
.B2(n_1014),
.C(n_1031),
.Y(n_1132)
);

OAI211xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1114),
.A2(n_984),
.B(n_903),
.C(n_910),
.Y(n_1133)
);

AOI211xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1116),
.A2(n_1011),
.B(n_984),
.C(n_903),
.Y(n_1134)
);

OAI211xp5_ASAP7_75t_L g1135 ( 
.A1(n_1112),
.A2(n_1114),
.B(n_1119),
.C(n_1122),
.Y(n_1135)
);

NAND4xp25_ASAP7_75t_L g1136 ( 
.A(n_1126),
.B(n_910),
.C(n_973),
.D(n_974),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1112),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1125),
.B(n_1124),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1118),
.A2(n_1031),
.B1(n_1018),
.B2(n_1014),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1127),
.B(n_191),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1120),
.B(n_949),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1117),
.B(n_907),
.C(n_974),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1114),
.B(n_1005),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_L g1144 ( 
.A(n_1130),
.B(n_1005),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1135),
.B(n_193),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1137),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1143),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1131),
.A2(n_1018),
.B1(n_1006),
.B2(n_995),
.C(n_993),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1141),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1140),
.A2(n_907),
.B1(n_920),
.B2(n_1006),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1134),
.A2(n_888),
.B(n_907),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1138),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1128),
.A2(n_888),
.B(n_875),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1139),
.B(n_949),
.Y(n_1154)
);

OA22x2_ASAP7_75t_L g1155 ( 
.A1(n_1152),
.A2(n_1129),
.B1(n_1128),
.B2(n_1133),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1146),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_L g1157 ( 
.A(n_1149),
.B(n_1147),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1145),
.B(n_1132),
.C(n_1136),
.Y(n_1158)
);

AOI211xp5_ASAP7_75t_L g1159 ( 
.A1(n_1153),
.A2(n_1142),
.B(n_909),
.C(n_875),
.Y(n_1159)
);

AO22x2_ASAP7_75t_L g1160 ( 
.A1(n_1154),
.A2(n_995),
.B1(n_822),
.B2(n_897),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1150),
.B(n_885),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1156),
.B(n_1148),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1161),
.B(n_1144),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_L g1164 ( 
.A(n_1157),
.B(n_1153),
.C(n_1151),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1158),
.B(n_889),
.C(n_909),
.Y(n_1165)
);

NOR3x1_ASAP7_75t_L g1166 ( 
.A(n_1155),
.B(n_889),
.C(n_897),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1159),
.B(n_194),
.Y(n_1167)
);

NAND4xp75_ASAP7_75t_L g1168 ( 
.A(n_1160),
.B(n_197),
.C(n_198),
.D(n_200),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1168),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_1164),
.B(n_203),
.Y(n_1170)
);

NAND4xp75_ASAP7_75t_L g1171 ( 
.A(n_1166),
.B(n_207),
.C(n_211),
.D(n_212),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1162),
.Y(n_1172)
);

NAND4xp75_ASAP7_75t_L g1173 ( 
.A(n_1167),
.B(n_213),
.C(n_214),
.D(n_215),
.Y(n_1173)
);

NAND4xp75_ASAP7_75t_L g1174 ( 
.A(n_1163),
.B(n_216),
.C(n_218),
.D(n_219),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1172),
.B(n_1165),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1169),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1171),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1170),
.B(n_221),
.C(n_225),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_SL g1179 ( 
.A(n_1174),
.B(n_1173),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1176),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1175),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1177),
.A2(n_893),
.B1(n_227),
.B2(n_231),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1179),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1180),
.A2(n_1178),
.B1(n_234),
.B2(n_239),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1183),
.A2(n_226),
.B1(n_240),
.B2(n_244),
.Y(n_1185)
);

AOI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1181),
.A2(n_245),
.B(n_246),
.Y(n_1186)
);

AO22x2_ASAP7_75t_SL g1187 ( 
.A1(n_1182),
.A2(n_250),
.B1(n_253),
.B2(n_256),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1184),
.A2(n_260),
.B1(n_262),
.B2(n_265),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1187),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1185),
.A2(n_266),
.B(n_267),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1189),
.A2(n_1186),
.B(n_271),
.Y(n_1191)
);

OAI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1188),
.A2(n_268),
.B(n_272),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1190),
.A2(n_275),
.B1(n_278),
.B2(n_283),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1191),
.B(n_292),
.Y(n_1194)
);

AO221x2_ASAP7_75t_L g1195 ( 
.A1(n_1192),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.C(n_297),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_313),
.B1(n_304),
.B2(n_305),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1194),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1197),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1198),
.A2(n_1195),
.B1(n_1196),
.B2(n_298),
.Y(n_1199)
);


endmodule