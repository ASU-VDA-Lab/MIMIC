module real_aes_2464_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_13;
wire n_7;
wire n_8;
wire n_12;
wire n_9;
wire n_14;
wire n_10;
wire n_11;
AOI221xp5_ASAP7_75t_L g6 ( .A1(n_0), .A2(n_2), .B1(n_7), .B2(n_12), .C(n_13), .Y(n_6) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_14), .Y(n_13) );
BUFx2_ASAP7_75t_SL g9 ( .A(n_4), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
INVx1_ASAP7_75t_SL g12 ( .A(n_7), .Y(n_12) );
NOR2xp33_ASAP7_75t_SL g7 ( .A(n_8), .B(n_10), .Y(n_7) );
CKINVDCx8_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
endmodule