module real_jpeg_24683_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

AO21x1_ASAP7_75t_SL g11 ( 
.A1(n_2),
.A2(n_12),
.B(n_14),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_19),
.B(n_21),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.C(n_33),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_16),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_12),
.A2(n_14),
.B(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_15),
.A2(n_38),
.B(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_21),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);


endmodule