module fake_jpeg_175_n_114 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_16),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_30),
.B1(n_35),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_72),
.B1(n_53),
.B2(n_44),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_40),
.C(n_31),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_14),
.A3(n_26),
.B1(n_15),
.B2(n_34),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_73),
.B(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_22),
.B2(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_10),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_89),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_71),
.B(n_67),
.C(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_65),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_67),
.C(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_78),
.B1(n_76),
.B2(n_82),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_53),
.A3(n_52),
.B1(n_13),
.B2(n_3),
.C1(n_9),
.C2(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_13),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_78),
.B1(n_58),
.B2(n_79),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_48),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_100),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_96),
.C(n_95),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_91),
.C(n_97),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_78),
.A3(n_64),
.B1(n_61),
.B2(n_75),
.C1(n_18),
.C2(n_50),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_60),
.C(n_56),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_102),
.B(n_50),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_103),
.B(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_102),
.B1(n_97),
.B2(n_92),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);

NAND4xp25_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_0),
.C(n_2),
.D(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_105),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_0),
.B(n_2),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_2),
.C(n_41),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_42),
.Y(n_114)
);


endmodule