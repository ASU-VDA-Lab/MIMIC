module fake_jpeg_9279_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_32),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_61),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_33),
.B1(n_34),
.B2(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_60),
.B1(n_34),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_27),
.B1(n_17),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_62),
.B1(n_65),
.B2(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_33),
.B1(n_24),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_22),
.B1(n_18),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_34),
.B1(n_23),
.B2(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_74),
.Y(n_105)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_88),
.B1(n_53),
.B2(n_49),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_34),
.B1(n_20),
.B2(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_72),
.B1(n_61),
.B2(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_0),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_59),
.C(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_20),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_2),
.Y(n_108)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_111),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_44),
.A3(n_56),
.B1(n_49),
.B2(n_53),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_71),
.B(n_69),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_119),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_89),
.B1(n_62),
.B2(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_4),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_4),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_66),
.B1(n_81),
.B2(n_80),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_141),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_110),
.B1(n_96),
.B2(n_118),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_83),
.B1(n_70),
.B2(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_128),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_122),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_67),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_107),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_133),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_86),
.C(n_93),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_139),
.C(n_100),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_68),
.B1(n_66),
.B2(n_76),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_146),
.B1(n_114),
.B2(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_111),
.C(n_97),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_97),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_103),
.B1(n_119),
.B2(n_95),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_66),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_108),
.B(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_90),
.B1(n_82),
.B2(n_74),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_171),
.B1(n_154),
.B2(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_148),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_107),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_157),
.C(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_162),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_158),
.B(n_173),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_103),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_117),
.B(n_116),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_123),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_134),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_104),
.B1(n_117),
.B2(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_125),
.B1(n_126),
.B2(n_121),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_153),
.B1(n_156),
.B2(n_160),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_160),
.B(n_7),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_127),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_138),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_132),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_5),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_152),
.B(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_145),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_174),
.B1(n_173),
.B2(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_162),
.C(n_148),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_104),
.C(n_7),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_171),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_168),
.B1(n_149),
.B2(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_215),
.B1(n_177),
.B2(n_191),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_219),
.B(n_192),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_216),
.C(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_104),
.B1(n_73),
.B2(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_198),
.B(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.C(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_201),
.B1(n_202),
.B2(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_188),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_228),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_184),
.Y(n_225)
);

BUFx12f_ASAP7_75t_SL g227 ( 
.A(n_211),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_229),
.B(n_219),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_183),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_189),
.Y(n_229)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_207),
.B(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_186),
.C(n_176),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_212),
.C(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_221),
.B(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_244),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_208),
.B(n_204),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_232),
.B(n_231),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_185),
.B1(n_197),
.B2(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_214),
.B1(n_215),
.B2(n_189),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_223),
.B(n_8),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_225),
.C(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_226),
.B(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_252),
.B(n_239),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_234),
.B(n_230),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_240),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_223),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_5),
.C(n_8),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_5),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_257),
.B1(n_252),
.B2(n_256),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_246),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_247),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_271),
.A3(n_259),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_9),
.Y(n_271)
);

AOI321xp33_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_259),
.A3(n_260),
.B1(n_12),
.B2(n_13),
.C(n_10),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.C(n_269),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.C(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_268),
.C(n_11),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_10),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_11),
.Y(n_280)
);


endmodule