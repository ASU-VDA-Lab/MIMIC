module fake_jpeg_2865_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g14 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx12_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_6),
.B1(n_11),
.B2(n_9),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_29),
.B1(n_20),
.B2(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_13),
.B(n_9),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_21),
.C(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_13),
.B1(n_16),
.B2(n_12),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_32),
.B(n_22),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_25),
.C(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_36),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_3),
.B(n_4),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_32),
.CI(n_33),
.CON(n_38),
.SN(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_3),
.B(n_5),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_38),
.C(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_40),
.B(n_38),
.Y(n_44)
);


endmodule