module fake_jpeg_31979_n_512 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_512);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_512;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_53),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_97),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_61),
.A2(n_45),
.B1(n_50),
.B2(n_31),
.Y(n_156)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_63),
.Y(n_146)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_19),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_21),
.B1(n_24),
.B2(n_34),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_2),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_96),
.Y(n_119)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_19),
.B(n_3),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_100),
.Y(n_126)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_3),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_21),
.B1(n_39),
.B2(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_108),
.A2(n_131),
.B1(n_136),
.B2(n_147),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_48),
.B(n_51),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g181 ( 
.A(n_112),
.B(n_73),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_123),
.B(n_133),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_139),
.B1(n_45),
.B2(n_27),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_67),
.B1(n_101),
.B2(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_62),
.B(n_38),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_32),
.B1(n_21),
.B2(n_26),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_52),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_142),
.B(n_148),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_89),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_70),
.A2(n_26),
.B1(n_40),
.B2(n_18),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_52),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_55),
.B(n_51),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_93),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_82),
.A2(n_26),
.B1(n_40),
.B2(n_50),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_23),
.B1(n_100),
.B2(n_96),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_27),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_165),
.B(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_167),
.B(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_141),
.Y(n_171)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_75),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_178),
.Y(n_233)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_175),
.A2(n_211),
.B1(n_108),
.B2(n_109),
.Y(n_227)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_176),
.Y(n_258)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_103),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_182),
.B(n_188),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_118),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_156),
.B(n_119),
.C(n_153),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_150),
.B1(n_146),
.B2(n_109),
.Y(n_240)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_56),
.B1(n_86),
.B2(n_23),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_30),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_31),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

BUFx16f_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_210),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_110),
.B(n_30),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_214),
.Y(n_249)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

AO22x1_ASAP7_75t_SL g215 ( 
.A1(n_136),
.A2(n_94),
.B1(n_71),
.B2(n_90),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_215),
.B(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_87),
.C(n_84),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_160),
.C(n_162),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_163),
.B1(n_122),
.B2(n_151),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_221),
.A2(n_240),
.B1(n_243),
.B2(n_250),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_225),
.B(n_191),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_227),
.A2(n_235),
.B1(n_256),
.B2(n_259),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_181),
.A2(n_131),
.B1(n_147),
.B2(n_151),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_184),
.A2(n_163),
.B1(n_150),
.B2(n_155),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_188),
.A2(n_114),
.B1(n_121),
.B2(n_115),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_189),
.B(n_146),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_193),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_121),
.C(n_115),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_217),
.C(n_167),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_182),
.A2(n_114),
.B1(n_130),
.B2(n_18),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_188),
.A2(n_93),
.B1(n_58),
.B2(n_18),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_167),
.A2(n_58),
.B1(n_130),
.B2(n_6),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_215),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_266),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_175),
.B(n_203),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_263),
.A2(n_270),
.B(n_279),
.Y(n_330)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_195),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_295),
.Y(n_325)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_212),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_276),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_203),
.B(n_183),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_271),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_261),
.B(n_253),
.C(n_259),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_242),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_273),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_274),
.A2(n_296),
.B1(n_267),
.B2(n_273),
.Y(n_313)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_192),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_171),
.B(n_198),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_187),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_281),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_185),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_284),
.A2(n_287),
.B1(n_290),
.B2(n_298),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_211),
.B(n_205),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_292),
.B(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_260),
.B(n_166),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_215),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_297),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_228),
.A2(n_190),
.B(n_179),
.C(n_194),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_169),
.C(n_210),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_228),
.C(n_247),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_224),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_238),
.B(n_255),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_214),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_253),
.B(n_240),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_296),
.Y(n_335)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_235),
.A3(n_227),
.B1(n_233),
.B2(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_320),
.B(n_326),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_313),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_236),
.B1(n_223),
.B2(n_226),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_314),
.A2(n_316),
.B1(n_333),
.B2(n_298),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_236),
.B1(n_223),
.B2(n_226),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_247),
.C(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_322),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_263),
.A2(n_222),
.B(n_241),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_266),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_220),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_220),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_329),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_220),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_279),
.A2(n_229),
.B(n_251),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_331),
.A2(n_292),
.B(n_289),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_272),
.A2(n_257),
.B1(n_201),
.B2(n_238),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_335),
.B(n_344),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_272),
.B1(n_280),
.B2(n_276),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_336),
.A2(n_342),
.B1(n_319),
.B2(n_306),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_271),
.B1(n_283),
.B2(n_265),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_343),
.B1(n_353),
.B2(n_355),
.Y(n_377)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

BUFx8_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_340),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_R g341 ( 
.A1(n_318),
.A2(n_285),
.B(n_281),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_299),
.B1(n_304),
.B2(n_311),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_302),
.B1(n_324),
.B2(n_312),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_307),
.A2(n_270),
.B(n_282),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_301),
.A2(n_277),
.B1(n_285),
.B2(n_289),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_331),
.B(n_332),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g395 ( 
.A1(n_345),
.A2(n_351),
.B(n_194),
.C(n_239),
.D(n_6),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_332),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_356),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_348),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_262),
.Y(n_349)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_330),
.A2(n_297),
.B(n_269),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_324),
.A2(n_289),
.B1(n_290),
.B2(n_284),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_326),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_287),
.B1(n_292),
.B2(n_294),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_364),
.B1(n_365),
.B2(n_288),
.Y(n_384)
);

OA22x2_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_275),
.B1(n_238),
.B2(n_251),
.Y(n_362)
);

AOI22x1_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_323),
.B1(n_320),
.B2(n_264),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_306),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_316),
.A2(n_275),
.B1(n_258),
.B2(n_176),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_258),
.B1(n_288),
.B2(n_257),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_325),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_389),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_369),
.A2(n_380),
.B1(n_337),
.B2(n_365),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_350),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_370),
.B(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

AOI22x1_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_325),
.B1(n_312),
.B2(n_311),
.Y(n_376)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_329),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_379),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_328),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_338),
.A2(n_309),
.B1(n_299),
.B2(n_315),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_322),
.C(n_229),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_348),
.C(n_355),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_346),
.B(n_315),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_384),
.A2(n_393),
.B1(n_362),
.B2(n_339),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_173),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_268),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_394),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_244),
.Y(n_391)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_356),
.A2(n_244),
.B1(n_239),
.B2(n_200),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_345),
.B(n_357),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_396),
.A2(n_17),
.B(n_5),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_363),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_399),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_400),
.A2(n_419),
.B1(n_398),
.B2(n_393),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_402),
.C(n_403),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_359),
.C(n_344),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_381),
.C(n_390),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_413),
.B1(n_415),
.B2(n_417),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_406),
.A2(n_408),
.B1(n_375),
.B2(n_380),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_335),
.C(n_344),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_394),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_384),
.A2(n_335),
.B1(n_344),
.B2(n_357),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_344),
.C(n_353),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_377),
.C(n_376),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_366),
.B(n_346),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_382),
.A2(n_358),
.B(n_360),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_416),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_391),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_362),
.B(n_364),
.C(n_340),
.Y(n_418)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_369),
.A2(n_362),
.B1(n_340),
.B2(n_6),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_428),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_425),
.A2(n_407),
.B1(n_405),
.B2(n_8),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_414),
.A2(n_377),
.B1(n_385),
.B2(n_388),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_434),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_389),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_432),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_395),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_406),
.B1(n_408),
.B2(n_412),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_402),
.B(n_375),
.CI(n_387),
.CON(n_434),
.SN(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_373),
.C(n_392),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_438),
.C(n_441),
.Y(n_449)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_437),
.Y(n_444)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_340),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_439),
.A2(n_418),
.B(n_414),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_440),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_16),
.Y(n_441)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g446 ( 
.A1(n_434),
.A2(n_400),
.B(n_396),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_451),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_423),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_454),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_450),
.B1(n_440),
.B2(n_437),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_409),
.B1(n_419),
.B2(n_404),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g452 ( 
.A(n_442),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_452),
.B(n_432),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_411),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_425),
.A2(n_429),
.B1(n_428),
.B2(n_409),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_424),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_401),
.C(n_410),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_438),
.C(n_431),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_405),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_457),
.B(n_458),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_424),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_468),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_456),
.A2(n_427),
.B(n_426),
.Y(n_461)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_465),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_470),
.C(n_471),
.Y(n_480)
);

INVx6_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_449),
.C(n_458),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_422),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_444),
.A2(n_439),
.B(n_433),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_472),
.A2(n_460),
.B(n_469),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_441),
.C(n_436),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_4),
.C(n_7),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_475),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_464),
.B(n_453),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_483),
.Y(n_496)
);

OAI211xp5_ASAP7_75t_L g477 ( 
.A1(n_462),
.A2(n_450),
.B(n_448),
.C(n_459),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_479),
.B(n_485),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_478),
.A2(n_482),
.B(n_12),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_472),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_4),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_470),
.A2(n_8),
.B(n_9),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_474),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_490),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_467),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_484),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_494),
.Y(n_503)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_486),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_12),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_495),
.B(n_497),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_478),
.A2(n_12),
.B(n_13),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_487),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_498),
.A2(n_479),
.B(n_15),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_487),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_502),
.A2(n_477),
.B(n_496),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_506),
.B(n_500),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_500),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_14),
.B(n_16),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_507),
.A2(n_508),
.B(n_501),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_503),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_14),
.C(n_16),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_511),
.Y(n_512)
);


endmodule