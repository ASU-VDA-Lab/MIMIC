module fake_netlist_6_1430_n_185 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_185);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_185;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_130;
wire n_84;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx4_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_16),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_1),
.C(n_4),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_5),
.Y(n_73)
);

AND3x2_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_5),
.C(n_7),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_42),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_45),
.B1(n_51),
.B2(n_42),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_62),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_54),
.B1(n_36),
.B2(n_40),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_41),
.B(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22x1_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_61),
.B1(n_63),
.B2(n_71),
.Y(n_95)
);

AO31x2_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_72),
.A3(n_69),
.B(n_68),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_65),
.B(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_74),
.B(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_72),
.B(n_69),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2x1_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_91),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_91),
.B(n_89),
.C(n_83),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_87),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_85),
.B(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_67),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_79),
.B1(n_64),
.B2(n_46),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_95),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_101),
.B(n_85),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_108),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_112),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_114),
.B1(n_90),
.B2(n_115),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_95),
.B(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_116),
.B(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_111),
.B1(n_61),
.B2(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_134),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_129),
.Y(n_143)
);

NAND4xp25_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_126),
.C(n_129),
.D(n_56),
.Y(n_144)
);

AOI321xp33_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_45),
.A3(n_133),
.B1(n_59),
.B2(n_60),
.C(n_68),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_74),
.C(n_75),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_33),
.B1(n_132),
.B2(n_75),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_60),
.C(n_59),
.Y(n_148)
);

O2A1O1Ixp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_130),
.B(n_62),
.C(n_69),
.Y(n_149)
);

OAI221xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_57),
.B1(n_75),
.B2(n_88),
.C(n_72),
.Y(n_150)
);

NAND2x1p5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_57),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_57),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_7),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_144),
.B1(n_145),
.B2(n_88),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_93),
.B(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_8),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_8),
.C(n_9),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_102),
.B(n_78),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_161),
.B1(n_156),
.B2(n_93),
.C(n_13),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_86),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_41),
.A3(n_86),
.B1(n_84),
.B2(n_78),
.C1(n_22),
.C2(n_28),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_84),
.A3(n_86),
.B1(n_19),
.B2(n_20),
.C1(n_14),
.C2(n_15),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_84),
.C(n_96),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

NOR4xp75_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_164),
.C(n_163),
.D(n_168),
.Y(n_177)
);

NAND4xp25_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_162),
.C(n_170),
.D(n_96),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_96),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_172),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_103),
.B1(n_178),
.B2(n_171),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_103),
.B(n_182),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_181),
.B1(n_183),
.B2(n_180),
.C(n_103),
.Y(n_185)
);


endmodule