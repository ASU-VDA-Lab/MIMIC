module fake_ibex_1239_n_1071 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1071);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1071;

wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1031;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_736;
wire n_550;
wire n_1055;
wire n_732;
wire n_673;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_496;
wire n_301;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_646;
wire n_448;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_580;
wire n_483;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_849;
wire n_765;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_648;
wire n_571;
wire n_472;
wire n_209;
wire n_229;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_947;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_195;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_912;
wire n_874;
wire n_890;
wire n_921;
wire n_1058;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_90),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_23),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_47),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g201 ( 
.A(n_97),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_86),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_29),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_98),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_0),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_78),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_100),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_99),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_13),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_159),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_65),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_131),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_150),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_5),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_92),
.B(n_180),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_29),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_121),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_55),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_25),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_81),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_157),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_88),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_144),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_132),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_26),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_72),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_79),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_58),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_87),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_40),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_37),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_46),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_42),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_89),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_50),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_147),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_154),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_152),
.B(n_165),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_25),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_42),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_26),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_117),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_11),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_155),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_83),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_127),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_146),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_136),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_137),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_69),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_124),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_10),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_20),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_169),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_46),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_108),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_64),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_33),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_52),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_9),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_35),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_179),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_59),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_118),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_8),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_107),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_114),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_156),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_19),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_143),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_142),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_22),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_76),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_148),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_182),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_50),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_15),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_103),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_133),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_19),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_106),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_171),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_158),
.B(n_140),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_134),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_16),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_123),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_70),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_96),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_61),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_232),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_232),
.B(n_2),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_258),
.B(n_211),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_199),
.B(n_191),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_221),
.B(n_3),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_200),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_221),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_208),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_242),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_224),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_187),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_242),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_187),
.A2(n_74),
.B(n_176),
.Y(n_348)
);

CKINVDCx8_ASAP7_75t_R g349 ( 
.A(n_185),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_199),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_192),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_209),
.B(n_288),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_200),
.B(n_6),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_233),
.B(n_6),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g357 ( 
.A1(n_192),
.A2(n_75),
.B(n_175),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_186),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_204),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_188),
.B(n_53),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_8),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_204),
.A2(n_80),
.B(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_236),
.B(n_235),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_259),
.B(n_9),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_186),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_214),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_280),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_183),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_207),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_242),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_209),
.B(n_14),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_242),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_190),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_207),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_274),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_193),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_208),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_243),
.B(n_17),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_261),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_311),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_253),
.B(n_18),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_214),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_274),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_250),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_189),
.B(n_21),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_288),
.B(n_24),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_203),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_261),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_219),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_262),
.B(n_27),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_325),
.B(n_30),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_262),
.B(n_30),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_239),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_230),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_241),
.Y(n_398)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_250),
.Y(n_399)
);

CKINVDCx8_ASAP7_75t_R g400 ( 
.A(n_201),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_247),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_251),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_269),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_251),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_325),
.B(n_255),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_249),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_230),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_252),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_255),
.B(n_31),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_276),
.B(n_34),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_274),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_269),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_276),
.A2(n_122),
.B(n_173),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_292),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_271),
.B(n_34),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_230),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_263),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_244),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_265),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_292),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_271),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_244),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_327),
.B(n_38),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_275),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_39),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_277),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_272),
.B(n_41),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_282),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_244),
.B(n_129),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_272),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_273),
.B(n_43),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_290),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_273),
.B(n_43),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_287),
.B(n_44),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_287),
.B(n_45),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_293),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_291),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_194),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_195),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_299),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_244),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_358),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_339),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_378),
.B(n_304),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_353),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_374),
.B(n_197),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_352),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_374),
.B(n_389),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_198),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_337),
.B(n_293),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_386),
.B(n_205),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_343),
.B(n_309),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_352),
.Y(n_468)
);

INVx4_ASAP7_75t_SL g469 ( 
.A(n_352),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_386),
.B(n_206),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_349),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_358),
.B(n_294),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_399),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_400),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_372),
.A2(n_312),
.B1(n_284),
.B2(n_227),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_362),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_362),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_350),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_382),
.B(n_184),
.Y(n_484)
);

NOR2x1p5_ASAP7_75t_L g485 ( 
.A(n_336),
.B(n_308),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_409),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_382),
.B(n_184),
.Y(n_489)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_342),
.B(n_316),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_380),
.B(n_317),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_410),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_412),
.B(n_196),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_341),
.B(n_305),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_345),
.B(n_210),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_389),
.B(n_394),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_394),
.B(n_212),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_305),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_368),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_381),
.B(n_248),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_403),
.B(n_196),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_349),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_425),
.B(n_213),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_425),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_365),
.B(n_217),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_405),
.B(n_215),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_381),
.B(n_248),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

INVx4_ASAP7_75t_SL g519 ( 
.A(n_338),
.Y(n_519)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_361),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_334),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_371),
.A2(n_324),
.B1(n_332),
.B2(n_330),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_424),
.B(n_220),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_357),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_334),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_393),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_424),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_424),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_376),
.B(n_215),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_427),
.B(n_223),
.Y(n_531)
);

AND3x2_ASAP7_75t_L g532 ( 
.A(n_356),
.B(n_216),
.C(n_264),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_379),
.B(n_218),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_357),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_395),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_427),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_356),
.B(n_366),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_390),
.A2(n_333),
.B1(n_323),
.B2(n_320),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_440),
.B(n_441),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_366),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_415),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_392),
.B(n_218),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

BUFx8_ASAP7_75t_SL g547 ( 
.A(n_432),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_434),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_435),
.B(n_436),
.C(n_384),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_396),
.B(n_225),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_222),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_346),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_348),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_348),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_361),
.A2(n_370),
.B1(n_383),
.B2(n_421),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_357),
.B(n_237),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_440),
.B(n_238),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_441),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_406),
.B(n_240),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_443),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_391),
.A2(n_286),
.B1(n_257),
.B2(n_314),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_351),
.B(n_245),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_408),
.B(n_248),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_359),
.B(n_246),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_417),
.B(n_254),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_556),
.A2(n_266),
.B1(n_285),
.B2(n_284),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_547),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_450),
.B(n_256),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_479),
.B(n_335),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_490),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_485),
.A2(n_266),
.B1(n_285),
.B2(n_227),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_493),
.A2(n_369),
.B1(n_385),
.B2(n_439),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_527),
.B(n_536),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_490),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_419),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_429),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_493),
.A2(n_387),
.B1(n_385),
.B2(n_439),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_530),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_530),
.Y(n_583)
);

BUFx5_ASAP7_75t_L g584 ( 
.A(n_452),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_560),
.B(n_433),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_518),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_514),
.A2(n_438),
.B1(n_442),
.B2(n_437),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_554),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_444),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_547),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_566),
.B(n_388),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_566),
.B(n_222),
.Y(n_592)
);

NAND2x1_ASAP7_75t_L g593 ( 
.A(n_477),
.B(n_363),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_534),
.B(n_226),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_473),
.B(n_354),
.Y(n_597)
);

A2O1A1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_446),
.A2(n_413),
.B(n_426),
.C(n_420),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_444),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_528),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

AO21x1_ASAP7_75t_L g603 ( 
.A1(n_525),
.A2(n_413),
.B(n_335),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_537),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_551),
.B(n_228),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_479),
.B(n_488),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_545),
.B(n_229),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_544),
.A2(n_401),
.B1(n_315),
.B2(n_329),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_364),
.Y(n_610)
);

AND2x6_ASAP7_75t_SL g611 ( 
.A(n_466),
.B(n_247),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_516),
.B(n_231),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_559),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_505),
.B(n_506),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_543),
.B(n_340),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_453),
.B(n_267),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_451),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_461),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_500),
.B(n_260),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_549),
.B(n_340),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_493),
.A2(n_387),
.B1(n_426),
.B2(n_420),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_283),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_447),
.A2(n_359),
.B1(n_414),
.B2(n_404),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_451),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_522),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_538),
.A2(n_369),
.B1(n_414),
.B2(n_404),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_546),
.B(n_283),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_526),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_451),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_542),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

NOR2x1p5_ASAP7_75t_L g635 ( 
.A(n_510),
.B(n_289),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_510),
.B(n_315),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

OR2x6_ASAP7_75t_SL g638 ( 
.A(n_478),
.B(n_268),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_464),
.A2(n_270),
.B1(n_402),
.B2(n_278),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_449),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_492),
.B(n_340),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_562),
.A2(n_360),
.B1(n_355),
.B2(n_367),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_520),
.B(n_504),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_492),
.B(n_355),
.Y(n_644)
);

OAI22xp33_ASAP7_75t_L g645 ( 
.A1(n_466),
.A2(n_355),
.B1(n_360),
.B2(n_367),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_508),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_457),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_467),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_484),
.B(n_360),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_489),
.B(n_367),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_496),
.B(n_281),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_468),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_468),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_511),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_469),
.B(n_279),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_469),
.B(n_296),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_462),
.A2(n_313),
.B1(n_310),
.B2(n_301),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_466),
.A2(n_307),
.B1(n_306),
.B2(n_302),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_463),
.B(n_295),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_511),
.B(n_303),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_557),
.B(n_326),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_504),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_480),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_598),
.A2(n_535),
.B(n_525),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_575),
.B(n_474),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_623),
.A2(n_502),
.B(n_524),
.C(n_531),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_593),
.A2(n_554),
.B(n_555),
.Y(n_670)
);

AO32x1_ASAP7_75t_L g671 ( 
.A1(n_629),
.A2(n_525),
.A3(n_535),
.B1(n_499),
.B2(n_498),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_633),
.B(n_578),
.Y(n_672)
);

BUFx6f_ASAP7_75t_SL g673 ( 
.A(n_664),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_600),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_588),
.A2(n_363),
.B(n_486),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_598),
.A2(n_555),
.B(n_535),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_582),
.A2(n_481),
.B(n_482),
.C(n_495),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_645),
.A2(n_562),
.B1(n_501),
.B2(n_550),
.C(n_487),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_614),
.B(n_520),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_617),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_663),
.A2(n_460),
.B(n_503),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_643),
.A2(n_521),
.B1(n_476),
.B2(n_562),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_620),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_582),
.A2(n_512),
.B(n_460),
.C(n_503),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_568),
.B(n_465),
.C(n_471),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_637),
.B(n_476),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_627),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_590),
.B(n_521),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_583),
.B(n_521),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_583),
.B(n_532),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_611),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_623),
.A2(n_512),
.B(n_491),
.C(n_509),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_607),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_580),
.B(n_540),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_648),
.B(n_454),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_585),
.B(n_491),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_642),
.B(n_507),
.C(n_517),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_620),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_632),
.B(n_491),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_587),
.A2(n_517),
.B(n_507),
.C(n_565),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_567),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_645),
.A2(n_565),
.B(n_466),
.C(n_494),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_591),
.A2(n_491),
.B1(n_509),
.B2(n_523),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_651),
.A2(n_494),
.B(n_430),
.C(n_564),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_646),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_647),
.Y(n_711)
);

CKINVDCx11_ASAP7_75t_R g712 ( 
.A(n_638),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_656),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_642),
.A2(n_491),
.B1(n_509),
.B2(n_494),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_630),
.B(n_509),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_640),
.A2(n_553),
.B1(n_561),
.B2(n_234),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_637),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_613),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_592),
.B(n_454),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_618),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_634),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_597),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_596),
.B(n_483),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_573),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_649),
.A2(n_561),
.B(n_553),
.C(n_430),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_606),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_652),
.A2(n_445),
.B(n_448),
.C(n_455),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_615),
.B(n_558),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_621),
.B(n_558),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_558),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_650),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_653),
.B(n_625),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_610),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_609),
.B(n_558),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_628),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_665),
.A2(n_298),
.B(n_319),
.C(n_338),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_639),
.B(n_563),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_660),
.A2(n_563),
.B1(n_319),
.B2(n_418),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_612),
.B(n_563),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_661),
.A2(n_456),
.B(n_458),
.C(n_459),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_571),
.B(n_563),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_601),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_588),
.A2(n_603),
.B(n_570),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_569),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_635),
.B(n_319),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_636),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_602),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_572),
.B(n_563),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_579),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_576),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_577),
.B(n_49),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_659),
.A2(n_574),
.B(n_581),
.C(n_624),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_672),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_694),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_733),
.A2(n_624),
.B(n_581),
.C(n_574),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_736),
.Y(n_761)
);

NAND2x1p5_ASAP7_75t_L g762 ( 
.A(n_696),
.B(n_586),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_704),
.A2(n_599),
.B1(n_662),
.B2(n_622),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_705),
.A2(n_626),
.B(n_616),
.C(n_657),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_743),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_674),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_670),
.A2(n_677),
.B(n_666),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_748),
.Y(n_768)
);

AO32x2_ASAP7_75t_L g769 ( 
.A1(n_716),
.A2(n_626),
.A3(n_422),
.B1(n_347),
.B2(n_373),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_755),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_680),
.B(n_657),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_732),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_756),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_717),
.B(n_595),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_683),
.A2(n_595),
.B1(n_619),
.B2(n_658),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_655),
.B(n_654),
.C(n_619),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_675),
.B(n_619),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_701),
.B(n_54),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_727),
.A2(n_458),
.B(n_470),
.C(n_456),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_721),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_750),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_679),
.B(n_695),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_679),
.A2(n_422),
.B1(n_344),
.B2(n_347),
.C(n_373),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_584),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_724),
.B(n_584),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_726),
.A2(n_533),
.A3(n_513),
.B(n_459),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_690),
.B(n_584),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_703),
.A2(n_422),
.B(n_338),
.C(n_375),
.Y(n_789)
);

OAI22x1_ASAP7_75t_L g790 ( 
.A1(n_692),
.A2(n_57),
.B1(n_63),
.B2(n_66),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_691),
.B(n_584),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_708),
.B(n_375),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_734),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_709),
.B(n_678),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_687),
.B(n_373),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_752),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_669),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_682),
.A2(n_347),
.B(n_344),
.C(n_338),
.Y(n_798)
);

OAI21x1_ASAP7_75t_SL g799 ( 
.A1(n_678),
.A2(n_67),
.B(n_71),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_737),
.A2(n_347),
.A3(n_344),
.B(n_519),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_SL g801 ( 
.A1(n_693),
.A2(n_73),
.B(n_85),
.C(n_93),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_681),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_757),
.A2(n_344),
.B1(n_539),
.B2(n_101),
.Y(n_803)
);

OAI222xp33_ASAP7_75t_L g804 ( 
.A1(n_714),
.A2(n_94),
.B1(n_95),
.B2(n_104),
.C1(n_110),
.C2(n_113),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_730),
.A2(n_344),
.B(n_539),
.C(n_130),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_688),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_687),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_722),
.B(n_168),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_178),
.Y(n_809)
);

AO31x2_ASAP7_75t_L g810 ( 
.A1(n_671),
.A2(n_170),
.A3(n_172),
.B(n_706),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_747),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_740),
.A2(n_715),
.B(n_671),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_685),
.A2(n_731),
.B(n_707),
.C(n_700),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_673),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_698),
.B(n_719),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_685),
.A2(n_738),
.B(n_699),
.C(n_686),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_SL g817 ( 
.A(n_669),
.B(n_697),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_739),
.B(n_741),
.C(n_746),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_753),
.A2(n_707),
.B(n_702),
.C(n_735),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_669),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_729),
.B(n_751),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_742),
.A2(n_741),
.B(n_728),
.C(n_749),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_745),
.B(n_720),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_712),
.B(n_689),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_710),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_673),
.A2(n_711),
.B1(n_713),
.B2(n_718),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_754),
.A2(n_733),
.B(n_705),
.C(n_668),
.Y(n_827)
);

AO31x2_ASAP7_75t_L g828 ( 
.A1(n_677),
.A2(n_598),
.A3(n_603),
.B(n_744),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_670),
.A2(n_677),
.B(n_588),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_672),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_672),
.B(n_667),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_677),
.A2(n_744),
.B(n_666),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_672),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_694),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_670),
.A2(n_677),
.B(n_588),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_672),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_677),
.A2(n_598),
.A3(n_603),
.B(n_744),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_670),
.A2(n_677),
.B(n_676),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_733),
.A2(n_705),
.B(n_668),
.C(n_703),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_672),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_694),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_674),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_672),
.B(n_667),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_672),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_694),
.B(n_600),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_675),
.Y(n_846)
);

AOI222xp33_ASAP7_75t_L g847 ( 
.A1(n_712),
.A2(n_556),
.B1(n_679),
.B2(n_538),
.C1(n_589),
.C2(n_600),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_672),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_667),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_831),
.B(n_843),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_849),
.B(n_833),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_844),
.B(n_830),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_836),
.B(n_840),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_758),
.B(n_848),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_759),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_758),
.B(n_848),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_772),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_847),
.A2(n_783),
.B1(n_794),
.B2(n_786),
.Y(n_858)
);

OA21x2_ASAP7_75t_L g859 ( 
.A1(n_838),
.A2(n_832),
.B(n_767),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_775),
.A2(n_784),
.B1(n_761),
.B2(n_773),
.Y(n_860)
);

AO31x2_ASAP7_75t_L g861 ( 
.A1(n_789),
.A2(n_813),
.A3(n_777),
.B(n_827),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_846),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_841),
.Y(n_863)
);

AO21x2_ASAP7_75t_L g864 ( 
.A1(n_798),
.A2(n_822),
.B(n_803),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_765),
.Y(n_865)
);

AOI221xp5_ASAP7_75t_L g866 ( 
.A1(n_768),
.A2(n_770),
.B1(n_816),
.B2(n_806),
.C(n_802),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_819),
.A2(n_760),
.B(n_764),
.C(n_779),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_779),
.A2(n_763),
.B1(n_815),
.B2(n_824),
.Y(n_868)
);

AOI221xp5_ASAP7_75t_L g869 ( 
.A1(n_807),
.A2(n_793),
.B1(n_826),
.B2(n_845),
.C(n_791),
.Y(n_869)
);

CKINVDCx6p67_ASAP7_75t_R g870 ( 
.A(n_811),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_796),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_797),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_771),
.B(n_834),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_823),
.B(n_774),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_825),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_766),
.B(n_842),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_823),
.B(n_774),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_778),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_821),
.B(n_785),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_808),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_762),
.B(n_782),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_799),
.A2(n_818),
.B1(n_795),
.B2(n_790),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_788),
.A2(n_809),
.B1(n_776),
.B2(n_782),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_792),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_828),
.B(n_837),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_797),
.B(n_820),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_804),
.A2(n_805),
.B(n_801),
.C(n_780),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_814),
.A2(n_820),
.B1(n_817),
.B2(n_837),
.Y(n_889)
);

OA21x2_ASAP7_75t_L g890 ( 
.A1(n_769),
.A2(n_810),
.B(n_787),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_800),
.B(n_834),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_800),
.B(n_831),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_833),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_758),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_847),
.A2(n_679),
.B1(n_642),
.B2(n_783),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_831),
.B(n_843),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_847),
.A2(n_679),
.B1(n_642),
.B2(n_783),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_759),
.B(n_841),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_831),
.B(n_843),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_SL g900 ( 
.A1(n_845),
.A2(n_444),
.B1(n_600),
.B2(n_704),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_758),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_849),
.B(n_843),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_839),
.A2(n_848),
.B(n_758),
.C(n_827),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_839),
.A2(n_848),
.B(n_758),
.C(n_827),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_812),
.A2(n_835),
.B(n_829),
.Y(n_905)
);

OAI22xp33_ASAP7_75t_L g906 ( 
.A1(n_831),
.A2(n_567),
.B1(n_849),
.B2(n_843),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_831),
.B(n_843),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_833),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_759),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_SL g910 ( 
.A1(n_845),
.A2(n_444),
.B1(n_600),
.B2(n_704),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_847),
.A2(n_679),
.B1(n_642),
.B2(n_783),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_812),
.A2(n_835),
.B(n_829),
.Y(n_912)
);

OAI221xp5_ASAP7_75t_L g913 ( 
.A1(n_847),
.A2(n_831),
.B1(n_849),
.B2(n_843),
.C(n_683),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_812),
.A2(n_835),
.B(n_829),
.Y(n_914)
);

CKINVDCx11_ASAP7_75t_R g915 ( 
.A(n_766),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_833),
.B(n_844),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_902),
.B(n_894),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_894),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_902),
.B(n_901),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_901),
.B(n_850),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_857),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_896),
.B(n_899),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_903),
.B(n_904),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_859),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_892),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_907),
.B(n_916),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_903),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_851),
.B(n_854),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_904),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_856),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_905),
.A2(n_914),
.B(n_912),
.Y(n_931)
);

OAI221xp5_ASAP7_75t_L g932 ( 
.A1(n_913),
.A2(n_911),
.B1(n_897),
.B2(n_895),
.C(n_858),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_887),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_858),
.B(n_895),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_SL g935 ( 
.A1(n_867),
.A2(n_888),
.B(n_887),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_891),
.B(n_867),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_865),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_883),
.B(n_868),
.C(n_911),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_871),
.Y(n_939)
);

AOI211x1_ASAP7_75t_L g940 ( 
.A1(n_906),
.A2(n_881),
.B(n_853),
.C(n_852),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_897),
.B(n_866),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_893),
.B(n_908),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_906),
.B(n_879),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_889),
.A2(n_884),
.B(n_883),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_862),
.Y(n_946)
);

OAI22xp33_ASAP7_75t_L g947 ( 
.A1(n_877),
.A2(n_909),
.B1(n_874),
.B2(n_862),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_861),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_861),
.Y(n_949)
);

OR2x2_ASAP7_75t_SL g950 ( 
.A(n_890),
.B(n_882),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_891),
.B(n_890),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_868),
.A2(n_910),
.B1(n_900),
.B2(n_869),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_891),
.B(n_880),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_861),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_873),
.B(n_885),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_955),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_941),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_941),
.B(n_890),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_944),
.B(n_861),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_925),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_925),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_936),
.B(n_873),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_924),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_948),
.B(n_864),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_921),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_921),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_955),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_944),
.B(n_860),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_955),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_930),
.B(n_860),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_920),
.B(n_875),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_948),
.B(n_876),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_918),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_930),
.B(n_872),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_936),
.B(n_935),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_931),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_965),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_963),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_956),
.B(n_863),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_971),
.B(n_950),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_958),
.B(n_954),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_957),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_962),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_958),
.B(n_954),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_958),
.B(n_949),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_965),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_971),
.B(n_919),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_957),
.B(n_950),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_972),
.B(n_936),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_959),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_982),
.B(n_985),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_981),
.B(n_959),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_977),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_982),
.B(n_964),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_978),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_987),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_983),
.B(n_973),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_973),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_977),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_979),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_980),
.B(n_870),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_L g1003 ( 
.A(n_989),
.B(n_975),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_985),
.B(n_964),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_986),
.B(n_964),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_991),
.B(n_989),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_994),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_997),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_998),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_984),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_998),
.B(n_947),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_991),
.B(n_983),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_999),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_993),
.B(n_992),
.Y(n_1015)
);

AOI222xp33_ASAP7_75t_L g1016 ( 
.A1(n_1002),
.A2(n_932),
.B1(n_938),
.B2(n_952),
.C1(n_934),
.C2(n_942),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_898),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_993),
.B(n_986),
.Y(n_1018)
);

OAI221xp5_ASAP7_75t_SL g1019 ( 
.A1(n_995),
.A2(n_932),
.B1(n_934),
.B2(n_975),
.C(n_942),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_1019),
.A2(n_980),
.B(n_975),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1008),
.Y(n_1021)
);

AOI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_946),
.B(n_938),
.Y(n_1022)
);

OAI222xp33_ASAP7_75t_L g1023 ( 
.A1(n_1017),
.A2(n_1012),
.B1(n_1018),
.B2(n_1015),
.C1(n_1006),
.C2(n_1013),
.Y(n_1023)
);

NAND4xp25_ASAP7_75t_L g1024 ( 
.A(n_1010),
.B(n_940),
.C(n_968),
.D(n_970),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1007),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_1017),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1009),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_1014),
.A2(n_940),
.B1(n_1005),
.B2(n_1004),
.C(n_995),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1008),
.B(n_1005),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1011),
.B(n_994),
.Y(n_1031)
);

OAI322xp33_ASAP7_75t_L g1032 ( 
.A1(n_1026),
.A2(n_970),
.A3(n_968),
.B1(n_953),
.B2(n_923),
.C1(n_966),
.C2(n_976),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1023),
.A2(n_1011),
.B1(n_966),
.B2(n_935),
.C(n_976),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_1028),
.A2(n_1011),
.B(n_975),
.Y(n_1034)
);

OAI211xp5_ASAP7_75t_L g1035 ( 
.A1(n_1022),
.A2(n_915),
.B(n_863),
.C(n_956),
.Y(n_1035)
);

OAI32xp33_ASAP7_75t_L g1036 ( 
.A1(n_1029),
.A2(n_956),
.A3(n_898),
.B1(n_953),
.B2(n_920),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1025),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1020),
.A2(n_975),
.B1(n_936),
.B2(n_956),
.Y(n_1038)
);

NAND2x1_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_975),
.Y(n_1039)
);

AOI221xp5_ASAP7_75t_SL g1040 ( 
.A1(n_1034),
.A2(n_1024),
.B1(n_1027),
.B2(n_1031),
.C(n_1030),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_1032),
.A2(n_922),
.B(n_1021),
.C(n_939),
.Y(n_1041)
);

OAI211xp5_ASAP7_75t_L g1042 ( 
.A1(n_1033),
.A2(n_855),
.B(n_923),
.C(n_956),
.Y(n_1042)
);

AOI321xp33_ASAP7_75t_L g1043 ( 
.A1(n_1038),
.A2(n_1021),
.A3(n_990),
.B1(n_917),
.B2(n_919),
.C(n_951),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1035),
.A2(n_975),
.B(n_922),
.Y(n_1044)
);

AOI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_1036),
.A2(n_960),
.B1(n_961),
.B2(n_939),
.C(n_990),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1039),
.A2(n_917),
.B(n_918),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1037),
.B(n_1000),
.Y(n_1047)
);

NAND4xp25_ASAP7_75t_SL g1048 ( 
.A(n_1040),
.B(n_928),
.C(n_951),
.D(n_929),
.Y(n_1048)
);

OAI31xp33_ASAP7_75t_L g1049 ( 
.A1(n_1042),
.A2(n_929),
.A3(n_927),
.B(n_967),
.Y(n_1049)
);

NAND5xp2_ASAP7_75t_L g1050 ( 
.A(n_1043),
.B(n_927),
.C(n_926),
.D(n_967),
.E(n_969),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_1041),
.B(n_1045),
.C(n_1046),
.Y(n_1051)
);

NAND5xp2_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_926),
.C(n_967),
.D(n_969),
.E(n_960),
.Y(n_1052)
);

NAND4xp75_ASAP7_75t_L g1053 ( 
.A(n_1047),
.B(n_878),
.C(n_945),
.D(n_943),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_937),
.C(n_974),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1048),
.B(n_1001),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1049),
.B(n_984),
.Y(n_1056)
);

NOR4xp25_ASAP7_75t_L g1057 ( 
.A(n_1053),
.B(n_1050),
.C(n_1052),
.D(n_937),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1056),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1057),
.A2(n_1053),
.B1(n_936),
.B2(n_945),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1054),
.A2(n_974),
.B(n_936),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1055),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1054),
.B(n_984),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_1059),
.Y(n_1064)
);

XNOR2xp5_ASAP7_75t_L g1065 ( 
.A(n_1060),
.B(n_928),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1066),
.B(n_1062),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1067),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1068),
.B(n_1064),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_1069),
.A2(n_1066),
.B(n_1065),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1070),
.A2(n_1063),
.B1(n_1061),
.B2(n_933),
.Y(n_1071)
);


endmodule