module fake_jpeg_1142_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_24),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_25),
.B1(n_11),
.B2(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_5),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_20),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_13),
.B1(n_17),
.B2(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_39),
.C(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_45),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B(n_43),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B(n_48),
.Y(n_52)
);

NAND4xp25_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_28),
.C(n_36),
.D(n_31),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.A3(n_9),
.B1(n_37),
.B2(n_32),
.C1(n_17),
.C2(n_46),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_27),
.B(n_29),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_29),
.C(n_19),
.Y(n_55)
);


endmodule