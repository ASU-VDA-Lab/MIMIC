module fake_jpeg_3007_n_492 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_52),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_56),
.Y(n_123)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_6),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_95),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_93),
.Y(n_132)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_29),
.B(n_0),
.CON(n_90),
.SN(n_90)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_98),
.Y(n_119)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_94),
.A2(n_97),
.B(n_49),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_14),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_6),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_38),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_31),
.B(n_8),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_18),
.B1(n_35),
.B2(n_23),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_108),
.A2(n_128),
.B(n_145),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_46),
.B1(n_35),
.B2(n_23),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_109),
.A2(n_54),
.B1(n_49),
.B2(n_51),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_84),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_39),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_126),
.B(n_153),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_18),
.B1(n_35),
.B2(n_46),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_38),
.B1(n_48),
.B2(n_42),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_98),
.B1(n_31),
.B2(n_43),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_162),
.C(n_116),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_37),
.C(n_39),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_119),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_69),
.A2(n_18),
.B1(n_17),
.B2(n_44),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_36),
.B1(n_42),
.B2(n_48),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_17),
.B1(n_36),
.B2(n_44),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_59),
.B(n_47),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_161),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_47),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_168),
.B1(n_179),
.B2(n_109),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_103),
.B1(n_100),
.B2(n_74),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_98),
.A3(n_70),
.B1(n_83),
.B2(n_50),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_22),
.B1(n_50),
.B2(n_91),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_173),
.A2(n_194),
.B1(n_202),
.B2(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_105),
.B(n_22),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_185),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_180),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_187),
.Y(n_221)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_77),
.B1(n_87),
.B2(n_80),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_43),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_0),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_197),
.Y(n_229)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_192),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_99),
.B1(n_93),
.B2(n_53),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_1),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_200),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_203),
.B1(n_207),
.B2(n_158),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_43),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_115),
.B(n_53),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_211),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_134),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_133),
.B(n_112),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_99),
.B1(n_93),
.B2(n_70),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_132),
.A2(n_78),
.B1(n_66),
.B2(n_65),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_209),
.B1(n_143),
.B2(n_111),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_247),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_163),
.B1(n_131),
.B2(n_139),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_238),
.B1(n_242),
.B2(n_171),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_175),
.A2(n_128),
.B1(n_108),
.B2(n_145),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_222),
.A2(n_200),
.B1(n_191),
.B2(n_207),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_144),
.C(n_157),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_236),
.C(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_163),
.C(n_131),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_139),
.B1(n_122),
.B2(n_113),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_187),
.A2(n_127),
.B1(n_122),
.B2(n_143),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_133),
.C(n_127),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_222),
.B1(n_167),
.B2(n_184),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_197),
.B(n_111),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_210),
.C(n_180),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_248),
.B(n_249),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_250),
.B(n_257),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_258),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_198),
.B(n_180),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_265),
.B(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_210),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_267),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_165),
.C(n_201),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_249),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_204),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_188),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_180),
.B(n_190),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_219),
.B(n_204),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_190),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_271),
.B1(n_276),
.B2(n_262),
.Y(n_288)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_212),
.B(n_240),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_212),
.B(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_203),
.B1(n_193),
.B2(n_183),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_215),
.B1(n_234),
.B2(n_231),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_216),
.A2(n_247),
.B1(n_219),
.B2(n_220),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_236),
.B1(n_247),
.B2(n_243),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_205),
.B1(n_199),
.B2(n_186),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_239),
.B1(n_225),
.B2(n_217),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_181),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_215),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_250),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_251),
.A2(n_242),
.B1(n_235),
.B2(n_246),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_295),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_287),
.A2(n_297),
.B1(n_301),
.B2(n_271),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_288),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_213),
.B1(n_246),
.B2(n_237),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_298),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_307),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_235),
.B1(n_213),
.B2(n_237),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_213),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_260),
.A2(n_226),
.B1(n_217),
.B2(n_225),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_226),
.B1(n_245),
.B2(n_239),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_245),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_218),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_260),
.B1(n_268),
.B2(n_251),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_332),
.B1(n_286),
.B2(n_285),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_248),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_321),
.C(n_324),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_315),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_290),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_294),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_336),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_261),
.C(n_267),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_264),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_325),
.C(n_331),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_296),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_266),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_334),
.B1(n_292),
.B2(n_287),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_248),
.C(n_270),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_254),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_279),
.A2(n_273),
.B1(n_276),
.B2(n_262),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_279),
.A2(n_255),
.B1(n_265),
.B2(n_262),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_284),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_309),
.A2(n_282),
.B(n_283),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g371 ( 
.A1(n_337),
.A2(n_365),
.B(n_334),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_362),
.B1(n_269),
.B2(n_218),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_297),
.B1(n_291),
.B2(n_305),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_345),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_341),
.B(n_329),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_336),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_343),
.B(n_357),
.Y(n_370)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_295),
.B1(n_302),
.B2(n_301),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_283),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_348),
.Y(n_382)
);

BUFx12f_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_361),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_304),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_335),
.A2(n_288),
.B(n_300),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_316),
.B(n_308),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_289),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_356),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_333),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_333),
.A2(n_286),
.B1(n_281),
.B2(n_257),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_272),
.C(n_286),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_364),
.C(n_329),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_230),
.C(n_285),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_SL g365 ( 
.A(n_327),
.B(n_274),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_345),
.B(n_361),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_322),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_332),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_384),
.B(n_12),
.Y(n_411)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_358),
.B(n_330),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_378),
.B(n_385),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_368),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_10),
.C(n_2),
.Y(n_413)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_381),
.A2(n_387),
.B1(n_390),
.B2(n_372),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_326),
.C(n_328),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_363),
.C(n_356),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_344),
.A2(n_328),
.B(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_312),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_339),
.A2(n_259),
.B1(n_269),
.B2(n_205),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_392),
.B1(n_195),
.B2(n_178),
.Y(n_404)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_395),
.B(n_397),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_390),
.A2(n_359),
.B1(n_365),
.B2(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_409),
.B(n_381),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_370),
.A2(n_341),
.B1(n_364),
.B2(n_346),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_407),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_412),
.Y(n_420)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_170),
.C(n_182),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_405),
.B(n_406),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_51),
.C(n_27),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_375),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_51),
.C(n_27),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_382),
.C(n_386),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_8),
.B(n_12),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_27),
.B1(n_8),
.B2(n_9),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_373),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_411),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_9),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_413),
.B(n_384),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_1),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g419 ( 
.A(n_396),
.B(n_380),
.CI(n_379),
.CON(n_419),
.SN(n_419)
);

FAx1_ASAP7_75t_SL g422 ( 
.A(n_413),
.B(n_373),
.CI(n_389),
.CON(n_422),
.SN(n_422)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_422),
.A2(n_388),
.B1(n_406),
.B2(n_3),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_376),
.C(n_366),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_423),
.B(n_425),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_376),
.C(n_366),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_427),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_374),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_432),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_369),
.Y(n_429)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_435),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_415),
.A2(n_401),
.B1(n_404),
.B2(n_409),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_434),
.A2(n_437),
.B1(n_430),
.B2(n_426),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_397),
.C(n_399),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_421),
.A2(n_411),
.B(n_393),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_436),
.B(n_446),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_415),
.A2(n_411),
.B1(n_410),
.B2(n_398),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_399),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_420),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_412),
.C(n_408),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_444),
.C(n_435),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_442),
.A2(n_430),
.B1(n_432),
.B2(n_414),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_1),
.C(n_2),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_1),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_414),
.B(n_417),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_451),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_427),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_453),
.B(n_454),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_424),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_458),
.Y(n_469)
);

NAND2x1_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_424),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_462),
.B(n_446),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_442),
.B1(n_422),
.B2(n_419),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_426),
.C(n_431),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_448),
.C(n_440),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_416),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_439),
.Y(n_464)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_438),
.A2(n_419),
.B(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_463),
.B(n_2),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_467),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_471),
.B1(n_473),
.B2(n_474),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_434),
.C(n_437),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_454),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_444),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_472),
.B(n_452),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_1),
.B(n_2),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_455),
.C(n_456),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_477),
.B(n_479),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_R g477 ( 
.A(n_470),
.B(n_462),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_478),
.B(n_461),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_453),
.C(n_459),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_466),
.B(n_468),
.Y(n_482)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_483),
.A2(n_484),
.B(n_4),
.Y(n_487)
);

NAND4xp25_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_470),
.C(n_475),
.D(n_479),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_485),
.A2(n_3),
.B(n_4),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_486),
.A2(n_487),
.B(n_4),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_5),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_490),
.A2(n_488),
.B(n_5),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_5),
.Y(n_492)
);


endmodule