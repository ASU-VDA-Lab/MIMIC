module fake_jpeg_32019_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_54),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_20),
.B1(n_17),
.B2(n_15),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_3),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_12),
.B(n_19),
.C(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_51),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_16),
.B1(n_10),
.B2(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_52),
.B1(n_41),
.B2(n_47),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_3),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_68),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_42),
.Y(n_74)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_70),
.B(n_77),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_60),
.C(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_85),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_64),
.B(n_55),
.Y(n_84)
);

NAND2xp67_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_88),
.C(n_92),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_79),
.B1(n_84),
.B2(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_94),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_55),
.C(n_73),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_97),
.B1(n_73),
.B2(n_69),
.Y(n_103)
);

AOI21x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_55),
.B(n_76),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_58),
.Y(n_105)
);


endmodule