module fake_jpeg_41_n_68 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_24),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_38)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_44),
.B(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_31),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_1),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_37),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_57),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_10),
.B1(n_19),
.B2(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_56),
.B1(n_58),
.B2(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_59),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_57),
.B(n_8),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_6),
.B(n_9),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_11),
.Y(n_68)
);


endmodule