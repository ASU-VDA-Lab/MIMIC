module real_jpeg_31865_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_297;
wire n_209;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_295;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_1),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_1),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_2),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_3),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_4),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_10),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_10),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_12),
.B(n_33),
.Y(n_200)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_15),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

AND2x4_ASAP7_75t_SL g94 ( 
.A(n_16),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_16),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_16),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_181),
.Y(n_17)
);

NAND2xp33_ASAP7_75t_R g18 ( 
.A(n_19),
.B(n_180),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_125),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_22),
.B(n_125),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.C(n_108),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_23),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_24),
.B(n_44),
.C(n_53),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.C(n_39),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_25),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_193)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_34),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_35),
.B(n_39),
.Y(n_191)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_52),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_49),
.Y(n_156)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_51),
.Y(n_285)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_52),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_54),
.B(n_61),
.C(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_60),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_65),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_65),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_67),
.B(n_109),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_84),
.C(n_97),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_68),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_73),
.C(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_84),
.B(n_97),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_85),
.A2(n_86),
.B1(n_94),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_90),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_94),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_103),
.Y(n_112)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.C(n_113),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_120),
.C(n_123),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_157),
.B2(n_158),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_147),
.B2(n_148),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_201),
.B(n_297),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_184),
.B(n_186),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_188),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2x2_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_228),
.B(n_296),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_225),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_203),
.B(n_225),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_221),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_221),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.C(n_217),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_208),
.B1(n_217),
.B2(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_246),
.B(n_295),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_244),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_230),
.B(n_244),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.C(n_242),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_234),
.B1(n_242),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_261),
.B(n_294),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_258),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_258),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_250),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_254),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_287),
.B(n_293),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_282),
.B(n_286),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_276),
.B1(n_277),
.B2(n_281),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_276),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);


endmodule