module fake_netlist_6_1921_n_1800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1800;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_78),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_40),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_3),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_37),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_105),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_74),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_24),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_64),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_113),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_65),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_59),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_81),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_170),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_30),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_15),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_98),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_100),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_71),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_45),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_140),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_15),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_5),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_43),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_85),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_108),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_111),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_47),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_130),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_84),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_5),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_149),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_75),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_102),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_128),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_17),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_119),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_61),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_73),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_42),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_28),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_36),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_151),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_31),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_82),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_22),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_107),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_23),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_31),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_49),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_63),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_104),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_118),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_169),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_53),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_55),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_10),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_54),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_69),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_110),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_167),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_132),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_40),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_35),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_18),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_34),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_67),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_138),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_148),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_51),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_158),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_23),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_34),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_94),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_131),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_87),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_66),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_135),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_95),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_125),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_7),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_47),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_86),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_20),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_60),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_124),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_83),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_90),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_114),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_99),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_33),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_62),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_35),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_89),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_32),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_155),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_58),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_159),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_10),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_93),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_12),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_91),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_97),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_12),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_59),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_145),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_46),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_54),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_144),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_1),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_193),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_197),
.B(n_0),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_183),
.B(n_1),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_173),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_178),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_208),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_181),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_200),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_197),
.B(n_202),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_221),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_223),
.B(n_2),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_186),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_193),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_207),
.B(n_3),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_292),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_189),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_193),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_183),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_192),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_192),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_218),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_199),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_218),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_176),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_289),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_301),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_6),
.Y(n_379)
);

BUFx2_ASAP7_75t_SL g380 ( 
.A(n_210),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_269),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_269),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_335),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_301),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_202),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_209),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_209),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_343),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_203),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_205),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_177),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_247),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_247),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_248),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_248),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_251),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_215),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_251),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_274),
.B(n_6),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_254),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_254),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_227),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_196),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_256),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_228),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_231),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_256),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_261),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_270),
.B(n_8),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_232),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_179),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_234),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_239),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_196),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_241),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_242),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_261),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_243),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_272),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_245),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_255),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_281),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_281),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_279),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_290),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_346),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_270),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_345),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_271),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_362),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_363),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_271),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_366),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_367),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_368),
.B(n_230),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_373),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_387),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_353),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_380),
.B(n_287),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_374),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_380),
.B(n_388),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_371),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_388),
.B(n_287),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_391),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_364),
.B(n_235),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_399),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_407),
.B(n_174),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_400),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_364),
.B(n_235),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_349),
.B(n_245),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_394),
.B(n_210),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_405),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_406),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_409),
.B(n_291),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_382),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_410),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_225),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_414),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_416),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_402),
.B(n_225),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_365),
.B(n_268),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_240),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_417),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_419),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_327),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_436),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_448),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_454),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_454),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_379),
.C(n_360),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_480),
.B(n_268),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_455),
.B(n_369),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_459),
.B(n_365),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_459),
.B(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_467),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_467),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_455),
.B(n_354),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_498),
.A2(n_376),
.B1(n_429),
.B2(n_425),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_473),
.B(n_352),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_441),
.B(n_177),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_347),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_422),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_436),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_473),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_455),
.B(n_240),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_185),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_443),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_488),
.B(n_430),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_505),
.A2(n_348),
.B1(n_274),
.B2(n_293),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_445),
.B(n_449),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_458),
.B(n_424),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_462),
.B(n_415),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_479),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_479),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_450),
.B(n_352),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_458),
.B(n_358),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_463),
.B(n_195),
.Y(n_551)
);

NOR2x1p5_ASAP7_75t_L g552 ( 
.A(n_453),
.B(n_348),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_435),
.B(n_398),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_490),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_435),
.B(n_426),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_490),
.Y(n_558)
);

INVx4_ASAP7_75t_SL g559 ( 
.A(n_505),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_447),
.B(n_185),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_492),
.B(n_497),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_466),
.A2(n_339),
.B1(n_252),
.B2(n_224),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_447),
.B(n_198),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_494),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_461),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_470),
.B(n_184),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_500),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_492),
.B(n_201),
.Y(n_570)
);

INVx4_ASAP7_75t_SL g571 ( 
.A(n_505),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_492),
.B(n_220),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

INVx4_ASAP7_75t_SL g575 ( 
.A(n_505),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_432),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_466),
.B(n_401),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_492),
.B(n_264),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_473),
.B(n_403),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_403),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_434),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_478),
.B(n_404),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_448),
.B(n_404),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_497),
.B(n_319),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_198),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_474),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_507),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_432),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_475),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_477),
.B(n_259),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_478),
.B(n_408),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_483),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_497),
.B(n_448),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_468),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_437),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_497),
.B(n_191),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_451),
.B(n_408),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_484),
.B(n_259),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_451),
.B(n_182),
.C(n_180),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_491),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_411),
.Y(n_608)
);

BUFx4f_ASAP7_75t_L g609 ( 
.A(n_505),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_432),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_499),
.B(n_411),
.Y(n_612)
);

OR2x2_ASAP7_75t_SL g613 ( 
.A(n_482),
.B(n_284),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_505),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_495),
.B(n_329),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_476),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_438),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_503),
.B(n_259),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_438),
.Y(n_619)
);

AND3x4_ASAP7_75t_L g620 ( 
.A(n_476),
.B(n_273),
.C(n_262),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_469),
.B(n_191),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_482),
.B(n_216),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_439),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_439),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_440),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_440),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_468),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_504),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_442),
.B(n_412),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_501),
.B(n_277),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_442),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_468),
.B(n_277),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_456),
.B(n_262),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_444),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_444),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_446),
.B(n_206),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_505),
.B(n_327),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_446),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_469),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_469),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_471),
.B(n_428),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_471),
.B(n_206),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_481),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_471),
.B(n_226),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_471),
.B(n_216),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_456),
.B(n_412),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_481),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_481),
.B(n_277),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_481),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_481),
.B(n_217),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_481),
.B(n_217),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_456),
.A2(n_253),
.B1(n_295),
.B2(n_265),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_460),
.A2(n_330),
.B1(n_341),
.B2(n_284),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_487),
.Y(n_657)
);

INVxp33_ASAP7_75t_L g658 ( 
.A(n_460),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_460),
.A2(n_286),
.B1(n_293),
.B2(n_304),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_561),
.B(n_487),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_608),
.B(n_356),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_561),
.B(n_487),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_524),
.B(n_327),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_612),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_508),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_530),
.B(n_487),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_524),
.B(n_327),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_530),
.B(n_615),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_615),
.B(n_520),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_511),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_600),
.B(n_487),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_524),
.B(n_614),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_548),
.B(n_244),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_512),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_538),
.A2(n_306),
.B1(n_246),
.B2(n_250),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_630),
.B(n_359),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_527),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_644),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_600),
.B(n_570),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_513),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_630),
.B(n_377),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_570),
.B(n_487),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_489),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_489),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_557),
.B(n_384),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_578),
.B(n_489),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_577),
.A2(n_286),
.B(n_304),
.C(n_324),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_524),
.B(n_299),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_527),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_515),
.A2(n_514),
.B1(n_510),
.B2(n_537),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_557),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_549),
.B(n_273),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_614),
.B(n_305),
.Y(n_693)
);

INVxp33_ASAP7_75t_L g694 ( 
.A(n_541),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_578),
.B(n_489),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_541),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_521),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_532),
.B(n_390),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_588),
.B(n_489),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_588),
.B(n_489),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_538),
.B(n_244),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_523),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_510),
.B(n_246),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_510),
.B(n_250),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_188),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_510),
.B(n_263),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_535),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_614),
.B(n_307),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_563),
.B(n_540),
.C(n_551),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_554),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_542),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_537),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_537),
.A2(n_263),
.B1(n_267),
.B2(n_276),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_529),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_522),
.B(n_190),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_614),
.B(n_309),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_635),
.B(n_266),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_543),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_515),
.A2(n_310),
.B1(n_311),
.B2(n_321),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_509),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_609),
.B(n_559),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_510),
.B(n_266),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_546),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_509),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_528),
.B(n_603),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_567),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_528),
.A2(n_320),
.B1(n_276),
.B2(n_278),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_558),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_658),
.B(n_562),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_609),
.B(n_322),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_565),
.B(n_267),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_568),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_595),
.B(n_323),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_526),
.B(n_238),
.C(n_257),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_536),
.B(n_204),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_569),
.B(n_580),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_288),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_544),
.B(n_211),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_212),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_605),
.B(n_213),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_517),
.A2(n_324),
.B(n_330),
.C(n_341),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_647),
.A2(n_642),
.B(n_641),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_613),
.A2(n_306),
.B1(n_278),
.B2(n_297),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_586),
.B(n_297),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_579),
.B(n_421),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_590),
.B(n_298),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_559),
.B(n_336),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_563),
.B(n_233),
.C(n_229),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_618),
.B(n_222),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_593),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_602),
.B(n_298),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_617),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_517),
.B(n_236),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_559),
.B(n_340),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_583),
.B(n_237),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_619),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_581),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_528),
.A2(n_302),
.B1(n_333),
.B2(n_325),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_623),
.B(n_300),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_632),
.B(n_249),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_550),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_624),
.B(n_300),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_598),
.A2(n_423),
.B(n_427),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_571),
.B(n_302),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_528),
.A2(n_320),
.B1(n_308),
.B2(n_314),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_571),
.B(n_308),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_635),
.B(n_314),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_550),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_625),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_325),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_598),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_650),
.A2(n_496),
.B(n_485),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_621),
.A2(n_331),
.B1(n_333),
.B2(n_258),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_518),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_571),
.B(n_331),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_464),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_525),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_637),
.B(n_464),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_531),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_648),
.A2(n_427),
.B(n_423),
.C(n_428),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_529),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_525),
.B(n_464),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_528),
.B(n_465),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_640),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_575),
.B(n_277),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_643),
.B(n_465),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_553),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_653),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_595),
.B(n_288),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_575),
.B(n_496),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_647),
.B(n_465),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_599),
.B(n_288),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_603),
.B(n_472),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_606),
.B(n_317),
.C(n_275),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_472),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_653),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_621),
.A2(n_318),
.B1(n_280),
.B2(n_282),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_518),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_599),
.B(n_288),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_654),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_603),
.B(n_472),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_575),
.B(n_496),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_604),
.B(n_485),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_648),
.A2(n_385),
.B(n_383),
.C(n_328),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_518),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_315),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_553),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_654),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_622),
.B(n_316),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_539),
.B(n_260),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_604),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_545),
.B(n_646),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_529),
.B(n_283),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_635),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_622),
.B(n_326),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_566),
.B(n_285),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_332),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_533),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_573),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_533),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_677),
.B(n_689),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_709),
.B(n_582),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_714),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_668),
.A2(n_679),
.B(n_796),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_691),
.A2(n_645),
.B(n_634),
.C(n_651),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_714),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_694),
.B(n_591),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_709),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_669),
.A2(n_552),
.B1(n_622),
.B2(n_628),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_714),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_785),
.B(n_631),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_696),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_785),
.B(n_631),
.Y(n_841)
);

AOI21xp33_ASAP7_75t_L g842 ( 
.A1(n_707),
.A2(n_607),
.B(n_616),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_677),
.B(n_516),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_689),
.B(n_516),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_712),
.B(n_585),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_690),
.A2(n_657),
.B1(n_652),
.B2(n_639),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_826),
.B(n_627),
.Y(n_847)
);

AO21x1_ASAP7_75t_L g848 ( 
.A1(n_704),
.A2(n_645),
.B(n_638),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_828),
.A2(n_759),
.B(n_744),
.C(n_754),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_664),
.B(n_655),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_701),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_660),
.A2(n_650),
.B(n_547),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_711),
.A2(n_620),
.B1(n_627),
.B2(n_629),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_662),
.A2(n_547),
.B(n_596),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_701),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_678),
.B(n_629),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_666),
.A2(n_596),
.B(n_601),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_671),
.A2(n_601),
.B(n_611),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_799),
.A2(n_672),
.B(n_682),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_698),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_804),
.A2(n_638),
.B(n_589),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_685),
.A2(n_589),
.B1(n_574),
.B2(n_610),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_678),
.A2(n_708),
.B1(n_724),
.B2(n_705),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_741),
.B(n_656),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_820),
.A2(n_534),
.B(n_560),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_790),
.B(n_573),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_675),
.A2(n_659),
.B1(n_656),
.B2(n_294),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_661),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_798),
.A2(n_564),
.B(n_560),
.C(n_534),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_672),
.A2(n_611),
.B(n_601),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_750),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_706),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_808),
.A2(n_564),
.B(n_594),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_761),
.B(n_659),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_790),
.B(n_594),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_706),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_683),
.A2(n_611),
.B(n_576),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_720),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_733),
.B(n_576),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_385),
.B(n_328),
.C(n_342),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_719),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_684),
.A2(n_344),
.B(n_338),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_702),
.A2(n_328),
.B1(n_337),
.B2(n_313),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_824),
.B(n_729),
.Y(n_885)
);

O2A1O1Ixp5_ASAP7_75t_L g886 ( 
.A1(n_734),
.A2(n_328),
.B(n_303),
.C(n_296),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_816),
.B(n_9),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_720),
.B(n_13),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_686),
.A2(n_171),
.B(n_168),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_728),
.B(n_13),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_728),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_695),
.A2(n_165),
.B(n_163),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_820),
.A2(n_160),
.B(n_146),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_747),
.A2(n_134),
.B(n_127),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_797),
.B(n_121),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_699),
.A2(n_120),
.B(n_116),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_736),
.B(n_14),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_736),
.B(n_14),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_SL g899 ( 
.A1(n_798),
.A2(n_16),
.B(n_19),
.C(n_21),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_700),
.A2(n_101),
.B(n_96),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_800),
.B(n_807),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_716),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_727),
.A2(n_88),
.B(n_80),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_727),
.A2(n_77),
.B(n_76),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_723),
.A2(n_72),
.B(n_70),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_791),
.A2(n_68),
.B(n_19),
.Y(n_906)
);

CKINVDCx10_ASAP7_75t_R g907 ( 
.A(n_719),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_743),
.A2(n_16),
.B(n_24),
.C(n_25),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_730),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_811),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_723),
.A2(n_36),
.B(n_39),
.Y(n_911)
);

BUFx2_ASAP7_75t_SL g912 ( 
.A(n_822),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_789),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_764),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_756),
.B(n_44),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_756),
.B(n_48),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_758),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_SL g918 ( 
.A1(n_810),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_758),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_762),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_673),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_794),
.A2(n_50),
.B(n_52),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_762),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_781),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_776),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_776),
.B(n_665),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_670),
.B(n_52),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_772),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_674),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_792),
.Y(n_931)
);

NOR2x1_ASAP7_75t_SL g932 ( 
.A(n_810),
.B(n_56),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_717),
.B(n_58),
.C(n_753),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_721),
.A2(n_778),
.B1(n_765),
.B2(n_763),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_680),
.B(n_697),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_801),
.A2(n_809),
.B(n_803),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_811),
.A2(n_819),
.B1(n_739),
.B2(n_818),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_703),
.B(n_713),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_748),
.A2(n_746),
.B(n_687),
.C(n_769),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_676),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_784),
.A2(n_786),
.B(n_740),
.Y(n_941)
);

O2A1O1Ixp5_ASAP7_75t_L g942 ( 
.A1(n_793),
.A2(n_752),
.B(n_760),
.C(n_718),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_681),
.A2(n_725),
.B1(n_755),
.B2(n_745),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_731),
.B(n_732),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_742),
.B(n_738),
.C(n_767),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_781),
.B(n_813),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_781),
.B(n_813),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_735),
.A2(n_757),
.B(n_766),
.C(n_751),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_806),
.B(n_813),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_806),
.A2(n_813),
.B(n_760),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_722),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_806),
.A2(n_752),
.B(n_827),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_821),
.B(n_802),
.C(n_805),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_792),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_806),
.A2(n_827),
.B(n_768),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_827),
.A2(n_726),
.B(n_775),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_822),
.B(n_782),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_692),
.B(n_673),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_770),
.B(n_737),
.C(n_780),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_673),
.B(n_749),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_777),
.B(n_795),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_814),
.A2(n_825),
.B1(n_823),
.B2(n_817),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_719),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_719),
.A2(n_774),
.B1(n_715),
.B2(n_793),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_722),
.A2(n_775),
.B(n_768),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_774),
.B(n_775),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_726),
.B(n_815),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_774),
.A2(n_771),
.B1(n_783),
.B2(n_773),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_688),
.A2(n_718),
.B(n_710),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_688),
.A2(n_693),
.B(n_710),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_774),
.Y(n_971)
);

OAI321xp33_ASAP7_75t_L g972 ( 
.A1(n_812),
.A2(n_788),
.A3(n_773),
.B1(n_771),
.B2(n_783),
.C(n_693),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_787),
.A2(n_663),
.B1(n_667),
.B2(n_779),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_663),
.A2(n_668),
.B(n_691),
.C(n_702),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_787),
.B(n_667),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_668),
.B(n_669),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_660),
.A2(n_609),
.B(n_662),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_701),
.Y(n_978)
);

BUFx8_ASAP7_75t_L g979 ( 
.A(n_698),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_714),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_691),
.B(n_696),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_701),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_701),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_668),
.B(n_669),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_668),
.A2(n_675),
.B1(n_691),
.B2(n_696),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_660),
.A2(n_609),
.B(n_662),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_668),
.B(n_785),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_668),
.B(n_785),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_668),
.A2(n_675),
.B1(n_691),
.B2(n_696),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_714),
.B(n_723),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_820),
.A2(n_747),
.B(n_726),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_714),
.Y(n_992)
);

CKINVDCx10_ASAP7_75t_R g993 ( 
.A(n_709),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_714),
.B(n_723),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_660),
.A2(n_609),
.B(n_662),
.Y(n_995)
);

INVx11_ASAP7_75t_L g996 ( 
.A(n_709),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_668),
.A2(n_669),
.B1(n_515),
.B2(n_679),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_714),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_820),
.A2(n_747),
.B(n_726),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_709),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_668),
.B(n_785),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_668),
.B(n_785),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_668),
.A2(n_675),
.B1(n_691),
.B2(n_696),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_714),
.B(n_723),
.Y(n_1004)
);

AO22x1_ASAP7_75t_L g1005 ( 
.A1(n_668),
.A2(n_669),
.B1(n_694),
.B2(n_753),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_698),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_709),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_668),
.A2(n_675),
.B1(n_691),
.B2(n_696),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_668),
.A2(n_691),
.B(n_702),
.C(n_696),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_677),
.B(n_689),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_996),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_997),
.A2(n_984),
.B(n_976),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_987),
.B(n_988),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_856),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1001),
.B(n_1002),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_978),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_SL g1017 ( 
.A1(n_887),
.A2(n_890),
.B(n_888),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_936),
.A2(n_860),
.B(n_960),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_872),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_952),
.A2(n_965),
.B(n_858),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_849),
.A2(n_832),
.B(n_942),
.C(n_1005),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_867),
.A2(n_876),
.B(n_862),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_851),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_928),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_832),
.B(n_875),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_937),
.A2(n_989),
.B1(n_1008),
.B2(n_985),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_928),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_941),
.A2(n_948),
.B(n_874),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_956),
.A2(n_859),
.B(n_855),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_839),
.B(n_841),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_865),
.B(n_985),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_989),
.A2(n_1008),
.B1(n_1003),
.B2(n_945),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_885),
.A2(n_958),
.B1(n_953),
.B2(n_1003),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_874),
.A2(n_864),
.B(n_853),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_878),
.A2(n_950),
.B(n_955),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_940),
.A2(n_943),
.B1(n_837),
.B2(n_840),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_921),
.B(n_957),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_1000),
.B(n_933),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_969),
.A2(n_970),
.B(n_967),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_957),
.B(n_829),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_981),
.B(n_1009),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_926),
.B(n_935),
.Y(n_1042)
);

O2A1O1Ixp5_ASAP7_75t_L g1043 ( 
.A1(n_922),
.A2(n_886),
.B(n_915),
.C(n_897),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_870),
.A2(n_962),
.B(n_974),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_938),
.B(n_944),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_SL g1046 ( 
.A(n_924),
.B(n_928),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_846),
.A2(n_857),
.B(n_847),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_833),
.A2(n_961),
.B(n_975),
.Y(n_1048)
);

NAND2x1_ASAP7_75t_L g1049 ( 
.A(n_951),
.B(n_831),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_871),
.A2(n_893),
.B(n_1004),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_924),
.B(n_831),
.Y(n_1051)
);

AND2x6_ASAP7_75t_L g1052 ( 
.A(n_966),
.B(n_951),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_873),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_880),
.A2(n_901),
.B(n_924),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_861),
.B(n_835),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_877),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_939),
.A2(n_863),
.B(n_854),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_861),
.B(n_869),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_982),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_879),
.A2(n_919),
.B(n_891),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_968),
.A2(n_923),
.B(n_920),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_990),
.A2(n_994),
.B(n_894),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_946),
.A2(n_947),
.B(n_949),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_924),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_834),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1006),
.B(n_845),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_964),
.A2(n_895),
.B(n_968),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_930),
.A2(n_1006),
.B1(n_925),
.B2(n_917),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_959),
.A2(n_829),
.B1(n_1010),
.B2(n_934),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_913),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_834),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1010),
.B(n_983),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_946),
.A2(n_947),
.B(n_949),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_903),
.A2(n_904),
.B(n_954),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_922),
.A2(n_916),
.B(n_898),
.C(n_906),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_842),
.B(n_850),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_964),
.A2(n_972),
.B(n_934),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_931),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_927),
.B(n_883),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_SL g1080 ( 
.A1(n_971),
.A2(n_972),
.B(n_899),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_908),
.A2(n_932),
.A3(n_914),
.B(n_909),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_905),
.A2(n_892),
.B(n_900),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_868),
.B(n_980),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1007),
.B(n_963),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_834),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_884),
.B(n_902),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_905),
.A2(n_881),
.B(n_889),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_836),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_838),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_838),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_SL g1091 ( 
.A1(n_998),
.A2(n_992),
.B(n_838),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_SL g1092 ( 
.A1(n_910),
.A2(n_843),
.B(n_844),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_868),
.B(n_852),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_912),
.B(n_852),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_852),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_896),
.A2(n_882),
.B(n_911),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_918),
.A2(n_929),
.B(n_914),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_882),
.A2(n_998),
.B(n_992),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_980),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_830),
.B(n_992),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_909),
.A2(n_929),
.B(n_979),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_979),
.A2(n_907),
.B(n_993),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_987),
.B(n_668),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_997),
.A2(n_668),
.B(n_694),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_872),
.B(n_691),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_987),
.B(n_668),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_987),
.B(n_668),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_848),
.A2(n_668),
.B(n_849),
.C(n_977),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_987),
.B(n_668),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_987),
.B(n_668),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_921),
.B(n_957),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_836),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_872),
.B(n_691),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_997),
.B(n_668),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_977),
.A2(n_995),
.B(n_986),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_872),
.B(n_691),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_921),
.B(n_957),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_830),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_856),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_849),
.A2(n_668),
.B(n_832),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_872),
.B(n_691),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_997),
.A2(n_668),
.B1(n_849),
.B2(n_987),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_851),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_997),
.A2(n_691),
.B1(n_696),
.B2(n_620),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_991),
.A2(n_999),
.B(n_866),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_869),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_976),
.B(n_668),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_987),
.B(n_668),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_991),
.A2(n_999),
.B(n_866),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_987),
.B(n_668),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_991),
.A2(n_999),
.B(n_866),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_887),
.A2(n_705),
.B(n_704),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_SL g1133 ( 
.A(n_997),
.B(n_668),
.C(n_849),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_836),
.B(n_709),
.Y(n_1134)
);

BUFx12f_ASAP7_75t_L g1135 ( 
.A(n_979),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_849),
.A2(n_668),
.B(n_832),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_849),
.A2(n_668),
.B(n_832),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_997),
.A2(n_668),
.B1(n_849),
.B2(n_987),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_836),
.B(n_709),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_997),
.B(n_668),
.C(n_480),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_987),
.B(n_668),
.Y(n_1141)
);

OAI22x1_ASAP7_75t_L g1142 ( 
.A1(n_997),
.A2(n_668),
.B1(n_696),
.B2(n_669),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_976),
.B(n_668),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_872),
.Y(n_1144)
);

AO21x1_ASAP7_75t_L g1145 ( 
.A1(n_997),
.A2(n_668),
.B(n_976),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_987),
.B(n_668),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_849),
.A2(n_668),
.B(n_832),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_848),
.A2(n_973),
.A3(n_986),
.B(n_977),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1026),
.A2(n_1077),
.B1(n_1107),
.B2(n_1130),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1040),
.B(n_1037),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1064),
.B(n_1024),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1077),
.A2(n_1108),
.B(n_1021),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1055),
.B(n_1105),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1127),
.B(n_1143),
.Y(n_1157)
);

NOR2xp67_ASAP7_75t_L g1158 ( 
.A(n_1011),
.B(n_1118),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1110),
.B(n_1128),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1064),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1112),
.Y(n_1161)
);

AOI222xp33_ASAP7_75t_L g1162 ( 
.A1(n_1032),
.A2(n_1114),
.B1(n_1140),
.B2(n_1031),
.C1(n_1076),
.C2(n_1142),
.Y(n_1162)
);

BUFx8_ASAP7_75t_SL g1163 ( 
.A(n_1135),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1033),
.A2(n_1146),
.B1(n_1141),
.B2(n_1139),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1025),
.B(n_1030),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1011),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1016),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1019),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1144),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1067),
.A2(n_1136),
.B(n_1147),
.C(n_1120),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1013),
.B(n_1015),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1172)
);

INVxp67_ASAP7_75t_SL g1173 ( 
.A(n_1046),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1028),
.A2(n_1082),
.B(n_1044),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1076),
.B(n_1104),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1027),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1126),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1040),
.B(n_1037),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1119),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_1064),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1078),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1121),
.B(n_1066),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1028),
.A2(n_1082),
.B(n_1044),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1111),
.B(n_1117),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1023),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1053),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1056),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1134),
.B(n_1058),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1059),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1070),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1064),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1123),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1034),
.A2(n_1042),
.B(n_1079),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1072),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_1137),
.B(n_1045),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1027),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1124),
.B(n_1086),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1122),
.A2(n_1138),
.B(n_1133),
.C(n_1041),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1145),
.B(n_1012),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1133),
.A2(n_1124),
.B1(n_1067),
.B2(n_1101),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1083),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1070),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1100),
.B(n_1111),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1093),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1117),
.B(n_1084),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1057),
.B(n_1069),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1088),
.B(n_1036),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1089),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1090),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1022),
.B(n_1052),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1094),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1051),
.Y(n_1212)
);

AND2x6_ASAP7_75t_L g1213 ( 
.A(n_1027),
.B(n_1065),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1092),
.B(n_1038),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1098),
.B(n_1094),
.Y(n_1215)
);

AOI211xp5_ASAP7_75t_L g1216 ( 
.A1(n_1087),
.A2(n_1068),
.B(n_1096),
.C(n_1061),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1060),
.A2(n_1094),
.B1(n_1022),
.B2(n_1096),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1021),
.A2(n_1043),
.B(n_1075),
.C(n_1108),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1098),
.B(n_1071),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1085),
.B(n_1081),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1052),
.B(n_1048),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1071),
.B(n_1095),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1102),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1065),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1027),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1115),
.A2(n_1047),
.B(n_1075),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1065),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1065),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1051),
.A2(n_1097),
.B(n_1054),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1081),
.B(n_1102),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1074),
.A2(n_1035),
.B(n_1020),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1099),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1097),
.A2(n_1054),
.B(n_1099),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1095),
.B(n_1024),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1043),
.A2(n_1029),
.B(n_1091),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1081),
.B(n_1099),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1099),
.Y(n_1237)
);

NAND2x1_ASAP7_75t_L g1238 ( 
.A(n_1052),
.B(n_1073),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1052),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1052),
.B(n_1081),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1063),
.B(n_1062),
.Y(n_1241)
);

O2A1O1Ixp5_ASAP7_75t_SL g1242 ( 
.A1(n_1017),
.A2(n_1132),
.B(n_1080),
.C(n_1148),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1049),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1080),
.A2(n_1017),
.B1(n_1132),
.B2(n_1148),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_SL g1245 ( 
.A(n_1050),
.B(n_1125),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1129),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1131),
.B(n_1055),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1039),
.A2(n_609),
.B(n_1018),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1040),
.B(n_1037),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1014),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1077),
.A2(n_668),
.B(n_669),
.C(n_997),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1127),
.B(n_668),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1027),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1112),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1135),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1055),
.B(n_1105),
.Y(n_1258)
);

BUFx2_ASAP7_75t_R g1259 ( 
.A(n_1102),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1014),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1026),
.A2(n_849),
.B(n_1032),
.C(n_1133),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_L g1262 ( 
.A(n_1135),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1027),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1040),
.B(n_1037),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1064),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1032),
.A2(n_563),
.B1(n_1026),
.B2(n_668),
.C(n_691),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1032),
.A2(n_668),
.B(n_984),
.C(n_976),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1032),
.A2(n_668),
.B1(n_515),
.B2(n_1140),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1026),
.A2(n_997),
.B1(n_668),
.B2(n_1077),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1014),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1027),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1026),
.A2(n_997),
.B1(n_668),
.B2(n_1077),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1127),
.B(n_668),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1014),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1026),
.A2(n_997),
.B1(n_668),
.B2(n_1077),
.Y(n_1280)
);

INVx8_ASAP7_75t_L g1281 ( 
.A(n_1064),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1032),
.A2(n_668),
.B1(n_515),
.B2(n_1140),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1014),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1144),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1064),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1135),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1236),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1169),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1220),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1175),
.A2(n_1268),
.B1(n_1253),
.B2(n_1278),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1240),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1257),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1157),
.A2(n_1280),
.B1(n_1277),
.B2(n_1273),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1155),
.B(n_1159),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1229),
.B(n_1233),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1281),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1251),
.Y(n_1298)
);

BUFx2_ASAP7_75t_SL g1299 ( 
.A(n_1196),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1272),
.A2(n_1282),
.B1(n_1171),
.B2(n_1248),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1286),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1166),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1273),
.A2(n_1280),
.B1(n_1277),
.B2(n_1206),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1171),
.A2(n_1270),
.B1(n_1266),
.B2(n_1248),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1235),
.A2(n_1231),
.B(n_1249),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1275),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1240),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1156),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1238),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1279),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1206),
.A2(n_1214),
.B1(n_1223),
.B2(n_1230),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1281),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1256),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1241),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1162),
.A2(n_1164),
.B1(n_1200),
.B2(n_1149),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1162),
.A2(n_1149),
.B1(n_1197),
.B2(n_1204),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1241),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1283),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1239),
.B(n_1247),
.Y(n_1319)
);

CKINVDCx16_ASAP7_75t_R g1320 ( 
.A(n_1161),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1284),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1151),
.A2(n_1274),
.B1(n_1254),
.B2(n_1270),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1165),
.B(n_1201),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1244),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1207),
.A2(n_1182),
.B1(n_1188),
.B2(n_1199),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1151),
.A2(n_1263),
.B1(n_1271),
.B2(n_1254),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1211),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1154),
.A2(n_1258),
.B1(n_1263),
.B2(n_1266),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1244),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_1168),
.Y(n_1330)
);

BUFx8_ASAP7_75t_SL g1331 ( 
.A(n_1163),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1217),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1165),
.B(n_1252),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1217),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1210),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1284),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1190),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1271),
.A2(n_1274),
.B1(n_1172),
.B2(n_1221),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1210),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1202),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1224),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1177),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1179),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1184),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1194),
.A2(n_1215),
.B1(n_1262),
.B2(n_1158),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1219),
.B(n_1246),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1170),
.B(n_1153),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1180),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1260),
.Y(n_1349)
);

INVxp33_ASAP7_75t_L g1350 ( 
.A(n_1205),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1261),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1180),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1187),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1262),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1281),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1215),
.B(n_1212),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1269),
.A2(n_1198),
.B(n_1195),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1203),
.B(n_1150),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1189),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1208),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1178),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1215),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1153),
.Y(n_1363)
);

AO21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1243),
.A2(n_1225),
.B(n_1227),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1178),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1208),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1267),
.Y(n_1367)
);

AO21x1_ASAP7_75t_L g1368 ( 
.A1(n_1216),
.A2(n_1174),
.B(n_1183),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1193),
.A2(n_1226),
.B(n_1242),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1250),
.A2(n_1265),
.B1(n_1173),
.B2(n_1192),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1218),
.Y(n_1372)
);

INVx6_ASAP7_75t_L g1373 ( 
.A(n_1267),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1267),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1250),
.A2(n_1265),
.B1(n_1186),
.B2(n_1181),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1246),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1209),
.A2(n_1185),
.B(n_1245),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1245),
.A2(n_1246),
.B(n_1222),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1212),
.A2(n_1234),
.B1(n_1232),
.B2(n_1285),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1246),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1259),
.A2(n_1228),
.B1(n_1196),
.B2(n_1237),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1160),
.B(n_1285),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1234),
.A2(n_1213),
.B(n_1259),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1191),
.B(n_1276),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1213),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1152),
.A2(n_1196),
.B(n_1228),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1176),
.A2(n_1255),
.B1(n_1264),
.B2(n_1276),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1226),
.A2(n_1235),
.B(n_1077),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1167),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1257),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1238),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1238),
.B(n_1239),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1253),
.A2(n_668),
.B1(n_1278),
.B2(n_997),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1236),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1236),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1290),
.B(n_1322),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_L g1397 ( 
.A(n_1348),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1321),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1370),
.A2(n_1305),
.B(n_1357),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1308),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1393),
.A2(n_1293),
.B1(n_1300),
.B2(n_1315),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1287),
.B(n_1395),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1360),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1332),
.B(n_1334),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1322),
.A2(n_1371),
.B1(n_1294),
.B2(n_1350),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1356),
.B(n_1314),
.Y(n_1406)
);

INVxp33_ASAP7_75t_SL g1407 ( 
.A(n_1313),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1287),
.B(n_1395),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1304),
.B(n_1326),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1378),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1394),
.B(n_1289),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1308),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1356),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1378),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1356),
.B(n_1314),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1324),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1356),
.B(n_1314),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1323),
.B(n_1328),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1329),
.Y(n_1419)
);

NOR2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1385),
.B(n_1348),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1323),
.B(n_1338),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1358),
.B(n_1313),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1291),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1355),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1366),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1332),
.B(n_1334),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1307),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1333),
.B(n_1336),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1288),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1309),
.A2(n_1391),
.B(n_1368),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_SL g1431 ( 
.A(n_1302),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1394),
.B(n_1289),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1388),
.A2(n_1372),
.B(n_1376),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1317),
.B(n_1362),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1343),
.Y(n_1435)
);

NOR2x1_ASAP7_75t_L g1436 ( 
.A(n_1345),
.B(n_1295),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1337),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1388),
.A2(n_1372),
.B(n_1376),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1388),
.A2(n_1380),
.B(n_1363),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1340),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1342),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1335),
.B(n_1339),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1295),
.B(n_1362),
.Y(n_1444)
);

AO21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1303),
.A2(n_1316),
.B(n_1347),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1377),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1319),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1377),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1377),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1335),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1355),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1339),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1347),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1333),
.A2(n_1351),
.B(n_1349),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1353),
.B(n_1359),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1330),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1344),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1319),
.B(n_1297),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1298),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1351),
.A2(n_1325),
.B(n_1359),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1373),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1353),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1298),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1306),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1409),
.B(n_1311),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_R g1466 ( 
.A(n_1454),
.B(n_1383),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1454),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1454),
.B(n_1383),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1383),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1444),
.B(n_1392),
.Y(n_1470)
);

INVx2_ASAP7_75t_R g1471 ( 
.A(n_1446),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1453),
.B(n_1310),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_L g1473 ( 
.A(n_1436),
.B(n_1383),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1440),
.B(n_1392),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1401),
.A2(n_1375),
.B1(n_1365),
.B2(n_1379),
.C(n_1302),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1399),
.B(n_1346),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1405),
.B(n_1396),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1403),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1410),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1433),
.B(n_1438),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1410),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1438),
.B(n_1318),
.Y(n_1482)
);

AND2x4_ASAP7_75t_SL g1483 ( 
.A(n_1444),
.B(n_1369),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1443),
.B(n_1310),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1443),
.B(n_1389),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1448),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1449),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1416),
.B(n_1364),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1429),
.B(n_1361),
.C(n_1387),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1299),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1414),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1419),
.B(n_1382),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1439),
.B(n_1384),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1478),
.B(n_1428),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1478),
.B(n_1425),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1473),
.B(n_1397),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1477),
.A2(n_1436),
.B(n_1381),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1437),
.Y(n_1501)
);

OAI221xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1465),
.A2(n_1418),
.B1(n_1421),
.B2(n_1442),
.C(n_1457),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1489),
.A2(n_1444),
.B1(n_1398),
.B2(n_1413),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1473),
.B(n_1397),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1493),
.B(n_1456),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1493),
.B(n_1441),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1484),
.B(n_1400),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1489),
.A2(n_1445),
.B1(n_1413),
.B2(n_1415),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1475),
.B(n_1400),
.C(n_1412),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1475),
.A2(n_1412),
.B1(n_1422),
.B2(n_1455),
.C(n_1458),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1469),
.A2(n_1444),
.B1(n_1447),
.B2(n_1404),
.C(n_1426),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1490),
.A2(n_1397),
.B1(n_1461),
.B2(n_1341),
.C(n_1451),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1488),
.A2(n_1420),
.B(n_1435),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1432),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_SL g1515 ( 
.A(n_1490),
.B(n_1398),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1488),
.A2(n_1420),
.B(n_1435),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1490),
.A2(n_1445),
.B1(n_1413),
.B2(n_1415),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1472),
.B(n_1413),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1466),
.B(n_1459),
.C(n_1460),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1460),
.C(n_1463),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1470),
.A2(n_1431),
.B1(n_1423),
.B2(n_1427),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1476),
.A2(n_1430),
.B(n_1460),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1485),
.B(n_1455),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1485),
.B(n_1455),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1490),
.A2(n_1415),
.B1(n_1417),
.B2(n_1406),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1472),
.B(n_1320),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1479),
.B(n_1481),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1479),
.B(n_1434),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1450),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1480),
.B(n_1460),
.C(n_1464),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1479),
.B(n_1434),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1481),
.B(n_1434),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1480),
.A2(n_1407),
.B(n_1402),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1492),
.B(n_1450),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1481),
.B(n_1434),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1483),
.A2(n_1415),
.B(n_1406),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1474),
.A2(n_1408),
.B1(n_1402),
.B2(n_1439),
.C(n_1462),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1492),
.B(n_1452),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1491),
.B(n_1408),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_1467),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1529),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1541),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1541),
.Y(n_1547)
);

AND2x4_ASAP7_75t_SL g1548 ( 
.A(n_1519),
.B(n_1490),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1471),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1482),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1514),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1486),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1555)
);

NAND2xp67_ASAP7_75t_L g1556 ( 
.A(n_1496),
.B(n_1483),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1536),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1540),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1516),
.B(n_1482),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1521),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1471),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1490),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1525),
.Y(n_1565)
);

NOR2xp67_ASAP7_75t_L g1566 ( 
.A(n_1521),
.B(n_1467),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1526),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1507),
.Y(n_1568)
);

INVxp33_ASAP7_75t_L g1569 ( 
.A(n_1528),
.Y(n_1569)
);

NOR2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1509),
.B(n_1292),
.Y(n_1570)
);

AND2x4_ASAP7_75t_SL g1571 ( 
.A(n_1533),
.B(n_1470),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1471),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1467),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1494),
.B(n_1539),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1506),
.B(n_1505),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1532),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1537),
.B(n_1474),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1520),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1554),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1570),
.A2(n_1515),
.B1(n_1503),
.B2(n_1499),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1576),
.B(n_1522),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1501),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1574),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1575),
.B(n_1511),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1554),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1544),
.B(n_1538),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1574),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1569),
.B(n_1502),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1566),
.Y(n_1593)
);

AOI31xp33_ASAP7_75t_L g1594 ( 
.A1(n_1562),
.A2(n_1499),
.A3(n_1509),
.B(n_1508),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1566),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1545),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1545),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1547),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1548),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1558),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1470),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1562),
.A2(n_1504),
.B(n_1498),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1576),
.A2(n_1535),
.B(n_1504),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1470),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1568),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1547),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1546),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1474),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1558),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1571),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1546),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1546),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1522),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1550),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1550),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1577),
.B(n_1487),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1535),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1594),
.A2(n_1577),
.B(n_1498),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1587),
.B(n_1579),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1551),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1544),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1596),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1591),
.B(n_1579),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1599),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1599),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1593),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1584),
.B(n_1551),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1597),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1581),
.A2(n_1592),
.B1(n_1588),
.B2(n_1603),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1598),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1555),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1557),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1602),
.B(n_1513),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1614),
.B(n_1561),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1607),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1586),
.B(n_1555),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1617),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1639)
);

NOR4xp25_ASAP7_75t_L g1640 ( 
.A(n_1614),
.B(n_1595),
.C(n_1618),
.D(n_1572),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_1563),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1580),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1555),
.Y(n_1643)
);

NAND2x2_ASAP7_75t_L g1644 ( 
.A(n_1611),
.B(n_1341),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1589),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1605),
.B(n_1564),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1582),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_SL g1648 ( 
.A(n_1582),
.B(n_1292),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1608),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1605),
.B(n_1564),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1585),
.B(n_1559),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1616),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1549),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1583),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1601),
.A2(n_1572),
.B(n_1563),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1549),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1601),
.A2(n_1548),
.B(n_1604),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1611),
.B(n_1549),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1601),
.B(n_1571),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1612),
.B(n_1559),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1583),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1601),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1641),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1633),
.B(n_1600),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1630),
.A2(n_1548),
.B1(n_1604),
.B2(n_1510),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1625),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1619),
.A2(n_1563),
.B1(n_1572),
.B2(n_1604),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1646),
.B(n_1604),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1627),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1623),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1626),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1610),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1623),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1610),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1654),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1621),
.B(n_1613),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1631),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1634),
.B(n_1542),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1620),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1648),
.B(n_1331),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1650),
.B(n_1578),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1615),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1622),
.B(n_1578),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1658),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1560),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_SL g1691 ( 
.A(n_1655),
.B(n_1354),
.C(n_1542),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1628),
.B(n_1561),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1628),
.B(n_1550),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1556),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1636),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1622),
.B(n_1573),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1659),
.B(n_1573),
.Y(n_1697)
);

AOI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1670),
.A2(n_1648),
.B(n_1635),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1666),
.A2(n_1644),
.B1(n_1542),
.B2(n_1635),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1689),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1667),
.B(n_1632),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1667),
.B(n_1636),
.Y(n_1703)
);

AOI322xp5_ASAP7_75t_L g1704 ( 
.A1(n_1691),
.A2(n_1643),
.A3(n_1637),
.B1(n_1632),
.B2(n_1658),
.C1(n_1656),
.C2(n_1653),
.Y(n_1704)
);

XOR2x2_ASAP7_75t_L g1705 ( 
.A(n_1683),
.B(n_1512),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1672),
.B(n_1301),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1691),
.A2(n_1644),
.B1(n_1659),
.B2(n_1642),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1672),
.B(n_1645),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1681),
.A2(n_1639),
.B1(n_1638),
.B2(n_1651),
.C(n_1637),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1671),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1671),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1670),
.A2(n_1661),
.B(n_1652),
.C(n_1649),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1673),
.B(n_1659),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_SL g1717 ( 
.A1(n_1673),
.A2(n_1556),
.B(n_1660),
.C(n_1652),
.Y(n_1717)
);

AOI322xp5_ASAP7_75t_L g1718 ( 
.A1(n_1682),
.A2(n_1643),
.A3(n_1656),
.B1(n_1653),
.B2(n_1552),
.C1(n_1543),
.C2(n_1649),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1688),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1682),
.A2(n_1542),
.B(n_1517),
.Y(n_1720)
);

NAND4xp25_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1523),
.C(n_1567),
.D(n_1565),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1684),
.B(n_1560),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1675),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1703),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1715),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1719),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1700),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1708),
.B(n_1662),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1701),
.A2(n_1663),
.B(n_1668),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1707),
.B(n_1684),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1662),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1709),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1722),
.B(n_1664),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1698),
.B(n_1686),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1699),
.A2(n_1694),
.B1(n_1669),
.B2(n_1688),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1710),
.A2(n_1694),
.B1(n_1699),
.B2(n_1720),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1698),
.B(n_1704),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1718),
.B(n_1686),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1688),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1723),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1743),
.B(n_1716),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1732),
.B(n_1301),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1724),
.A2(n_1717),
.B1(n_1720),
.B2(n_1713),
.C(n_1663),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1663),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1738),
.A2(n_1721),
.B(n_1664),
.C(n_1690),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1725),
.B(n_1677),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1737),
.A2(n_1680),
.B(n_1675),
.C(n_1676),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1725),
.B(n_1696),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_L g1752 ( 
.A(n_1733),
.B(n_1680),
.C(n_1676),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_L g1753 ( 
.A(n_1733),
.B(n_1320),
.C(n_1695),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1727),
.B(n_1696),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1736),
.A2(n_1694),
.B1(n_1692),
.B2(n_1669),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1740),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1746),
.A2(n_1735),
.B(n_1732),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1751),
.B(n_1727),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_L g1760 ( 
.A(n_1747),
.B(n_1730),
.C(n_1726),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1756),
.Y(n_1761)
);

OA22x2_ASAP7_75t_L g1762 ( 
.A1(n_1755),
.A2(n_1728),
.B1(n_1754),
.B2(n_1739),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1748),
.B(n_1728),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1750),
.A2(n_1745),
.B(n_1744),
.C(n_1753),
.Y(n_1764)
);

INVxp33_ASAP7_75t_SL g1765 ( 
.A(n_1752),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1746),
.B(n_1734),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1755),
.A2(n_1694),
.B1(n_1730),
.B2(n_1741),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1756),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1765),
.B(n_1740),
.Y(n_1769)
);

O2A1O1Ixp5_ASAP7_75t_SL g1770 ( 
.A1(n_1761),
.A2(n_1726),
.B(n_1729),
.C(n_1742),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1760),
.B(n_1729),
.Y(n_1771)
);

NOR4xp75_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1690),
.C(n_1685),
.D(n_1730),
.Y(n_1772)
);

NOR4xp75_ASAP7_75t_L g1773 ( 
.A(n_1763),
.B(n_1685),
.C(n_1730),
.D(n_1740),
.Y(n_1773)
);

AO221x1_ASAP7_75t_L g1774 ( 
.A1(n_1768),
.A2(n_1742),
.B1(n_1695),
.B2(n_1762),
.C(n_1687),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1771),
.Y(n_1775)
);

NAND2x1_ASAP7_75t_L g1776 ( 
.A(n_1774),
.B(n_1740),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1769),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1773),
.A2(n_1764),
.B(n_1757),
.C(n_1767),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1772),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1770),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1778),
.A2(n_1759),
.B(n_1758),
.C(n_1734),
.Y(n_1781)
);

XNOR2xp5_ASAP7_75t_L g1782 ( 
.A(n_1777),
.B(n_1779),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1775),
.A2(n_1694),
.B1(n_1678),
.B2(n_1687),
.Y(n_1783)
);

XNOR2xp5_ASAP7_75t_L g1784 ( 
.A(n_1776),
.B(n_1390),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1780),
.Y(n_1785)
);

AOI22x1_ASAP7_75t_L g1786 ( 
.A1(n_1784),
.A2(n_1390),
.B1(n_1778),
.B2(n_1327),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1782),
.Y(n_1787)
);

AND3x4_ASAP7_75t_L g1788 ( 
.A(n_1785),
.B(n_1687),
.C(n_1678),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1787),
.A2(n_1783),
.B1(n_1327),
.B2(n_1781),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1788),
.B1(n_1786),
.B2(n_1678),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1790),
.A2(n_1665),
.B1(n_1679),
.B2(n_1692),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1665),
.B1(n_1679),
.B2(n_1693),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1791),
.A2(n_1693),
.B1(n_1697),
.B2(n_1543),
.Y(n_1793)
);

OAI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1792),
.A2(n_1697),
.B(n_1451),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1794),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1793),
.B(n_1296),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1796),
.B(n_1312),
.Y(n_1797)
);

AOI322xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1513),
.A3(n_1517),
.B1(n_1312),
.B2(n_1296),
.C1(n_1573),
.C2(n_1367),
.Y(n_1798)
);

OAI31xp33_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1424),
.A3(n_1367),
.B(n_1374),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1386),
.B(n_1424),
.C(n_1352),
.Y(n_1800)
);


endmodule