module fake_ariane_510_n_30 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_30);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_30;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_27;
wire n_29;
wire n_17;
wire n_18;
wire n_28;
wire n_11;
wire n_26;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_4),
.A2(n_0),
.B1(n_3),
.B2(n_7),
.Y(n_10)
);

A2O1A1Ixp33_ASAP7_75t_L g11 ( 
.A1(n_0),
.A2(n_5),
.B(n_1),
.C(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_3),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

AO31x2_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_2),
.A3(n_6),
.B(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_16),
.B(n_9),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_11),
.B(n_12),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_15),
.B1(n_13),
.B2(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_14),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_16),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_18),
.B(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_25),
.B1(n_14),
.B2(n_21),
.C(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_21),
.B1(n_14),
.B2(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_17),
.B(n_28),
.Y(n_30)
);


endmodule