module fake_jpeg_25439_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_31;
wire n_17;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_SL g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_17),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_34),
.B(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_25),
.B1(n_27),
.B2(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_10),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.C(n_25),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_8),
.C(n_6),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_35),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_38),
.B1(n_40),
.B2(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_31),
.B1(n_15),
.B2(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_44),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_16),
.C(n_13),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_45),
.C(n_16),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_61),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_46),
.A3(n_13),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_1),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_54),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_2),
.B(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_56),
.B1(n_52),
.B2(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_13),
.C(n_4),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_64),
.C(n_65),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_13),
.B1(n_5),
.B2(n_2),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_71),
.B(n_5),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_9),
.B(n_13),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_9),
.Y(n_76)
);


endmodule