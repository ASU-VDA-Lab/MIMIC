module fake_jpeg_15496_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_25),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_28),
.B1(n_33),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_60),
.B1(n_46),
.B2(n_44),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_33),
.B1(n_16),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_62),
.B1(n_42),
.B2(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_33),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_23),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_16),
.B1(n_25),
.B2(n_32),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_75),
.B1(n_99),
.B2(n_100),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_30),
.B1(n_17),
.B2(n_26),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_70),
.B1(n_89),
.B2(n_46),
.Y(n_109)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_42),
.B1(n_44),
.B2(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_73),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_76),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_31),
.B1(n_20),
.B2(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_17),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_23),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_34),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_61),
.B1(n_50),
.B2(n_53),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_44),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_79),
.B1(n_63),
.B2(n_99),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_46),
.C(n_36),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_38),
.C(n_36),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_18),
.A3(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_124),
.B1(n_70),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_18),
.B1(n_27),
.B2(n_21),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_132),
.B(n_67),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_81),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_101),
.B(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_157),
.B1(n_158),
.B2(n_77),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_146),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_148),
.B(n_150),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_78),
.CI(n_91),
.CON(n_143),
.SN(n_143)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_153),
.B1(n_120),
.B2(n_117),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_93),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_90),
.B(n_94),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_108),
.B1(n_133),
.B2(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_72),
.B1(n_95),
.B2(n_119),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_0),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_110),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_27),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_100),
.B1(n_64),
.B2(n_87),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_113),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_19),
.B(n_21),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_127),
.B(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_71),
.B1(n_82),
.B2(n_84),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_107),
.A2(n_133),
.B1(n_116),
.B2(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_104),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_166),
.B1(n_175),
.B2(n_184),
.Y(n_206)
);

HAxp5_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_103),
.CON(n_163),
.SN(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_129),
.B1(n_128),
.B2(n_124),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_125),
.B(n_128),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_170),
.B(n_190),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_103),
.B(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_179),
.C(n_180),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_155),
.B1(n_159),
.B2(n_119),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_148),
.B1(n_143),
.B2(n_160),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_85),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_122),
.C(n_112),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_122),
.C(n_131),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_127),
.B1(n_112),
.B2(n_131),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_19),
.B1(n_21),
.B2(n_38),
.Y(n_214)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_197),
.C(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_196),
.A2(n_161),
.B1(n_190),
.B2(n_199),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_150),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_137),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_210),
.C(n_216),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_134),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_134),
.B(n_1),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_168),
.B(n_186),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_172),
.B1(n_178),
.B2(n_162),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_29),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_177),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_29),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_227),
.B1(n_229),
.B2(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_226),
.B(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_162),
.B1(n_165),
.B2(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_213),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_180),
.C(n_173),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_238),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_173),
.B(n_165),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_166),
.B1(n_176),
.B2(n_19),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_193),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_102),
.C(n_37),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_244),
.C(n_204),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_102),
.C(n_37),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_29),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_3),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_205),
.B1(n_3),
.B2(n_4),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_201),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_241),
.B1(n_222),
.B2(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_222),
.B1(n_204),
.B2(n_205),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_263),
.C(n_265),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_221),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_266),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_197),
.B1(n_203),
.B2(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_249),
.B1(n_264),
.B2(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_2),
.C(n_3),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_3),
.C(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_9),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_245),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_236),
.B1(n_244),
.B2(n_243),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_233),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.C(n_279),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_225),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_232),
.B(n_252),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_283),
.B(n_284),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_231),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_227),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_265),
.C(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_235),
.B(n_247),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_224),
.B(n_246),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_246),
.B1(n_248),
.B2(n_254),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_261),
.B(n_246),
.C(n_263),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_276),
.B1(n_281),
.B2(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_299),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_274),
.B(n_11),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_7),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_287),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_271),
.C(n_275),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_287),
.C(n_294),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_292),
.B1(n_289),
.B2(n_6),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_308),
.B1(n_292),
.B2(n_14),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_279),
.B1(n_272),
.B2(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_290),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_310),
.B(n_296),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_288),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_296),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_318),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_303),
.C(n_292),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_301),
.B(n_289),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_314),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_326),
.A2(n_327),
.B(n_310),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_322),
.B(n_324),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_329),
.CI(n_7),
.CON(n_330),
.SN(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_15),
.B(n_5),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_330),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_330),
.Y(n_333)
);


endmodule