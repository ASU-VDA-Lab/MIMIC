module fake_jpeg_17821_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx5_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_11),
.B1(n_13),
.B2(n_8),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_13),
.B(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_15),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_9),
.B1(n_13),
.B2(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_12),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_31),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_28),
.B(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_46),
.B(n_7),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_38),
.B1(n_10),
.B2(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_0),
.B1(n_2),
.B2(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_43),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_7),
.B(n_21),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_12),
.Y(n_54)
);

OAI31xp33_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_0),
.A3(n_2),
.B(n_12),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_21),
.C(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_18),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_21),
.B(n_17),
.Y(n_57)
);


endmodule