module fake_jpeg_24316_n_71 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_25;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_16),
.B1(n_2),
.B2(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_29),
.B(n_27),
.C(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_44),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_49),
.C(n_46),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_52),
.B(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_23),
.B1(n_30),
.B2(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_51),
.C(n_43),
.Y(n_65)
);

AOI321xp33_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_29),
.A3(n_34),
.B1(n_37),
.B2(n_41),
.C(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_63),
.C(n_22),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_34),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_41),
.B(n_53),
.C(n_48),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_53),
.B(n_48),
.Y(n_71)
);


endmodule