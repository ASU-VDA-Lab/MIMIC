module fake_jpeg_20839_n_162 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_6),
.B(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_63),
.B1(n_67),
.B2(n_15),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_27),
.B1(n_22),
.B2(n_15),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_14),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_77),
.B1(n_87),
.B2(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_14),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_83),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_95),
.B(n_0),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_27),
.B1(n_16),
.B2(n_14),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_27),
.B1(n_19),
.B2(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_27),
.B1(n_1),
.B2(n_3),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_97),
.B1(n_70),
.B2(n_60),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_27),
.B(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_70),
.B(n_45),
.C(n_69),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_6),
.B(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_61),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_108),
.C(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_110),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_97),
.B(n_90),
.C(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_9),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_5),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_112),
.A2(n_81),
.B1(n_75),
.B2(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_81),
.C(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_126),
.C(n_108),
.Y(n_131)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_92),
.CI(n_85),
.CON(n_123),
.SN(n_123)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

OAI211xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_92),
.B(n_93),
.C(n_69),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_5),
.C(n_6),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_99),
.B(n_113),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_135),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_100),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_137),
.C(n_126),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_123),
.C(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_121),
.B1(n_119),
.B2(n_125),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_129),
.B(n_128),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_141),
.B(n_127),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_121),
.B(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_144),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_103),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_123),
.Y(n_145)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_8),
.B(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_139),
.B1(n_143),
.B2(n_147),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_154),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_114),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_153),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_157),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.Y(n_162)
);


endmodule