module fake_jpeg_5954_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.C(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_38),
.CON(n_52),
.SN(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_20),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_25),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_49),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_75),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_28),
.B1(n_22),
.B2(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_46),
.B1(n_60),
.B2(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_27),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_43),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_57),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_65),
.C(n_24),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_57),
.C(n_45),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_65),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.C(n_76),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_47),
.B1(n_55),
.B2(n_48),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_73),
.B1(n_75),
.B2(n_66),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_75),
.B1(n_66),
.B2(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_61),
.B1(n_71),
.B2(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_110),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_58),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_79),
.B(n_25),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_83),
.C(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_24),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_19),
.C(n_23),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_120),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_100),
.B1(n_106),
.B2(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_97),
.Y(n_120)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_79),
.B1(n_85),
.B2(n_94),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_79),
.B(n_30),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_43),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_99),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_98),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_64),
.C(n_15),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_149),
.B1(n_21),
.B2(n_26),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_128),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_115),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_143),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_107),
.B(n_108),
.C(n_100),
.D(n_106),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_16),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_16),
.B1(n_26),
.B2(n_21),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_60),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_58),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_158),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_128),
.C(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_154),
.C(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_39),
.B1(n_35),
.B2(n_16),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_161),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_26),
.C(n_21),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_145),
.B1(n_142),
.B2(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_135),
.B1(n_146),
.B2(n_138),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_157),
.C(n_156),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_151),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_7),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_173),
.B(n_164),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.C(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_9),
.C(n_10),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_194),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_168),
.C(n_7),
.D(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_184),
.C(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_167),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_10),
.C(n_12),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_190),
.B(n_192),
.C(n_14),
.D(n_12),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_13),
.C(n_197),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_199),
.Y(n_201)
);


endmodule