module real_aes_8417_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI222xp33_ASAP7_75t_L g167 ( .A1(n_0), .A2(n_13), .B1(n_39), .B2(n_168), .C1(n_171), .C2(n_176), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_1), .A2(n_228), .B(n_230), .C(n_305), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_2), .A2(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_3), .B(n_266), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_4), .Y(n_141) );
AOI221xp5_ASAP7_75t_L g145 ( .A1(n_5), .A2(n_17), .B1(n_146), .B2(n_150), .C(n_152), .Y(n_145) );
AOI221xp5_ASAP7_75t_L g87 ( .A1(n_6), .A2(n_66), .B1(n_88), .B2(n_106), .C(n_110), .Y(n_87) );
INVx1_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
AND2x6_ASAP7_75t_L g228 ( .A(n_7), .B(n_203), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_7), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g330 ( .A(n_8), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_9), .B(n_239), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_10), .A2(n_54), .B1(n_188), .B2(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_10), .Y(n_189) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_11), .A2(n_30), .B1(n_95), .B2(n_100), .Y(n_103) );
INVx1_ASAP7_75t_L g221 ( .A(n_12), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_14), .A2(n_27), .B1(n_124), .B2(n_131), .C(n_136), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_15), .A2(n_274), .B(n_315), .C(n_317), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_16), .B(n_266), .Y(n_318) );
AO22x2_ASAP7_75t_L g105 ( .A1(n_18), .A2(n_32), .B1(n_95), .B2(n_96), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_19), .B(n_362), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_20), .A2(n_260), .B(n_291), .C(n_294), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_21), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_22), .B(n_239), .Y(n_275) );
OAI22xp5_ASAP7_75t_SL g82 ( .A1(n_23), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_23), .Y(n_85) );
INVx1_ASAP7_75t_L g272 ( .A(n_24), .Y(n_272) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_25), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_26), .Y(n_303) );
INVx1_ASAP7_75t_L g359 ( .A(n_28), .Y(n_359) );
INVx2_ASAP7_75t_L g226 ( .A(n_29), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_31), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g196 ( .A1(n_32), .A2(n_44), .B1(n_55), .B2(n_197), .C(n_198), .Y(n_196) );
INVxp67_ASAP7_75t_L g199 ( .A(n_32), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_33), .A2(n_260), .B(n_261), .C(n_263), .Y(n_259) );
INVxp67_ASAP7_75t_L g360 ( .A(n_34), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g257 ( .A(n_35), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_36), .A2(n_230), .B(n_271), .C(n_278), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_37), .A2(n_241), .B(n_328), .C(n_329), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_38), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_40), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_41), .Y(n_356) );
INVx1_ASAP7_75t_L g289 ( .A(n_42), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_43), .Y(n_159) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_44), .A2(n_67), .B1(n_95), .B2(n_96), .Y(n_94) );
INVxp67_ASAP7_75t_L g200 ( .A(n_44), .Y(n_200) );
CKINVDCx14_ASAP7_75t_R g326 ( .A(n_45), .Y(n_326) );
INVx1_ASAP7_75t_L g203 ( .A(n_46), .Y(n_203) );
INVx1_ASAP7_75t_L g220 ( .A(n_47), .Y(n_220) );
INVx1_ASAP7_75t_SL g262 ( .A(n_48), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_49), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_50), .B(n_266), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_51), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_52), .A2(n_75), .B1(n_185), .B2(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_52), .Y(n_186) );
INVx1_ASAP7_75t_L g234 ( .A(n_53), .Y(n_234) );
INVx1_ASAP7_75t_L g188 ( .A(n_54), .Y(n_188) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_55), .A2(n_72), .B1(n_95), .B2(n_100), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_56), .A2(n_182), .B1(n_191), .B2(n_192), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g191 ( .A(n_56), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_57), .A2(n_255), .B(n_325), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_58), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_59), .Y(n_246) );
INVx1_ASAP7_75t_L g84 ( .A(n_60), .Y(n_84) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_60), .A2(n_255), .B(n_312), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_61), .A2(n_354), .B(n_355), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_62), .Y(n_269) );
AOI22xp5_ASAP7_75t_SL g531 ( .A1(n_62), .A2(n_86), .B1(n_180), .B2(n_269), .Y(n_531) );
INVx1_ASAP7_75t_L g313 ( .A(n_63), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_64), .A2(n_255), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g316 ( .A(n_65), .Y(n_316) );
INVx2_ASAP7_75t_L g218 ( .A(n_68), .Y(n_218) );
INVx1_ASAP7_75t_L g306 ( .A(n_69), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_70), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_71), .A2(n_230), .B(n_233), .C(n_243), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_73), .B(n_216), .Y(n_331) );
INVx1_ASAP7_75t_L g95 ( .A(n_74), .Y(n_95) );
INVx1_ASAP7_75t_L g97 ( .A(n_74), .Y(n_97) );
INVx1_ASAP7_75t_L g185 ( .A(n_75), .Y(n_185) );
INVx2_ASAP7_75t_L g292 ( .A(n_76), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_77), .A2(n_86), .B1(n_180), .B2(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_77), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_193), .B1(n_206), .B2(n_526), .C(n_530), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_181), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_86), .B2(n_180), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_84), .Y(n_83) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_85), .A2(n_223), .B(n_229), .Y(n_222) );
INVx1_ASAP7_75t_L g180 ( .A(n_86), .Y(n_180) );
AND4x1_ASAP7_75t_L g86 ( .A(n_87), .B(n_123), .C(n_145), .D(n_167), .Y(n_86) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx3_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_101), .Y(n_91) );
AND2x6_ASAP7_75t_L g128 ( .A(n_92), .B(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g140 ( .A(n_92), .B(n_114), .Y(n_140) );
AND2x6_ASAP7_75t_L g170 ( .A(n_92), .B(n_164), .Y(n_170) );
AND2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_98), .Y(n_92) );
AND2x2_ASAP7_75t_L g135 ( .A(n_93), .B(n_99), .Y(n_135) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_94), .B(n_99), .Y(n_109) );
AND2x2_ASAP7_75t_L g115 ( .A(n_94), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g157 ( .A(n_94), .B(n_103), .Y(n_157) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g100 ( .A(n_97), .Y(n_100) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
INVx1_ASAP7_75t_L g175 ( .A(n_99), .Y(n_175) );
AND2x4_ASAP7_75t_L g107 ( .A(n_101), .B(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g134 ( .A(n_101), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_101), .B(n_115), .Y(n_144) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
AND2x2_ASAP7_75t_L g114 ( .A(n_102), .B(n_105), .Y(n_114) );
OR2x2_ASAP7_75t_L g130 ( .A(n_102), .B(n_105), .Y(n_130) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g164 ( .A(n_103), .B(n_105), .Y(n_164) );
INVx1_ASAP7_75t_L g158 ( .A(n_104), .Y(n_158) );
AND2x2_ASAP7_75t_L g174 ( .A(n_104), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x6_ASAP7_75t_L g121 ( .A(n_109), .B(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B1(n_117), .B2(n_118), .Y(n_110) );
BUFx2_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x6_ASAP7_75t_L g151 ( .A(n_114), .B(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx6_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx11_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g149 ( .A(n_129), .B(n_135), .Y(n_149) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_141), .B2(n_142), .Y(n_136) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx4f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_159), .B2(n_160), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2x1p5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x4_ASAP7_75t_L g173 ( .A(n_157), .B(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g178 ( .A(n_157), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_162), .Y(n_161) );
OR2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_165), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g179 ( .A(n_175), .Y(n_179) );
BUFx4f_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
BUFx12f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_182), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_187), .B2(n_190), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g190 ( .A(n_187), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
AND3x1_ASAP7_75t_SL g195 ( .A(n_196), .B(n_201), .C(n_204), .Y(n_195) );
INVxp67_ASAP7_75t_L g535 ( .A(n_196), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_SL g537 ( .A(n_201), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_201), .A2(n_528), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g546 ( .A(n_201), .Y(n_546) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_202), .B(n_205), .Y(n_540) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_SL g545 ( .A(n_204), .B(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_208), .B(n_481), .Y(n_207) );
NOR4xp25_ASAP7_75t_L g208 ( .A(n_209), .B(n_418), .C(n_452), .D(n_468), .Y(n_208) );
NAND4xp25_ASAP7_75t_SL g209 ( .A(n_210), .B(n_344), .C(n_382), .D(n_398), .Y(n_209) );
AOI222xp33_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_281), .B1(n_319), .B2(n_332), .C1(n_337), .C2(n_343), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI31xp33_ASAP7_75t_L g514 ( .A1(n_212), .A2(n_515), .A3(n_516), .B(n_518), .Y(n_514) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_249), .Y(n_212) );
AND2x2_ASAP7_75t_L g489 ( .A(n_213), .B(n_251), .Y(n_489) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_SL g336 ( .A(n_214), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_214), .B(n_267), .Y(n_343) );
AND2x2_ASAP7_75t_L g403 ( .A(n_214), .B(n_252), .Y(n_403) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_222), .B(n_245), .Y(n_214) );
INVx3_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_215), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_215), .B(n_309), .Y(n_308) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g352 ( .A(n_217), .Y(n_352) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x2_ASAP7_75t_SL g248 ( .A(n_218), .B(n_219), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_223), .A2(n_248), .B(n_269), .C(n_270), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_223), .A2(n_303), .B(n_304), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
AND2x4_ASAP7_75t_L g255 ( .A(n_224), .B(n_228), .Y(n_255) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g231 ( .A(n_226), .Y(n_231) );
INVx1_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
INVx1_ASAP7_75t_L g232 ( .A(n_227), .Y(n_232) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_227), .Y(n_237) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
INVx3_ASAP7_75t_L g274 ( .A(n_227), .Y(n_274) );
INVx4_ASAP7_75t_SL g244 ( .A(n_228), .Y(n_244) );
BUFx3_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
INVx5_ASAP7_75t_L g258 ( .A(n_230), .Y(n_258) );
AND2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
BUFx3_ASAP7_75t_L g242 ( .A(n_231), .Y(n_242) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_238), .C(n_240), .Y(n_233) );
O2A1O1Ixp5_ASAP7_75t_L g305 ( .A1(n_235), .A2(n_240), .B(n_306), .C(n_307), .Y(n_305) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_235), .Y(n_529) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx4_ASAP7_75t_L g293 ( .A(n_237), .Y(n_293) );
INVx4_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
INVx2_ASAP7_75t_L g328 ( .A(n_239), .Y(n_328) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g317 ( .A(n_242), .Y(n_317) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_244), .A2(n_257), .B(n_258), .C(n_259), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g288 ( .A1(n_244), .A2(n_258), .B(n_289), .C(n_290), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_SL g312 ( .A1(n_244), .A2(n_258), .B(n_313), .C(n_314), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_SL g325 ( .A1(n_244), .A2(n_258), .B(n_326), .C(n_327), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g355 ( .A1(n_244), .A2(n_258), .B(n_356), .C(n_357), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g362 ( .A(n_247), .Y(n_362) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g301 ( .A(n_248), .Y(n_301) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_248), .A2(n_324), .B(n_331), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_249), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_250), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_250), .B(n_347), .Y(n_393) );
AND2x2_ASAP7_75t_L g486 ( .A(n_250), .B(n_426), .Y(n_486) );
OAI321xp33_ASAP7_75t_L g520 ( .A1(n_250), .A2(n_336), .A3(n_493), .B1(n_521), .B2(n_523), .C(n_524), .Y(n_520) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_250), .B(n_322), .C(n_433), .D(n_525), .Y(n_524) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_267), .Y(n_250) );
AND2x2_ASAP7_75t_L g388 ( .A(n_251), .B(n_334), .Y(n_388) );
AND2x2_ASAP7_75t_L g407 ( .A(n_251), .B(n_336), .Y(n_407) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g335 ( .A(n_252), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g363 ( .A(n_252), .B(n_267), .Y(n_363) );
AND2x2_ASAP7_75t_L g449 ( .A(n_252), .B(n_334), .Y(n_449) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_265), .Y(n_252) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_253), .A2(n_287), .B(n_296), .Y(n_286) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_253), .A2(n_311), .B(n_318), .Y(n_310) );
BUFx2_ASAP7_75t_L g354 ( .A(n_255), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_260), .B(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_SL g334 ( .A(n_267), .Y(n_334) );
AND2x2_ASAP7_75t_L g381 ( .A(n_267), .B(n_368), .Y(n_381) );
OR2x2_ASAP7_75t_L g414 ( .A(n_267), .B(n_336), .Y(n_414) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_267), .Y(n_421) );
AND2x2_ASAP7_75t_L g450 ( .A(n_267), .B(n_335), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_267), .B(n_423), .Y(n_465) );
AND2x2_ASAP7_75t_L g497 ( .A(n_267), .B(n_489), .Y(n_497) );
AND2x2_ASAP7_75t_L g506 ( .A(n_267), .B(n_348), .Y(n_506) );
OR2x6_ASAP7_75t_L g267 ( .A(n_268), .B(n_279), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B(n_275), .C(n_276), .Y(n_271) );
OAI322xp33_ASAP7_75t_L g530 ( .A1(n_272), .A2(n_531), .A3(n_532), .B1(n_536), .B2(n_538), .C1(n_541), .C2(n_543), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_273), .A2(n_293), .B1(n_359), .B2(n_360), .Y(n_358) );
INVx5_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_274), .B(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_276), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_277), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_278), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_297), .Y(n_282) );
INVx1_ASAP7_75t_SL g474 ( .A(n_283), .Y(n_474) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g339 ( .A(n_284), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g321 ( .A(n_285), .B(n_299), .Y(n_321) );
AND2x2_ASAP7_75t_L g410 ( .A(n_285), .B(n_323), .Y(n_410) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g380 ( .A(n_286), .B(n_310), .Y(n_380) );
OR2x2_ASAP7_75t_L g391 ( .A(n_286), .B(n_323), .Y(n_391) );
AND2x2_ASAP7_75t_L g417 ( .A(n_286), .B(n_323), .Y(n_417) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_286), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_293), .B(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_297), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_297), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g390 ( .A(n_298), .B(n_391), .Y(n_390) );
AOI322xp5_ASAP7_75t_L g476 ( .A1(n_298), .A2(n_380), .A3(n_386), .B1(n_417), .B2(n_467), .C1(n_477), .C2(n_479), .Y(n_476) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_310), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_322), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_299), .B(n_323), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_299), .B(n_340), .Y(n_397) );
AND2x2_ASAP7_75t_L g451 ( .A(n_299), .B(n_417), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_299), .Y(n_455) );
AND2x2_ASAP7_75t_L g467 ( .A(n_299), .B(n_310), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_299), .B(n_339), .Y(n_499) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g364 ( .A(n_300), .B(n_310), .Y(n_364) );
BUFx3_ASAP7_75t_L g378 ( .A(n_300), .Y(n_378) );
AND3x2_ASAP7_75t_L g460 ( .A(n_300), .B(n_440), .C(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_308), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_310), .B(n_321), .C(n_322), .Y(n_320) );
INVx1_ASAP7_75t_SL g340 ( .A(n_310), .Y(n_340) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_310), .Y(n_445) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g439 ( .A(n_321), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g446 ( .A(n_321), .Y(n_446) );
AND2x2_ASAP7_75t_L g484 ( .A(n_322), .B(n_462), .Y(n_484) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
AND2x2_ASAP7_75t_L g440 ( .A(n_323), .B(n_340), .Y(n_440) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g384 ( .A(n_334), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g503 ( .A(n_334), .B(n_403), .Y(n_503) );
AND2x2_ASAP7_75t_L g517 ( .A(n_334), .B(n_336), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_335), .B(n_348), .Y(n_458) );
AND2x2_ASAP7_75t_L g505 ( .A(n_335), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g368 ( .A(n_336), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g385 ( .A(n_336), .B(n_348), .Y(n_385) );
INVx1_ASAP7_75t_L g395 ( .A(n_336), .Y(n_395) );
AND2x2_ASAP7_75t_L g426 ( .A(n_336), .B(n_348), .Y(n_426) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_338), .A2(n_469), .B1(n_473), .B2(n_475), .C(n_476), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g372 ( .A(n_339), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_342), .B(n_379), .Y(n_522) );
AOI322xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_364), .A3(n_365), .B1(n_366), .B2(n_372), .C1(n_374), .C2(n_381), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_363), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_347), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_347), .B(n_413), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_347), .A2(n_363), .B(n_437), .C(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_347), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_347), .B(n_407), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_347), .B(n_489), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_347), .B(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_348), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_348), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g478 ( .A(n_348), .B(n_365), .Y(n_478) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B(n_361), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_350), .A2(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g370 ( .A(n_353), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_361), .Y(n_371) );
INVx1_ASAP7_75t_L g453 ( .A(n_363), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g463 ( .A1(n_363), .A2(n_388), .A3(n_464), .B(n_466), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_363), .B(n_369), .Y(n_515) );
INVx1_ASAP7_75t_SL g376 ( .A(n_364), .Y(n_376) );
AND2x2_ASAP7_75t_L g409 ( .A(n_364), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g490 ( .A(n_364), .B(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g375 ( .A(n_365), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g400 ( .A(n_365), .Y(n_400) );
AND2x2_ASAP7_75t_L g427 ( .A(n_365), .B(n_380), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_365), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g519 ( .A(n_365), .B(n_467), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_367), .B(n_437), .Y(n_510) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g406 ( .A(n_369), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g424 ( .A(n_369), .Y(n_424) );
NAND2xp33_ASAP7_75t_SL g374 ( .A(n_375), .B(n_377), .Y(n_374) );
OAI211xp5_ASAP7_75t_SL g418 ( .A1(n_376), .A2(n_419), .B(n_425), .C(n_441), .Y(n_418) );
OR2x2_ASAP7_75t_L g493 ( .A(n_376), .B(n_474), .Y(n_493) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_378), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_378), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g399 ( .A(n_380), .B(n_400), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B(n_389), .C(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g433 ( .A(n_385), .Y(n_433) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_388), .B(n_426), .Y(n_431) );
INVx1_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g396 ( .A(n_391), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g429 ( .A(n_391), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g491 ( .A(n_391), .Y(n_491) );
AOI21xp33_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B(n_396), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_394), .A2(n_405), .B(n_408), .Y(n_404) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_404), .C(n_411), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_399), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_402), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g415 ( .A(n_403), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_405), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_410), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g435 ( .A(n_410), .Y(n_435) );
AOI21xp33_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_415), .B(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g466 ( .A(n_417), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_423), .B(n_449), .Y(n_475) );
AND2x2_ASAP7_75t_L g488 ( .A(n_423), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g502 ( .A(n_423), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g512 ( .A(n_423), .B(n_450), .Y(n_512) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_428), .C(n_436), .Y(n_425) );
INVx1_ASAP7_75t_L g472 ( .A(n_426), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_432), .B2(n_434), .Y(n_428) );
OR2x2_ASAP7_75t_L g434 ( .A(n_430), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_430), .B(n_491), .Y(n_513) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_447), .B1(n_450), .B2(n_451), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g471 ( .A(n_449), .Y(n_471) );
OAI211xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B(n_456), .C(n_463), .Y(n_452) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_471), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR5xp2_ASAP7_75t_L g481 ( .A(n_482), .B(n_500), .C(n_508), .D(n_514), .E(n_520), .Y(n_481) );
OAI211xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_485), .B(n_487), .C(n_494), .Y(n_482) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_492), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_497), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_SL g523 ( .A(n_503), .Y(n_523) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_511), .B(n_513), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
endmodule