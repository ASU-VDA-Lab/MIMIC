module real_aes_2001_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_786, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_786;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g532 ( .A(n_0), .B(n_158), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_1), .B(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_2), .B(n_140), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_3), .B(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g147 ( .A(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_5), .B(n_140), .Y(n_488) );
NAND2xp33_ASAP7_75t_SL g524 ( .A(n_6), .B(n_146), .Y(n_524) );
INVx1_ASAP7_75t_L g517 ( .A(n_7), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g781 ( .A(n_9), .Y(n_781) );
AND2x2_ASAP7_75t_L g486 ( .A(n_10), .B(n_171), .Y(n_486) );
AND2x2_ASAP7_75t_L g205 ( .A(n_11), .B(n_190), .Y(n_205) );
AND2x2_ASAP7_75t_L g213 ( .A(n_12), .B(n_134), .Y(n_213) );
INVx2_ASAP7_75t_L g137 ( .A(n_13), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_14), .B(n_156), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_16), .A2(n_134), .B1(n_149), .B2(n_521), .C(n_523), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_17), .B(n_140), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_18), .B(n_140), .Y(n_184) );
INVx1_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_20), .A2(n_87), .B1(n_140), .B2(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_21), .A2(n_149), .B(n_490), .Y(n_489) );
AOI221xp5_ASAP7_75t_SL g499 ( .A1(n_22), .A2(n_37), .B1(n_140), .B2(n_149), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_23), .B(n_158), .Y(n_491) );
INVxp33_ASAP7_75t_L g783 ( .A(n_24), .Y(n_783) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_25), .A2(n_86), .B(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g161 ( .A(n_25), .B(n_86), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_26), .B(n_156), .Y(n_511) );
INVxp67_ASAP7_75t_L g519 ( .A(n_27), .Y(n_519) );
AND2x2_ASAP7_75t_L g548 ( .A(n_28), .B(n_175), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_29), .A2(n_149), .B(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_30), .A2(n_134), .B(n_138), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_31), .B(n_156), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_32), .A2(n_149), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_33), .B(n_156), .Y(n_168) );
AND2x2_ASAP7_75t_L g146 ( .A(n_34), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g150 ( .A(n_34), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g229 ( .A(n_34), .Y(n_229) );
OR2x6_ASAP7_75t_L g113 ( .A(n_35), .B(n_114), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_35), .B(n_111), .C(n_780), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_36), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_38), .B(n_140), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_39), .A2(n_79), .B1(n_149), .B2(n_227), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_40), .B(n_156), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_41), .B(n_140), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_42), .B(n_158), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_43), .A2(n_149), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_44), .B(n_158), .Y(n_252) );
AND2x2_ASAP7_75t_L g535 ( .A(n_45), .B(n_175), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_46), .B(n_175), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_47), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g143 ( .A(n_48), .Y(n_143) );
INVx1_ASAP7_75t_L g153 ( .A(n_48), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_49), .B(n_156), .Y(n_211) );
AND2x2_ASAP7_75t_L g174 ( .A(n_50), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_51), .B(n_140), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_52), .B(n_158), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_53), .B(n_158), .Y(n_167) );
AND2x2_ASAP7_75t_L g482 ( .A(n_54), .B(n_175), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_55), .B(n_140), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_56), .B(n_156), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_57), .B(n_140), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_58), .A2(n_149), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_59), .B(n_158), .Y(n_480) );
AND2x2_ASAP7_75t_SL g512 ( .A(n_60), .B(n_171), .Y(n_512) );
AND2x2_ASAP7_75t_L g191 ( .A(n_61), .B(n_171), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_62), .A2(n_149), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_63), .B(n_156), .Y(n_492) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_64), .B(n_190), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_65), .B(n_158), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_66), .B(n_158), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_67), .A2(n_90), .B1(n_149), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_68), .B(n_156), .Y(n_187) );
INVx1_ASAP7_75t_L g145 ( .A(n_69), .Y(n_145) );
INVx1_ASAP7_75t_L g151 ( .A(n_69), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_70), .B(n_158), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_71), .A2(n_149), .B(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_72), .A2(n_149), .B(n_250), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_73), .A2(n_149), .B(n_154), .Y(n_148) );
AND2x2_ASAP7_75t_L g170 ( .A(n_74), .B(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_75), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_75), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_76), .B(n_175), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_77), .B(n_140), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_78), .A2(n_81), .B1(n_140), .B2(n_221), .Y(n_583) );
INVx1_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_80), .B(n_115), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_82), .B(n_158), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_83), .B(n_158), .Y(n_502) );
AND2x2_ASAP7_75t_L g253 ( .A(n_84), .B(n_190), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_85), .A2(n_149), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_88), .B(n_156), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_89), .A2(n_149), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_91), .B(n_156), .Y(n_251) );
BUFx2_ASAP7_75t_L g189 ( .A(n_92), .Y(n_189) );
INVxp67_ASAP7_75t_L g522 ( .A(n_93), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_94), .B(n_140), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_95), .A2(n_149), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_96), .B(n_156), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_97), .A2(n_119), .B1(n_758), .B2(n_760), .Y(n_757) );
BUFx2_ASAP7_75t_L g105 ( .A(n_98), .Y(n_105) );
BUFx2_ASAP7_75t_SL g764 ( .A(n_98), .Y(n_764) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_773), .B(n_782), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_118), .B(n_762), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_107), .A2(n_766), .B(n_770), .Y(n_765) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_117), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g772 ( .A(n_110), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x6_ASAP7_75t_SL g125 ( .A(n_111), .B(n_112), .Y(n_125) );
AND2x6_ASAP7_75t_SL g466 ( .A(n_111), .B(n_113), .Y(n_466) );
OR2x2_ASAP7_75t_L g761 ( .A(n_111), .B(n_113), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B(n_757), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_126), .B(n_463), .Y(n_121) );
BUFx4f_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
CKINVDCx11_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_125), .A2(n_127), .B1(n_467), .B2(n_759), .Y(n_758) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND3x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_341), .C(n_437), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_283), .C(n_310), .Y(n_128) );
OAI211xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_192), .B(n_232), .C(n_256), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_172), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_131), .A2(n_234), .B(n_238), .C(n_244), .Y(n_233) );
OR2x2_ASAP7_75t_L g356 ( .A(n_131), .B(n_293), .Y(n_356) );
INVx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g323 ( .A(n_132), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_132), .B(n_294), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_132), .B(n_439), .Y(n_454) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_162), .Y(n_132) );
AND2x2_ASAP7_75t_L g240 ( .A(n_133), .B(n_173), .Y(n_240) );
INVx1_ASAP7_75t_L g260 ( .A(n_133), .Y(n_260) );
OR2x2_ASAP7_75t_L g275 ( .A(n_133), .B(n_182), .Y(n_275) );
INVx2_ASAP7_75t_L g281 ( .A(n_133), .Y(n_281) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_133), .Y(n_336) );
INVx1_ASAP7_75t_L g413 ( .A(n_133), .Y(n_413) );
INVx3_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_135), .A2(n_207), .B(n_213), .Y(n_206) );
AOI21x1_ASAP7_75t_L g528 ( .A1(n_135), .A2(n_529), .B(n_535), .Y(n_528) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx4f_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
AND2x4_ASAP7_75t_L g160 ( .A(n_137), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_137), .B(n_161), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_148), .B(n_160), .Y(n_138) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g525 ( .A(n_141), .Y(n_525) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
AND2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g156 ( .A(n_144), .B(n_153), .Y(n_156) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
AND2x2_ASAP7_75t_L g152 ( .A(n_147), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
BUFx3_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
INVx2_ASAP7_75t_L g231 ( .A(n_151), .Y(n_231) );
AND2x4_ASAP7_75t_L g227 ( .A(n_152), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g223 ( .A(n_153), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_158), .B(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_159), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_159), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_159), .A2(n_251), .B(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_159), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_159), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_159), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_159), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_159), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_159), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_160), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_160), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_160), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_160), .B(n_522), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_160), .B(n_524), .C(n_525), .Y(n_523) );
NOR2x1_ASAP7_75t_SL g262 ( .A(n_162), .B(n_182), .Y(n_262) );
AND2x2_ASAP7_75t_L g292 ( .A(n_162), .B(n_281), .Y(n_292) );
AO21x1_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B(n_170), .Y(n_162) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_163), .A2(n_164), .B(n_170), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_169), .Y(n_164) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_171), .Y(n_175) );
OR2x2_ASAP7_75t_L g286 ( .A(n_172), .B(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_172), .B(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g414 ( .A(n_172), .Y(n_414) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_173), .B(n_182), .Y(n_172) );
OR2x2_ASAP7_75t_SL g274 ( .A(n_173), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
INVx4_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
OR2x2_ASAP7_75t_L g309 ( .A(n_173), .B(n_242), .Y(n_309) );
AND2x2_ASAP7_75t_L g348 ( .A(n_173), .B(n_262), .Y(n_348) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_173), .Y(n_360) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_176), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_175), .Y(n_198) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_175), .A2(n_220), .B(n_226), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_175), .A2(n_248), .B(n_249), .Y(n_247) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_175), .A2(n_499), .B(n_503), .Y(n_498) );
AND2x2_ASAP7_75t_L g241 ( .A(n_182), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g293 ( .A(n_182), .B(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g308 ( .A(n_182), .Y(n_308) );
AND2x2_ASAP7_75t_L g324 ( .A(n_182), .B(n_294), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_182), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g369 ( .A(n_182), .B(n_281), .Y(n_369) );
INVx2_ASAP7_75t_SL g439 ( .A(n_182), .Y(n_439) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_191), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_190), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_190), .A2(n_507), .B(n_508), .Y(n_506) );
INVx2_ASAP7_75t_SL g581 ( .A(n_190), .Y(n_581) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp67_ASAP7_75t_L g193 ( .A(n_194), .B(n_214), .Y(n_193) );
OAI211xp5_ASAP7_75t_L g310 ( .A1(n_194), .A2(n_311), .B(n_315), .C(n_331), .Y(n_310) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g406 ( .A(n_195), .B(n_245), .Y(n_406) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
INVx2_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
AND2x4_ASAP7_75t_SL g266 ( .A(n_196), .B(n_246), .Y(n_266) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
AND2x2_ASAP7_75t_L g328 ( .A(n_196), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g402 ( .A(n_196), .Y(n_402) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_197), .Y(n_304) );
AND2x2_ASAP7_75t_L g347 ( .A(n_197), .B(n_206), .Y(n_347) );
AOI21x1_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_205), .Y(n_197) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_198), .A2(n_476), .B(n_482), .Y(n_475) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_198), .A2(n_542), .B(n_548), .Y(n_541) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_198), .A2(n_542), .B(n_548), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_204), .Y(n_199) );
INVx2_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
AND2x2_ASAP7_75t_L g297 ( .A(n_206), .B(n_246), .Y(n_297) );
INVx2_ASAP7_75t_L g329 ( .A(n_206), .Y(n_329) );
OR2x2_ASAP7_75t_L g352 ( .A(n_206), .B(n_217), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_214), .B(n_269), .Y(n_376) );
AND2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_346), .Y(n_410) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OAI31xp33_ASAP7_75t_SL g331 ( .A1(n_215), .A2(n_312), .A3(n_332), .B(n_339), .Y(n_331) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_216), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx3_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
AND2x2_ASAP7_75t_L g282 ( .A(n_217), .B(n_245), .Y(n_282) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x4_ASAP7_75t_L g272 ( .A(n_218), .B(n_219), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_221), .A2(n_227), .B1(n_516), .B2(n_518), .Y(n_515) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_225), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2x1p5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g417 ( .A(n_235), .Y(n_417) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_237), .B(n_246), .Y(n_299) );
AND2x2_ASAP7_75t_L g340 ( .A(n_237), .B(n_255), .Y(n_340) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g320 ( .A(n_241), .B(n_278), .Y(n_320) );
AND2x2_ASAP7_75t_L g279 ( .A(n_242), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
INVx2_ASAP7_75t_L g338 ( .A(n_242), .Y(n_338) );
AND2x2_ASAP7_75t_L g428 ( .A(n_242), .B(n_413), .Y(n_428) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g434 ( .A(n_244), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_245), .B(n_304), .Y(n_373) );
AND2x2_ASAP7_75t_L g421 ( .A(n_245), .B(n_347), .Y(n_421) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g330 ( .A(n_246), .B(n_302), .Y(n_330) );
AND2x2_ASAP7_75t_L g339 ( .A(n_246), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g351 ( .A(n_246), .Y(n_351) );
BUFx2_ASAP7_75t_L g367 ( .A(n_246), .Y(n_367) );
AND2x4_ASAP7_75t_L g401 ( .A(n_246), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g446 ( .A(n_246), .B(n_347), .Y(n_446) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_253), .Y(n_246) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AOI222xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_263), .B1(n_267), .B2(n_273), .C1(n_276), .C2(n_282), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_258), .A2(n_322), .B1(n_325), .B2(n_330), .Y(n_321) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g305 ( .A(n_259), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_SL g319 ( .A(n_259), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_259), .B(n_324), .Y(n_457) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g418 ( .A(n_260), .B(n_324), .Y(n_418) );
OR2x2_ASAP7_75t_L g395 ( .A(n_261), .B(n_277), .Y(n_395) );
OR2x2_ASAP7_75t_L g403 ( .A(n_261), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g387 ( .A(n_262), .B(n_280), .Y(n_387) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g295 ( .A(n_265), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g445 ( .A(n_265), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g396 ( .A(n_266), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_266), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_SL g431 ( .A(n_266), .Y(n_431) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx2_ASAP7_75t_L g416 ( .A(n_269), .Y(n_416) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_297), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_271), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g317 ( .A(n_271), .Y(n_317) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_271), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g420 ( .A(n_271), .B(n_292), .Y(n_420) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g354 ( .A(n_272), .B(n_340), .Y(n_354) );
AND2x2_ASAP7_75t_L g397 ( .A(n_272), .B(n_329), .Y(n_397) );
AND2x4_ASAP7_75t_L g312 ( .A(n_273), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g453 ( .A(n_275), .B(n_309), .Y(n_453) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_277), .B(n_292), .Y(n_436) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_278), .B(n_292), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_278), .A2(n_319), .B(n_420), .C(n_421), .Y(n_419) );
AND2x2_ASAP7_75t_L g450 ( .A(n_278), .B(n_428), .Y(n_450) );
INVx1_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_282), .B(n_346), .Y(n_345) );
OAI21xp33_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_295), .B(n_298), .Y(n_283) );
NOR2x1_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_286), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_294), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g386 ( .A(n_294), .Y(n_386) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_305), .Y(n_298) );
INVx1_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_321), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OR2x2_ASAP7_75t_L g362 ( .A(n_317), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g399 ( .A(n_317), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_317), .B(n_347), .Y(n_435) );
INVx1_ASAP7_75t_L g455 ( .A(n_318), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_320), .A2(n_423), .B1(n_426), .B2(n_429), .C(n_432), .Y(n_422) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI321xp33_ASAP7_75t_L g443 ( .A1(n_325), .A2(n_360), .A3(n_444), .B1(n_447), .B2(n_449), .C(n_451), .Y(n_443) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_337), .A2(n_365), .B1(n_369), .B2(n_370), .C(n_375), .Y(n_364) );
INVxp67_ASAP7_75t_L g393 ( .A(n_338), .Y(n_393) );
INVx1_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
NOR2xp67_ASAP7_75t_L g341 ( .A(n_342), .B(n_388), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_364), .C(n_379), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_349), .B2(n_355), .C(n_357), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g462 ( .A(n_347), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_353), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_351), .B(n_397), .Y(n_442) );
INVx2_ASAP7_75t_SL g374 ( .A(n_352), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_353), .A2(n_358), .B1(n_359), .B2(n_362), .Y(n_357) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_361), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_362), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g368 ( .A(n_363), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g407 ( .A1(n_365), .A2(n_408), .B1(n_410), .B2(n_411), .C1(n_415), .C2(n_418), .Y(n_407) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_366), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g441 ( .A(n_366), .B(n_420), .Y(n_441) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_374), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_374), .B(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_378), .Y(n_375) );
NAND2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_385), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_385), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND4xp25_ASAP7_75t_SL g388 ( .A(n_389), .B(n_407), .C(n_419), .D(n_422), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_394), .B(n_396), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_395), .A2(n_399), .B1(n_403), .B2(n_405), .Y(n_398) );
INVx1_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_414), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_431), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_436), .Y(n_432) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_443), .C(n_456), .D(n_458), .Y(n_437) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
CKINVDCx11_ASAP7_75t_R g759 ( .A(n_466), .Y(n_759) );
INVx4_ASAP7_75t_L g768 ( .A(n_467), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_467), .Y(n_769) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_696), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_589), .C(n_640), .Y(n_468) );
OAI211xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_493), .B(n_536), .C(n_567), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_483), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_474), .B(n_541), .Y(n_704) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g549 ( .A(n_475), .B(n_485), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_475), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g566 ( .A(n_475), .B(n_556), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_475), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_475), .B(n_579), .Y(n_603) );
INVx2_ASAP7_75t_L g629 ( .A(n_475), .Y(n_629) );
AND2x4_ASAP7_75t_L g638 ( .A(n_475), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g743 ( .A(n_475), .B(n_610), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
AND2x2_ASAP7_75t_L g627 ( .A(n_483), .B(n_628), .Y(n_627) );
OAI32xp33_ASAP7_75t_L g710 ( .A1(n_483), .A2(n_632), .A3(n_636), .B1(n_643), .B2(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_483), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g564 ( .A(n_484), .B(n_565), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_484), .B(n_559), .C(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g663 ( .A(n_484), .B(n_566), .Y(n_663) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
INVx5_ASAP7_75t_L g588 ( .A(n_485), .Y(n_588) );
AND2x4_ASAP7_75t_L g644 ( .A(n_485), .B(n_556), .Y(n_644) );
OR2x2_ASAP7_75t_L g659 ( .A(n_485), .B(n_579), .Y(n_659) );
OR2x2_ASAP7_75t_L g685 ( .A(n_485), .B(n_541), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_485), .B(n_639), .Y(n_693) );
AND2x4_ASAP7_75t_SL g718 ( .A(n_485), .B(n_638), .Y(n_718) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_494), .B(n_638), .Y(n_714) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_495), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x6_ASAP7_75t_SL g538 ( .A(n_496), .B(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g563 ( .A(n_497), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_497), .B(n_598), .Y(n_616) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_497), .Y(n_754) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AND2x2_ASAP7_75t_L g596 ( .A(n_498), .B(n_527), .Y(n_596) );
INVx2_ASAP7_75t_L g624 ( .A(n_498), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_498), .B(n_505), .Y(n_665) );
BUFx3_ASAP7_75t_L g689 ( .A(n_498), .Y(n_689) );
OR2x2_ASAP7_75t_L g701 ( .A(n_498), .B(n_505), .Y(n_701) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_498), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_504), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_731) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx1_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
OR2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g577 ( .A(n_505), .Y(n_577) );
AND2x4_ASAP7_75t_SL g594 ( .A(n_505), .B(n_514), .Y(n_594) );
AND2x4_ASAP7_75t_L g599 ( .A(n_505), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g608 ( .A(n_505), .Y(n_608) );
OR2x2_ASAP7_75t_L g614 ( .A(n_505), .B(n_514), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_505), .B(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_505), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_505), .B(n_596), .Y(n_730) );
OR2x2_ASAP7_75t_L g746 ( .A(n_505), .B(n_649), .Y(n_746) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_513), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g572 ( .A(n_513), .Y(n_572) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_513), .B(n_563), .Y(n_679) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_526), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_514), .B(n_527), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_514), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_514), .B(n_571), .Y(n_575) );
INVx3_ASAP7_75t_L g600 ( .A(n_514), .Y(n_600) );
INVx1_ASAP7_75t_L g633 ( .A(n_514), .Y(n_633) );
AND2x2_ASAP7_75t_L g713 ( .A(n_514), .B(n_577), .Y(n_713) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_527), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g598 ( .A(n_527), .Y(n_598) );
AND2x2_ASAP7_75t_L g623 ( .A(n_527), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g649 ( .A(n_527), .B(n_571), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_527), .B(n_600), .Y(n_666) );
INVx1_ASAP7_75t_L g672 ( .A(n_527), .Y(n_672) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
AOI222xp33_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_540), .B1(n_550), .B2(n_557), .C1(n_560), .C2(n_564), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_549), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_541), .B(n_610), .Y(n_661) );
AND2x4_ASAP7_75t_L g677 ( .A(n_541), .B(n_588), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_603), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_554), .A2(n_568), .B1(n_573), .B2(n_578), .C1(n_586), .C2(n_786), .Y(n_567) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g706 ( .A(n_555), .B(n_610), .Y(n_706) );
OR2x2_ASAP7_75t_L g749 ( .A(n_555), .B(n_655), .Y(n_749) );
AND2x2_ASAP7_75t_L g578 ( .A(n_556), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g639 ( .A(n_556), .Y(n_639) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_556), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_557), .A2(n_668), .B(n_673), .C(n_674), .Y(n_667) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g695 ( .A(n_559), .Y(n_695) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g625 ( .A(n_564), .Y(n_625) );
AND2x2_ASAP7_75t_L g609 ( .A(n_565), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_565), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_568), .A2(n_586), .A3(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_569), .A2(n_619), .B(n_663), .C(n_664), .Y(n_662) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
OR2x2_ASAP7_75t_L g651 ( .A(n_570), .B(n_600), .Y(n_651) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
BUFx2_ASAP7_75t_L g619 ( .A(n_579), .Y(n_619) );
AND2x2_ASAP7_75t_L g628 ( .A(n_579), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_580), .Y(n_610) );
AOI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_585), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_588), .B(n_645), .Y(n_737) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_601), .B(n_604), .C(n_626), .Y(n_589) );
INVxp33_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_592), .B(n_597), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g630 ( .A(n_594), .B(n_623), .Y(n_630) );
OR2x2_ASAP7_75t_L g606 ( .A(n_595), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_610), .Y(n_636) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g712 ( .A(n_596), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g735 ( .A(n_597), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_599), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_599), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g747 ( .A(n_599), .B(n_623), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_599), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g690 ( .A(n_600), .B(n_672), .Y(n_690) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g744 ( .A1(n_603), .A2(n_623), .A3(n_677), .B1(n_702), .B2(n_745), .C1(n_747), .C2(n_748), .Y(n_744) );
AOI211xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_609), .B(n_611), .C(n_620), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_607), .B(n_635), .Y(n_657) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g622 ( .A(n_608), .B(n_623), .Y(n_622) );
NOR2x1p5_ASAP7_75t_L g688 ( .A(n_608), .B(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_608), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_609), .A2(n_627), .B(n_630), .C(n_631), .Y(n_626) );
AND2x4_ASAP7_75t_L g645 ( .A(n_610), .B(n_629), .Y(n_645) );
INVx2_ASAP7_75t_L g655 ( .A(n_610), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_610), .B(n_644), .Y(n_675) );
AND2x2_ASAP7_75t_L g717 ( .A(n_610), .B(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_610), .B(n_734), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_610), .B(n_638), .Y(n_756) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B(n_617), .Y(n_611) );
AND2x2_ASAP7_75t_L g707 ( .A(n_613), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g635 ( .A(n_616), .Y(n_635) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_628), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g722 ( .A(n_628), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_634), .B(n_636), .C(n_637), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_635), .Y(n_719) );
INVx3_ASAP7_75t_SL g734 ( .A(n_638), .Y(n_734) );
NAND5xp2_ASAP7_75t_L g640 ( .A(n_641), .B(n_660), .C(n_667), .D(n_680), .E(n_691), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_646), .B1(n_650), .B2(n_652), .C1(n_656), .C2(n_658), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_643), .A2(n_724), .B1(n_728), .B2(n_729), .Y(n_723) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g673 ( .A(n_644), .B(n_645), .Y(n_673) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_654), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_655), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g692 ( .A(n_655), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g703 ( .A(n_655), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g733 ( .A(n_659), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g681 ( .A(n_666), .Y(n_681) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_677), .A2(n_681), .B1(n_682), .B2(n_686), .Y(n_680) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_677), .Y(n_728) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g694 ( .A(n_679), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g699 ( .A(n_681), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_SL g727 ( .A(n_690), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_715), .C(n_738), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_698), .B(n_714), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_710), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g739 ( .A(n_701), .B(n_727), .Y(n_739) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OAI321xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .A3(n_720), .B1(n_722), .B2(n_723), .C(n_731), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_729), .A2(n_751), .B1(n_755), .B2(n_756), .Y(n_750) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_740), .B(n_744), .C(n_750), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g784 ( .A(n_776), .Y(n_784) );
INVx3_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_SL g777 ( .A(n_778), .B(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
endmodule