module fake_jpeg_7645_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_2),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_30),
.C(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_18),
.C(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_60),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_23),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_29),
.B1(n_15),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_22),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_22),
.B1(n_18),
.B2(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_28),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_76),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_81),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_22),
.B(n_18),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_19),
.B(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_64),
.B1(n_53),
.B2(n_46),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_63),
.B1(n_19),
.B2(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_102),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_49),
.B(n_53),
.C(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_104),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_108),
.B(n_25),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_101),
.B1(n_68),
.B2(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_39),
.B(n_41),
.C(n_42),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_39),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_81),
.C(n_78),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_66),
.B(n_71),
.C(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_123),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_80),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_105),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_86),
.B1(n_113),
.B2(n_119),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_71),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_91),
.B(n_104),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_105),
.B(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_65),
.C(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_77),
.B1(n_73),
.B2(n_41),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_3),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_87),
.B(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_136),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_147),
.B(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_149),
.B1(n_58),
.B2(n_45),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_25),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_101),
.B1(n_108),
.B2(n_91),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_109),
.B1(n_120),
.B2(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_115),
.C(n_98),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_97),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_126),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_153),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_151),
.B1(n_135),
.B2(n_131),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_129),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_42),
.C(n_95),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_168),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_58),
.C(n_45),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_179),
.B1(n_58),
.B2(n_27),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_149),
.B1(n_151),
.B2(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_158),
.C(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_182),
.B(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_179),
.B1(n_153),
.B2(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_192),
.B1(n_195),
.B2(n_170),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_190),
.C(n_6),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_189),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_169),
.B1(n_155),
.B2(n_157),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_6),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_14),
.B1(n_13),
.B2(n_19),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_14),
.C(n_4),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_174),
.C(n_173),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_198),
.C(n_203),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_195),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_198),
.B1(n_9),
.B2(n_10),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_3),
.B(n_4),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_202),
.B(n_205),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_8),
.C(n_9),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_196),
.C(n_190),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_186),
.B(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_212),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_8),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_11),
.B(n_9),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_221),
.A2(n_10),
.B(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_223),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_227),
.Y(n_228)
);


endmodule