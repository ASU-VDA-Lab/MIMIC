module fake_jpeg_2604_n_442 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_57),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_59),
.B(n_90),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_68),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_5),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_91),
.Y(n_123)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_87),
.Y(n_151)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_34),
.B(n_8),
.Y(n_90)
);

CKINVDCx11_ASAP7_75t_R g91 ( 
.A(n_19),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_95),
.Y(n_180)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_26),
.Y(n_133)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_109),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_34),
.Y(n_103)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_107),
.B1(n_55),
.B2(n_57),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_108),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

NAND2xp67_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_54),
.Y(n_136)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_4),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_112),
.B(n_113),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_115),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_35),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_50),
.B1(n_47),
.B2(n_52),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_142),
.B1(n_160),
.B2(n_169),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_119),
.A2(n_135),
.B1(n_140),
.B2(n_153),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_126),
.A2(n_119),
.B1(n_118),
.B2(n_140),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_188),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_55),
.A2(n_43),
.B1(n_49),
.B2(n_28),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_134),
.A2(n_148),
.B1(n_157),
.B2(n_159),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_43),
.B1(n_53),
.B2(n_45),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_53),
.B1(n_45),
.B2(n_44),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_86),
.A2(n_44),
.B1(n_28),
.B2(n_51),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_82),
.A2(n_54),
.B1(n_51),
.B2(n_2),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_93),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_60),
.A2(n_99),
.B1(n_92),
.B2(n_89),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_95),
.A2(n_10),
.B1(n_13),
.B2(n_3),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_164),
.A2(n_165),
.B1(n_174),
.B2(n_175),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_71),
.A2(n_0),
.B1(n_12),
.B2(n_17),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_77),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_97),
.A2(n_101),
.B1(n_112),
.B2(n_110),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_73),
.B(n_85),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_113),
.A2(n_65),
.B1(n_81),
.B2(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_104),
.A2(n_107),
.B1(n_65),
.B2(n_81),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_74),
.A2(n_96),
.B1(n_56),
.B2(n_106),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_177),
.A2(n_187),
.B1(n_130),
.B2(n_185),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_56),
.B(n_64),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_64),
.B(n_59),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_64),
.B(n_59),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_176),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_68),
.A2(n_37),
.B1(n_25),
.B2(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_193),
.B(n_212),
.Y(n_259)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_196),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_139),
.C(n_125),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_221),
.Y(n_270)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_201),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_151),
.B(n_123),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_151),
.B(n_137),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_203),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_117),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_204),
.B(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_134),
.B1(n_126),
.B2(n_135),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_206),
.A2(n_236),
.B1(n_247),
.B2(n_219),
.Y(n_293)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_116),
.B(n_143),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_218),
.Y(n_258)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_213),
.B(n_237),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_127),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_221),
.B(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_226),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_159),
.A2(n_177),
.B(n_128),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_228),
.B(n_233),
.C(n_210),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_148),
.A2(n_164),
.B(n_157),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_229),
.A2(n_238),
.B1(n_247),
.B2(n_199),
.Y(n_292)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_232),
.Y(n_263)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_165),
.A2(n_132),
.B(n_120),
.C(n_158),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_167),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_235),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_172),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_130),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_156),
.A2(n_185),
.B1(n_179),
.B2(n_173),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_153),
.B(n_166),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_146),
.B(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_120),
.B(n_131),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_246),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_120),
.B(n_131),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_175),
.A2(n_37),
.B1(n_55),
.B2(n_25),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_122),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_121),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_133),
.B(n_178),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_207),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_261),
.B(n_259),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_217),
.A2(n_214),
.B1(n_228),
.B2(n_218),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_269),
.A2(n_284),
.B1(n_281),
.B2(n_271),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_286),
.C(n_262),
.Y(n_326)
);

AOI32xp33_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_195),
.A3(n_197),
.B1(n_189),
.B2(n_233),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_196),
.B(n_216),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_217),
.A2(n_214),
.B1(n_218),
.B2(n_227),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_210),
.Y(n_287)
);

OR2x4_ASAP7_75t_L g288 ( 
.A(n_195),
.B(n_229),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_252),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_245),
.B1(n_288),
.B2(n_284),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_238),
.B1(n_191),
.B2(n_211),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_297),
.A2(n_305),
.B1(n_308),
.B2(n_310),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_313),
.Y(n_335)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_260),
.B(n_208),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_303),
.B(n_311),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_223),
.B1(n_215),
.B2(n_243),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_304),
.A2(n_278),
.B1(n_282),
.B2(n_283),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_258),
.A2(n_194),
.B1(n_226),
.B2(n_231),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_306),
.A2(n_323),
.B(n_324),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_258),
.A2(n_291),
.B1(n_293),
.B2(n_269),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_258),
.A2(n_267),
.B1(n_252),
.B2(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_321),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_253),
.A2(n_294),
.B1(n_287),
.B2(n_270),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_314),
.A2(n_325),
.B1(n_308),
.B2(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_257),
.B(n_254),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_316),
.B(n_319),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_329),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_261),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_255),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_255),
.B(n_273),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_326),
.C(n_289),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_277),
.A2(n_281),
.B1(n_264),
.B2(n_280),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_281),
.A2(n_256),
.B1(n_272),
.B2(n_290),
.Y(n_325)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_327),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_289),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_278),
.Y(n_339)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_296),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_331),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_333),
.B(n_351),
.Y(n_362)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_345),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_295),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_341),
.B(n_338),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_328),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_283),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_301),
.C(n_309),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_300),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_348),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_312),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_298),
.Y(n_346)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_298),
.B(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_351),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_303),
.Y(n_352)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_352),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_324),
.A2(n_313),
.B(n_331),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_327),
.B(n_302),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_322),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_369),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_357),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_361),
.B(n_363),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_357),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_325),
.B1(n_309),
.B2(n_329),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_376),
.B1(n_352),
.B2(n_353),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_332),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_373),
.C(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_375),
.B(n_350),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_343),
.C(n_348),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_354),
.A2(n_349),
.B(n_340),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g377 ( 
.A(n_345),
.B(n_346),
.CI(n_344),
.CON(n_377),
.SN(n_377)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_377),
.B(n_344),
.CI(n_342),
.CON(n_380),
.SN(n_380)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_378),
.B(n_379),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_338),
.B(n_335),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_383),
.A2(n_367),
.B(n_359),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_368),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_389),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

NOR4xp25_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_355),
.C(n_356),
.D(n_335),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_393),
.C(n_369),
.Y(n_398)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_391),
.B(n_371),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_364),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_392),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_347),
.C(n_334),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_375),
.A2(n_337),
.B1(n_336),
.B2(n_347),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_394),
.A2(n_372),
.B1(n_366),
.B2(n_359),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_396),
.A2(n_401),
.B1(n_394),
.B2(n_391),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_362),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_382),
.B(n_378),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_387),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_381),
.A2(n_375),
.B1(n_360),
.B2(n_364),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_405),
.Y(n_413)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

XOR2x2_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_370),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_399),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_393),
.C(n_387),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_411),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_406),
.B(n_358),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_416),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_395),
.B(n_356),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_414),
.B(n_415),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_403),
.B(n_386),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_382),
.C(n_383),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_411),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_397),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g418 ( 
.A(n_416),
.B(n_400),
.CI(n_380),
.CON(n_418),
.SN(n_418)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_407),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_L g421 ( 
.A1(n_413),
.A2(n_402),
.B(n_403),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_401),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_408),
.Y(n_427)
);

AOI211xp5_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_397),
.B(n_409),
.C(n_384),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_426),
.B(n_430),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_428),
.A2(n_429),
.B1(n_422),
.B2(n_420),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_388),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_422),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_426),
.A2(n_428),
.B(n_417),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_432),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_434),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_418),
.Y(n_438)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_435),
.C(n_437),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_439),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_423),
.Y(n_442)
);


endmodule