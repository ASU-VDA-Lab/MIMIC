module fake_jpeg_27925_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_2),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_10),
.C(n_4),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_20),
.B1(n_16),
.B2(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_15),
.B1(n_20),
.B2(n_16),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_11),
.B(n_21),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_14),
.B1(n_36),
.B2(n_31),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_11),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_49),
.B1(n_50),
.B2(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_67),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_63),
.B1(n_60),
.B2(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_80),
.B1(n_71),
.B2(n_51),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_60),
.A3(n_56),
.B1(n_58),
.B2(n_3),
.C1(n_5),
.C2(n_6),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_69),
.C(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_53),
.C(n_61),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_24),
.C(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_70),
.B1(n_64),
.B2(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_73),
.B1(n_80),
.B2(n_36),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_44),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.C(n_43),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_17),
.A3(n_18),
.B1(n_40),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_43),
.C(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_10),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_89),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_2),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_17),
.C(n_18),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_97),
.C(n_101),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule