module fake_netlist_6_3695_n_1765 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1765);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1765;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_61),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_28),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_8),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_68),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_50),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_60),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_47),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_100),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_46),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_36),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_8),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_6),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_38),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_35),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_98),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_24),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_40),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_130),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_0),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_34),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_118),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_24),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_35),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_113),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_43),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_26),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_45),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_64),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_52),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_33),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_28),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_80),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_7),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_84),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_135),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_66),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_4),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_73),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_42),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_145),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_137),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_69),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_30),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_99),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_36),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_42),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_76),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_48),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_87),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_79),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_58),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_17),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_27),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_128),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_78),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_72),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_12),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_117),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_18),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_34),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_70),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_63),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_147),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_20),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_14),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_107),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_96),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_104),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_125),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_151),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_115),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_77),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_105),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_86),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_67),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_93),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_106),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_9),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_120),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_23),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_108),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_55),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_146),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_51),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_59),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_20),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_81),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_23),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_33),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_136),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_6),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_184),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_184),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_157),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_192),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_194),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_187),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_184),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_189),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_179),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_208),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_208),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_208),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_276),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_160),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_160),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_191),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_202),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_230),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_176),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_203),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_204),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_212),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_213),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_217),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_225),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_207),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_215),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_273),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_222),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_169),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_280),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_232),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_268),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_166),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_231),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_185),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_163),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_186),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_164),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_170),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_183),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_239),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_190),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_169),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_188),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_241),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_244),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_190),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_352),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_372),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_317),
.A2(n_272),
.B1(n_250),
.B2(n_238),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_366),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_237),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_318),
.A2(n_236),
.B1(n_308),
.B2(n_307),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_285),
.B(n_247),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_237),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_310),
.B1(n_308),
.B2(n_307),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_259),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_379),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_199),
.B(n_168),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_322),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_259),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_321),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_314),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_316),
.B(n_262),
.Y(n_428)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_319),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_320),
.B(n_168),
.Y(n_431)
);

BUFx8_ASAP7_75t_L g432 ( 
.A(n_339),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_315),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_156),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_313),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_342),
.B(n_156),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_322),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_337),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_377),
.B(n_175),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_325),
.B(n_193),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_325),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_343),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_336),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_338),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_197),
.B(n_195),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_445),
.B(n_338),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_331),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_368),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_340),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_424),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_390),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_200),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_385),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_429),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_199),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_346),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_340),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_429),
.B(n_220),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_432),
.B(n_344),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_431),
.A2(n_262),
.B1(n_285),
.B2(n_247),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_432),
.B(n_344),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_404),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_383),
.B1(n_234),
.B2(n_220),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_387),
.B(n_391),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_429),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_432),
.B(n_354),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_396),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

CKINVDCx6p67_ASAP7_75t_R g503 ( 
.A(n_435),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_384),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_431),
.A2(n_266),
.B1(n_234),
.B2(n_264),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_412),
.B(n_354),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_345),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_405),
.B(n_356),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_426),
.B(n_347),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_407),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_388),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_432),
.B(n_356),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_441),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_426),
.B(n_349),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_414),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

BUFx6f_ASAP7_75t_SL g525 ( 
.A(n_431),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_440),
.B(n_358),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_446),
.B(n_358),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_438),
.B(n_369),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_408),
.B(n_369),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_396),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_415),
.B(n_376),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_401),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_415),
.B(n_313),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_401),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_411),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_437),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_411),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_408),
.B(n_376),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_430),
.B(n_380),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_403),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_403),
.B(n_380),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_398),
.A2(n_299),
.B1(n_177),
.B2(n_180),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_410),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_398),
.A2(n_299),
.B1(n_295),
.B2(n_182),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_420),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_390),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_397),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_420),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_386),
.B(n_392),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_418),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_437),
.B(n_381),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_418),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_395),
.B(n_381),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_418),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_397),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_428),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_421),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_418),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_421),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_418),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_442),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_395),
.B(n_353),
.C(n_360),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_386),
.B(n_243),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_386),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_428),
.A2(n_305),
.B1(n_295),
.B2(n_310),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_442),
.B(n_175),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_392),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_434),
.Y(n_588)
);

CKINVDCx6p67_ASAP7_75t_R g589 ( 
.A(n_421),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_427),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_392),
.B(n_289),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_409),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_434),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_442),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_427),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_590),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_498),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_534),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_450),
.A2(n_341),
.B1(n_306),
.B2(n_209),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_545),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_531),
.B(n_421),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_449),
.A2(n_409),
.B(n_422),
.Y(n_606)
);

INVx8_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_596),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_572),
.B(n_158),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_545),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_534),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_544),
.B(n_422),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_482),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_169),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_158),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_549),
.B(n_434),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_455),
.B(n_159),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_508),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_548),
.B(n_159),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_576),
.B(n_544),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_532),
.A2(n_266),
.B1(n_257),
.B2(n_264),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_449),
.B(n_399),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_456),
.B(n_161),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_561),
.B(n_161),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_453),
.B(n_399),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_453),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_561),
.B(n_162),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_490),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_451),
.B(n_248),
.C(n_267),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_490),
.Y(n_633)
);

NAND3x1_ASAP7_75t_L g634 ( 
.A(n_554),
.B(n_350),
.C(n_351),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_551),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_470),
.B(n_399),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_470),
.B(n_221),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

BUFx5_ASAP7_75t_L g640 ( 
.A(n_461),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_468),
.B(n_221),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_561),
.B(n_162),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_468),
.B(n_257),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_538),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_492),
.B(n_211),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_517),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_457),
.A2(n_198),
.B1(n_201),
.B2(n_205),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_492),
.B(n_214),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_493),
.B(n_216),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_553),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_461),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_461),
.A2(n_543),
.B1(n_452),
.B2(n_546),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_546),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_476),
.B(n_509),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_561),
.B(n_165),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_494),
.B(n_219),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_552),
.B(n_165),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_494),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_500),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_500),
.B(n_223),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_229),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_464),
.A2(n_472),
.B(n_463),
.C(n_505),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_559),
.A2(n_196),
.B1(n_260),
.B2(n_180),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_570),
.B(n_167),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_515),
.B(n_245),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_508),
.B(n_355),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_510),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_515),
.B(n_249),
.Y(n_672)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_256),
.C(n_294),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_546),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_454),
.B(n_167),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_546),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_523),
.B(n_255),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_543),
.A2(n_175),
.B1(n_309),
.B2(n_169),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_524),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_542),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_523),
.B(n_284),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_528),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_589),
.B(n_275),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_528),
.B(n_292),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_452),
.A2(n_175),
.B1(n_309),
.B2(n_169),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_507),
.B(n_171),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_520),
.B(n_171),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_530),
.B(n_174),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_542),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_530),
.B(n_293),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_533),
.B(n_300),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_546),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_533),
.B(n_303),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_542),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_478),
.B(n_361),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_504),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_537),
.B(n_304),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_463),
.A2(n_363),
.B(n_362),
.C(n_439),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_537),
.B(n_539),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_475),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_539),
.B(n_174),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_520),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_463),
.B(n_169),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_527),
.B(n_286),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_588),
.B(n_309),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_475),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_562),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_585),
.B(n_286),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_583),
.B(n_433),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_460),
.B(n_506),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_582),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_433),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_488),
.B(n_253),
.C(n_274),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_522),
.B(n_433),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_479),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_469),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_503),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_460),
.B(n_301),
.C(n_287),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_529),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_479),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_541),
.B(n_287),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_481),
.B(n_290),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_525),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_522),
.B(n_439),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_582),
.B(n_444),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_525),
.A2(n_269),
.B1(n_206),
.B2(n_218),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_526),
.B(n_444),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_526),
.B(n_447),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_562),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_535),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_554),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_495),
.B(n_513),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_483),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_535),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_536),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_491),
.B(n_290),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_536),
.B(n_447),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_511),
.B(n_227),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_480),
.B(n_291),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_557),
.B(n_291),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_589),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_593),
.B(n_228),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_595),
.B(n_301),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_594),
.B(n_265),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_564),
.B(n_246),
.C(n_252),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_555),
.B(n_169),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_564),
.B(n_282),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_483),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_504),
.B(n_302),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_512),
.B(n_302),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_568),
.B(n_263),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_574),
.B(n_240),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_595),
.B(n_297),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_574),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_540),
.B(n_242),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_469),
.A2(n_261),
.B1(n_233),
.B2(n_235),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_540),
.B(n_254),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_550),
.B(n_281),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_512),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_550),
.B(n_297),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_555),
.B(n_258),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_558),
.B(n_309),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_709),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_732),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_556),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_734),
.A2(n_452),
.B1(n_469),
.B2(n_477),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_736),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_600),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_736),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_733),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_738),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_607),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_606),
.A2(n_558),
.B(n_563),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_739),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_603),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_600),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_598),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_623),
.B(n_556),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_610),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_646),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_629),
.B(n_563),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_469),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_608),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_613),
.B(n_503),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_496),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_599),
.Y(n_792)
);

AO22x1_ASAP7_75t_L g793 ( 
.A1(n_744),
.A2(n_579),
.B1(n_577),
.B2(n_182),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_674),
.Y(n_794)
);

INVx5_ASAP7_75t_L g795 ( 
.A(n_674),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_671),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_614),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_629),
.B(n_496),
.Y(n_798)
);

INVx8_ASAP7_75t_L g799 ( 
.A(n_607),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_615),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_SL g801 ( 
.A(n_666),
.B(n_305),
.C(n_277),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_656),
.B(n_497),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_720),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_656),
.B(n_497),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_698),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_620),
.A2(n_595),
.B(n_566),
.C(n_501),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_631),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_651),
.B(n_501),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_617),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_635),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_763),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_674),
.Y(n_812)
);

NAND2x2_ASAP7_75t_L g813 ( 
.A(n_722),
.B(n_612),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_644),
.B(n_577),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_639),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_600),
.B(n_579),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_607),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_654),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_704),
.B(n_469),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_654),
.B(n_677),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_650),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_726),
.B(n_670),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_633),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_677),
.B(n_514),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_694),
.B(n_606),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_637),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_680),
.A2(n_477),
.B1(n_169),
.B2(n_309),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_671),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_702),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_694),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_597),
.Y(n_831)
);

AND2x6_ASAP7_75t_SL g832 ( 
.A(n_753),
.B(n_477),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_618),
.Y(n_833)
);

CKINVDCx11_ASAP7_75t_R g834 ( 
.A(n_697),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_670),
.A2(n_477),
.B(n_586),
.C(n_487),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_640),
.B(n_514),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_680),
.A2(n_477),
.B1(n_458),
.B2(n_459),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_SL g838 ( 
.A(n_605),
.B(n_279),
.C(n_283),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_597),
.B(n_601),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_719),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_719),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_661),
.Y(n_842)
);

NAND2x1p5_ASAP7_75t_L g843 ( 
.A(n_726),
.B(n_581),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_669),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_601),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_618),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_754),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_728),
.B(n_571),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_708),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_662),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_620),
.A2(n_665),
.B(n_740),
.C(n_725),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_713),
.A2(n_474),
.B1(n_458),
.B2(n_473),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_665),
.A2(n_740),
.B(n_713),
.C(n_706),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_SL g854 ( 
.A1(n_712),
.A2(n_275),
.B1(n_5),
.B2(n_10),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_705),
.A2(n_581),
.B(n_518),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_718),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_719),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_712),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_675),
.B(n_571),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_640),
.B(n_516),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_678),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_640),
.B(n_581),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_640),
.B(n_516),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_697),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_660),
.A2(n_518),
.B(n_578),
.C(n_569),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_687),
.A2(n_473),
.B1(n_459),
.B2(n_462),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_723),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

INVx5_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_689),
.B(n_462),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_684),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_652),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_655),
.B(n_581),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_681),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_687),
.A2(n_467),
.B1(n_474),
.B2(n_487),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_737),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_735),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_718),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_640),
.B(n_569),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_735),
.B(n_571),
.Y(n_881)
);

AND2x6_ASAP7_75t_L g882 ( 
.A(n_625),
.B(n_578),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_735),
.B(n_565),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_640),
.B(n_486),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_602),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_758),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_659),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_727),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_673),
.B(n_565),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_724),
.B(n_275),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_673),
.B(n_565),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_730),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_752),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_701),
.B(n_486),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_731),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_682),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_653),
.B(n_489),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_741),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_SL g899 ( 
.A1(n_745),
.A2(n_690),
.B1(n_703),
.B2(n_685),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_691),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_667),
.B(n_467),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_653),
.B(n_489),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_609),
.A2(n_573),
.B1(n_587),
.B2(n_584),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_632),
.B(n_573),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_696),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_716),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_634),
.B(n_580),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_659),
.B(n_587),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_710),
.B(n_580),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_659),
.B(n_587),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_688),
.B(n_485),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_628),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_624),
.A2(n_584),
.B1(n_442),
.B2(n_573),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_742),
.B(n_499),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_707),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_636),
.B(n_584),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_659),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_SL g918 ( 
.A1(n_715),
.A2(n_729),
.B1(n_666),
.B2(n_647),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_619),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_624),
.A2(n_485),
.B1(n_465),
.B2(n_466),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_690),
.A2(n_465),
.B(n_466),
.C(n_471),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_638),
.B(n_465),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_749),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_641),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_676),
.B(n_485),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_659),
.B(n_502),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_643),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_766),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_747),
.B(n_502),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_721),
.B(n_499),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_757),
.B(n_502),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_624),
.A2(n_442),
.B1(n_484),
.B2(n_466),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_616),
.A2(n_442),
.B1(n_484),
.B2(n_471),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_746),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_627),
.B(n_471),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_645),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_711),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_659),
.B(n_499),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_714),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_649),
.A2(n_484),
.B1(n_519),
.B2(n_580),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_648),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_658),
.Y(n_942)
);

CKINVDCx6p67_ASAP7_75t_R g943 ( 
.A(n_626),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_707),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_707),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_663),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_707),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_664),
.B(n_580),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_668),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_672),
.B(n_519),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_679),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_748),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_700),
.A2(n_502),
.B(n_499),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_833),
.A2(n_622),
.B(n_630),
.C(n_642),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_833),
.A2(n_657),
.B(n_703),
.C(n_721),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_937),
.B(n_764),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_846),
.B(n_764),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_887),
.A2(n_700),
.B(n_765),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_887),
.A2(n_762),
.B(n_761),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_822),
.B(n_743),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_897),
.A2(n_902),
.B(n_804),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_795),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_846),
.A2(n_699),
.B(n_686),
.C(n_692),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_851),
.A2(n_695),
.B(n_683),
.C(n_693),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_918),
.A2(n_759),
.B1(n_751),
.B2(n_756),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_834),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_769),
.B(n_755),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_829),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_849),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_827),
.A2(n_760),
.B1(n_519),
.B2(n_502),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_855),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_844),
.B(n_499),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_817),
.B(n_519),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_781),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_853),
.A2(n_750),
.B(n_519),
.C(n_502),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_917),
.A2(n_948),
.B(n_863),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_799),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_859),
.B(n_4),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_917),
.A2(n_499),
.B(n_397),
.Y(n_979)
);

BUFx10_ASAP7_75t_L g980 ( 
.A(n_814),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_854),
.A2(n_10),
.B(n_11),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_890),
.A2(n_11),
.B(n_13),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_948),
.A2(n_397),
.B(n_567),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_795),
.A2(n_397),
.B(n_567),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_783),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_827),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_799),
.B(n_575),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_939),
.B(n_19),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_899),
.A2(n_21),
.B(n_22),
.C(n_25),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_868),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_811),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_888),
.B(n_21),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_892),
.B(n_25),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_895),
.B(n_898),
.Y(n_994)
);

AO32x1_ASAP7_75t_L g995 ( 
.A1(n_940),
.A2(n_31),
.A3(n_32),
.B1(n_39),
.B2(n_41),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_788),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_847),
.B(n_31),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_946),
.B(n_951),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_789),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_797),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_805),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_817),
.B(n_575),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_838),
.A2(n_39),
.B(n_41),
.C(n_44),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_782),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_795),
.A2(n_397),
.B(n_567),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_799),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_SL g1007 ( 
.A(n_795),
.B(n_575),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_812),
.A2(n_575),
.B(n_567),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_785),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_812),
.A2(n_575),
.B(n_567),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_L g1011 ( 
.A(n_801),
.B(n_44),
.C(n_560),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_790),
.B(n_560),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_800),
.Y(n_1013)
);

AOI222xp33_ASAP7_75t_L g1014 ( 
.A1(n_885),
.A2(n_49),
.B1(n_57),
.B2(n_62),
.C1(n_82),
.C2(n_88),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_946),
.B(n_89),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_907),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_812),
.A2(n_560),
.B(n_109),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_912),
.B(n_90),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_838),
.A2(n_110),
.B(n_111),
.C(n_112),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_822),
.B(n_560),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_839),
.B(n_560),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_777),
.A2(n_124),
.B(n_127),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_807),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_831),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_845),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_877),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_812),
.A2(n_132),
.B(n_133),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_796),
.Y(n_1029)
);

BUFx8_ASAP7_75t_L g1030 ( 
.A(n_792),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_796),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_794),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_854),
.A2(n_134),
.B1(n_144),
.B2(n_148),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_828),
.B(n_149),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_779),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_787),
.B(n_150),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_897),
.A2(n_902),
.B(n_804),
.Y(n_1037)
);

BUFx4f_ASAP7_75t_L g1038 ( 
.A(n_943),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_871),
.A2(n_154),
.B(n_906),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_857),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_823),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_819),
.A2(n_787),
.B1(n_923),
.B2(n_949),
.Y(n_1042)
);

AOI221xp5_ASAP7_75t_L g1043 ( 
.A1(n_801),
.A2(n_793),
.B1(n_828),
.B2(n_865),
.C(n_869),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_942),
.A2(n_927),
.B(n_802),
.C(n_941),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_857),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_884),
.A2(n_856),
.B(n_880),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_784),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_879),
.B(n_934),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_776),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_776),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_809),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_810),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_879),
.B(n_952),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_794),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_878),
.B(n_883),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_883),
.B(n_881),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_815),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_819),
.B(n_826),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_842),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_803),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_SL g1061 ( 
.A(n_816),
.B(n_862),
.C(n_872),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_772),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_772),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_802),
.B(n_850),
.Y(n_1064)
);

CKINVDCx16_ASAP7_75t_R g1065 ( 
.A(n_930),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_901),
.B(n_881),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_908),
.A2(n_910),
.B(n_825),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_919),
.B(n_886),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_840),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_884),
.A2(n_856),
.B(n_880),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_767),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_780),
.B(n_907),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_835),
.A2(n_911),
.B(n_924),
.C(n_768),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_780),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_840),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_770),
.A2(n_837),
.B1(n_786),
.B2(n_867),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_813),
.A2(n_936),
.B1(n_907),
.B2(n_909),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_774),
.Y(n_1078)
);

CKINVDCx8_ASAP7_75t_R g1079 ( 
.A(n_832),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_936),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_836),
.A2(n_861),
.B(n_864),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_936),
.Y(n_1082)
);

CKINVDCx6p67_ASAP7_75t_R g1083 ( 
.A(n_909),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_848),
.B(n_860),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_848),
.B(n_860),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_821),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_771),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_894),
.B(n_775),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_925),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_806),
.A2(n_921),
.B(n_825),
.C(n_866),
.Y(n_1090)
);

BUFx12f_ASAP7_75t_L g1091 ( 
.A(n_925),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_778),
.B(n_875),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_818),
.B(n_841),
.Y(n_1093)
);

AO32x2_ASAP7_75t_L g1094 ( 
.A1(n_940),
.A2(n_932),
.A3(n_913),
.B1(n_777),
.B2(n_882),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_836),
.A2(n_861),
.B(n_864),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_873),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_914),
.A2(n_950),
.B(n_904),
.C(n_928),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_770),
.A2(n_837),
.B1(n_786),
.B2(n_867),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_1004),
.A2(n_891),
.B1(n_889),
.B2(n_904),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_959),
.A2(n_950),
.B(n_894),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1025),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_1014),
.B(n_955),
.C(n_967),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1004),
.B(n_900),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_1030),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_962),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1009),
.Y(n_1107)
);

BUFx5_ASAP7_75t_L g1108 ( 
.A(n_1078),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_958),
.A2(n_830),
.B(n_910),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_962),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_976),
.A2(n_830),
.B(n_818),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1070),
.A2(n_824),
.B(n_808),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1030),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_985),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_991),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_SL g1116 ( 
.A1(n_1039),
.A2(n_905),
.B(n_875),
.C(n_858),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_1082),
.B(n_858),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1067),
.A2(n_808),
.B(n_820),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1064),
.B(n_798),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1081),
.A2(n_820),
.B(n_953),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_L g1121 ( 
.A(n_1049),
.B(n_843),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1095),
.A2(n_953),
.B(n_835),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_996),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_981),
.A2(n_798),
.B1(n_891),
.B2(n_889),
.C(n_841),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_956),
.B(n_818),
.Y(n_1125)
);

AND2x2_ASAP7_75t_SL g1126 ( 
.A(n_1065),
.B(n_1038),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_999),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1000),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_994),
.B(n_998),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_954),
.A2(n_935),
.B(n_896),
.C(n_905),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_964),
.A2(n_876),
.B(n_852),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1090),
.A2(n_818),
.B(n_938),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1076),
.A2(n_1098),
.B(n_1073),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_1001),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_961),
.A2(n_909),
.B(n_926),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1056),
.B(n_773),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1088),
.B(n_852),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1076),
.A2(n_874),
.B(n_931),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_957),
.B(n_873),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_965),
.A2(n_876),
.B(n_913),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1056),
.B(n_873),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1013),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1098),
.A2(n_975),
.B(n_1044),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_981),
.A2(n_932),
.B1(n_920),
.B2(n_933),
.C(n_944),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_986),
.A2(n_933),
.B1(n_915),
.B2(n_843),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1037),
.A2(n_929),
.B(n_931),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1024),
.Y(n_1147)
);

CKINVDCx16_ASAP7_75t_R g1148 ( 
.A(n_1060),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1055),
.B(n_791),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1066),
.B(n_882),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_986),
.A2(n_915),
.B1(n_929),
.B2(n_874),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1023),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1058),
.B(n_903),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1041),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_960),
.A2(n_1042),
.B1(n_1036),
.B2(n_1014),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_965),
.A2(n_882),
.B(n_922),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1039),
.A2(n_947),
.B(n_945),
.C(n_944),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1018),
.A2(n_947),
.B(n_945),
.C(n_791),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_960),
.A2(n_882),
.B1(n_922),
.B2(n_791),
.Y(n_1160)
);

AO22x2_ASAP7_75t_L g1161 ( 
.A1(n_1011),
.A2(n_882),
.B1(n_922),
.B2(n_916),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1029),
.B(n_1045),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_963),
.A2(n_870),
.B(n_922),
.C(n_916),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_1049),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1097),
.A2(n_922),
.B(n_916),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_970),
.A2(n_870),
.B(n_791),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_SL g1167 ( 
.A(n_1006),
.B(n_870),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1079),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1048),
.B(n_916),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1022),
.A2(n_916),
.B(n_791),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1053),
.B(n_870),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1059),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_966),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1071),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_983),
.A2(n_1072),
.B(n_1010),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1068),
.B(n_1092),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_997),
.A2(n_1016),
.B1(n_1011),
.B2(n_1080),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_992),
.B(n_993),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_988),
.B(n_968),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_970),
.A2(n_987),
.B(n_1015),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_978),
.B(n_1040),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_982),
.B(n_1077),
.C(n_1033),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1084),
.A2(n_1085),
.B(n_973),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_969),
.B(n_971),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_982),
.B(n_989),
.C(n_1003),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1061),
.A2(n_1019),
.B(n_1043),
.C(n_1034),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1021),
.A2(n_972),
.B(n_979),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_980),
.B(n_1089),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_977),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1055),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_SL g1191 ( 
.A1(n_995),
.A2(n_1075),
.B(n_1069),
.C(n_1032),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1007),
.A2(n_1012),
.B(n_1017),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1027),
.A2(n_1087),
.B(n_1086),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_990),
.Y(n_1194)
);

AO32x2_ASAP7_75t_L g1195 ( 
.A1(n_1033),
.A2(n_995),
.A3(n_1094),
.B1(n_1062),
.B2(n_1054),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1049),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1047),
.B(n_1028),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1035),
.B(n_1051),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1052),
.B(n_1057),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1200)
);

CKINVDCx11_ASAP7_75t_R g1201 ( 
.A(n_1050),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1008),
.A2(n_984),
.B(n_1005),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1093),
.A2(n_1002),
.B(n_1032),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1096),
.B(n_1062),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_980),
.B(n_1074),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1094),
.A2(n_1083),
.B(n_1016),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_977),
.B(n_1050),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1096),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_SL g1209 ( 
.A1(n_995),
.A2(n_1094),
.B(n_1016),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1038),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1050),
.B(n_1091),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1063),
.B(n_1096),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_977),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1054),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1020),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_987),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1020),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_987),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1046),
.A2(n_1070),
.B(n_1067),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1046),
.A2(n_1070),
.B(n_1067),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_959),
.A2(n_917),
.B(n_887),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_955),
.A2(n_851),
.B(n_967),
.C(n_899),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1056),
.B(n_1055),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_SL g1225 ( 
.A(n_981),
.B(n_1065),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_974),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_974),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_SL g1228 ( 
.A1(n_1073),
.A2(n_851),
.B(n_853),
.C(n_1039),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_959),
.A2(n_917),
.B(n_887),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1046),
.A2(n_1070),
.B(n_1067),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_991),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_975),
.A2(n_851),
.A3(n_853),
.B(n_964),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_959),
.A2(n_917),
.B(n_887),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_SL g1234 ( 
.A1(n_957),
.A2(n_890),
.B(n_992),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_967),
.B(n_994),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_967),
.B(n_994),
.Y(n_1236)
);

O2A1O1Ixp5_ASAP7_75t_L g1237 ( 
.A1(n_967),
.A2(n_851),
.B(n_605),
.C(n_853),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1046),
.A2(n_1070),
.B(n_1067),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1230),
.A2(n_1238),
.B(n_1122),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1231),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1165),
.A2(n_1157),
.B(n_1163),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1225),
.A2(n_1103),
.B1(n_1236),
.B2(n_1235),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1182),
.A2(n_1225),
.B1(n_1185),
.B2(n_1156),
.Y(n_1244)
);

BUFx4f_ASAP7_75t_SL g1245 ( 
.A(n_1134),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1170),
.A2(n_1112),
.B(n_1109),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1237),
.A2(n_1223),
.B(n_1178),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1185),
.A2(n_1228),
.B1(n_1133),
.B2(n_1186),
.C(n_1177),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1128),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1224),
.B(n_1190),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1224),
.B(n_1126),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1143),
.A2(n_1158),
.A3(n_1101),
.B(n_1124),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1131),
.A2(n_1140),
.B(n_1145),
.C(n_1157),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1206),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_SL g1256 ( 
.A(n_1125),
.B(n_1171),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1131),
.A2(n_1140),
.B1(n_1176),
.B2(n_1100),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1183),
.B(n_1180),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1222),
.A2(n_1233),
.B(n_1229),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1139),
.B(n_1154),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1145),
.A2(n_1152),
.B1(n_1176),
.B2(n_1148),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1164),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1162),
.B(n_1149),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1099),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1136),
.B(n_1181),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1119),
.A2(n_1144),
.B(n_1138),
.C(n_1137),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1165),
.A2(n_1118),
.B(n_1146),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1202),
.A2(n_1175),
.B(n_1135),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1164),
.B(n_1102),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1119),
.A2(n_1137),
.B1(n_1179),
.B2(n_1226),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1179),
.A2(n_1194),
.B1(n_1227),
.B2(n_1172),
.Y(n_1272)
);

AOI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1169),
.A2(n_1151),
.B(n_1193),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1166),
.A2(n_1111),
.B(n_1187),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1193),
.A2(n_1132),
.B(n_1116),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1217),
.A2(n_1188),
.B1(n_1123),
.B2(n_1127),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1234),
.A2(n_1192),
.B(n_1209),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1142),
.A2(n_1153),
.B1(n_1174),
.B2(n_1155),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1160),
.A2(n_1152),
.B(n_1219),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1144),
.A2(n_1130),
.B(n_1121),
.C(n_1197),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1210),
.A2(n_1218),
.B1(n_1147),
.B2(n_1107),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1201),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1198),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1200),
.A2(n_1199),
.B(n_1232),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1189),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1141),
.B(n_1205),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1200),
.B(n_1216),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1161),
.A2(n_1117),
.B1(n_1115),
.B2(n_1108),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1189),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1161),
.A2(n_1203),
.B(n_1215),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1232),
.A2(n_1191),
.B(n_1214),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1211),
.A2(n_1150),
.B1(n_1213),
.B2(n_1141),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1204),
.A2(n_1208),
.B(n_1212),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1108),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1204),
.A2(n_1150),
.B(n_1106),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1108),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1106),
.A2(n_1110),
.B(n_1108),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1105),
.A2(n_1113),
.B(n_1196),
.C(n_1211),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1108),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1207),
.B(n_1211),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1207),
.B(n_1189),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1232),
.A2(n_1195),
.B(n_1110),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1168),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1195),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1173),
.B(n_1195),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1114),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1308)
);

INVx6_ASAP7_75t_L g1309 ( 
.A(n_1164),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1231),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1201),
.Y(n_1311)
);

AO221x2_ASAP7_75t_L g1312 ( 
.A1(n_1185),
.A2(n_1033),
.B1(n_986),
.B2(n_1177),
.C(n_1103),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1162),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1165),
.A2(n_1157),
.B(n_1163),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1201),
.Y(n_1316)
);

OA21x2_ASAP7_75t_L g1317 ( 
.A1(n_1143),
.A2(n_1221),
.B(n_1220),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1114),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1223),
.A2(n_1186),
.B(n_1103),
.C(n_851),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1183),
.A2(n_1157),
.B(n_1178),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1135),
.A2(n_1138),
.B(n_1109),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1103),
.A2(n_981),
.B1(n_1182),
.B2(n_854),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_SL g1323 ( 
.A(n_1134),
.Y(n_1323)
);

INVx5_ASAP7_75t_L g1324 ( 
.A(n_1164),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1167),
.B(n_1016),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1231),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1114),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1201),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1135),
.A2(n_1138),
.B(n_1109),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1231),
.Y(n_1331)
);

OAI222xp33_ASAP7_75t_L g1332 ( 
.A1(n_1156),
.A2(n_854),
.B1(n_986),
.B2(n_899),
.C1(n_734),
.C2(n_744),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1165),
.A2(n_1157),
.B(n_1163),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_L g1334 ( 
.A(n_1104),
.B(n_805),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1150),
.B(n_1141),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1223),
.A2(n_1186),
.B(n_1103),
.C(n_851),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1165),
.A2(n_1157),
.B(n_1163),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1162),
.B(n_1149),
.Y(n_1339)
);

BUFx2_ASAP7_75t_SL g1340 ( 
.A(n_1164),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1114),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1114),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1143),
.A2(n_1158),
.A3(n_1163),
.B(n_851),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1149),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1235),
.B(n_859),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1201),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1114),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1206),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1114),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1103),
.A2(n_885),
.B1(n_605),
.B2(n_315),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1162),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1150),
.B(n_1141),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1231),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1223),
.A2(n_1186),
.B(n_1103),
.C(n_851),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1103),
.A2(n_1223),
.B(n_605),
.C(n_1186),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1235),
.B(n_859),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1120),
.A2(n_1221),
.B(n_1220),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1261),
.B(n_1347),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1359),
.B(n_1266),
.Y(n_1362)
);

O2A1O1Ixp5_ASAP7_75t_L g1363 ( 
.A1(n_1243),
.A2(n_1332),
.B(n_1247),
.C(n_1321),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1353),
.A2(n_1322),
.B1(n_1244),
.B2(n_1283),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1257),
.B(n_1313),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1265),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_1283),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1287),
.B(n_1251),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1301),
.B(n_1296),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1358),
.A2(n_1357),
.B(n_1337),
.C(n_1319),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1325),
.A2(n_1280),
.B(n_1249),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1372)
);

CKINVDCx6p67_ASAP7_75t_R g1373 ( 
.A(n_1311),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1252),
.B(n_1264),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1354),
.B(n_1264),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1322),
.A2(n_1244),
.B1(n_1243),
.B2(n_1276),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1335),
.B(n_1355),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1335),
.B(n_1355),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1311),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1334),
.B(n_1250),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1271),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1281),
.B(n_1284),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1263),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1255),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1272),
.B(n_1248),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1335),
.B(n_1355),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1319),
.A2(n_1337),
.B(n_1357),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1306),
.B(n_1241),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1278),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1263),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1262),
.A2(n_1258),
.B1(n_1289),
.B2(n_1272),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1254),
.A2(n_1271),
.B(n_1259),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1301),
.B(n_1318),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1255),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1329),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1310),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1254),
.A2(n_1259),
.B(n_1280),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1258),
.A2(n_1331),
.B1(n_1326),
.B2(n_1356),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1349),
.B(n_1352),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1351),
.A2(n_1312),
.B(n_1320),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1267),
.A2(n_1312),
.B(n_1273),
.C(n_1291),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1267),
.A2(n_1299),
.B(n_1279),
.C(n_1293),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1294),
.A2(n_1282),
.B(n_1259),
.C(n_1307),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1260),
.A2(n_1274),
.B(n_1317),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1324),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1260),
.A2(n_1274),
.B(n_1317),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1304),
.A2(n_1323),
.B1(n_1245),
.B2(n_1270),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1328),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_SL g1409 ( 
.A1(n_1351),
.A2(n_1256),
.B(n_1292),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1341),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1329),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1240),
.A2(n_1239),
.B(n_1350),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1344),
.B(n_1302),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1275),
.A2(n_1324),
.B(n_1277),
.C(n_1305),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1309),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_1277),
.B(n_1360),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1239),
.A2(n_1360),
.B(n_1350),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1303),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1242),
.A2(n_1338),
.B1(n_1333),
.B2(n_1315),
.C(n_1316),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1285),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1308),
.A2(n_1343),
.B(n_1314),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1316),
.Y(n_1424)
);

AOI221x1_ASAP7_75t_SL g1425 ( 
.A1(n_1305),
.A2(n_1300),
.B1(n_1295),
.B2(n_1323),
.C(n_1245),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1345),
.B(n_1340),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_L g1427 ( 
.A(n_1348),
.B(n_1297),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1345),
.B(n_1242),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1348),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1292),
.B(n_1345),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1246),
.A2(n_1308),
.B(n_1343),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1292),
.B(n_1288),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1345),
.B(n_1333),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1298),
.B(n_1253),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1330),
.A2(n_1253),
.B(n_1269),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1268),
.A2(n_1327),
.B1(n_1336),
.B2(n_1314),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1342),
.A2(n_851),
.B(n_1319),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1342),
.A2(n_1358),
.B(n_1103),
.C(n_981),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1261),
.B(n_1347),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1358),
.A2(n_1103),
.B(n_1332),
.C(n_1223),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1301),
.B(n_1296),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1353),
.A2(n_1322),
.B1(n_1244),
.B2(n_885),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1261),
.B(n_1347),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1306),
.A2(n_1178),
.B(n_890),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1319),
.A2(n_851),
.B(n_1337),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1353),
.A2(n_1322),
.B1(n_1244),
.B2(n_885),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1392),
.B(n_1397),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1384),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1419),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1412),
.A2(n_1418),
.B(n_1423),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1394),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1370),
.A2(n_1441),
.B(n_1387),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1419),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1381),
.B(n_1401),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1421),
.Y(n_1459)
);

OAI33xp33_ASAP7_75t_L g1460 ( 
.A1(n_1443),
.A2(n_1447),
.A3(n_1376),
.B1(n_1364),
.B2(n_1398),
.B3(n_1441),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1428),
.B(n_1435),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1363),
.A2(n_1446),
.B(n_1439),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1424),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1401),
.B(n_1366),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1371),
.B(n_1438),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1404),
.A2(n_1406),
.B(n_1436),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1420),
.B(n_1414),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1363),
.A2(n_1439),
.B(n_1426),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1410),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1379),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1408),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1399),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1370),
.A2(n_1391),
.B1(n_1402),
.B2(n_1375),
.C(n_1365),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1417),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1372),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1437),
.A2(n_1385),
.B(n_1382),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1369),
.B(n_1442),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1417),
.B(n_1388),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1369),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1431),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1402),
.B(n_1403),
.C(n_1380),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1431),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1442),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1396),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1405),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1413),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1393),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1374),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1361),
.B(n_1444),
.Y(n_1489)
);

BUFx4f_ASAP7_75t_SL g1490 ( 
.A(n_1395),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1425),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1440),
.B(n_1362),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1459),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1478),
.B(n_1368),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1450),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1459),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1480),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1461),
.B(n_1427),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1452),
.B(n_1415),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1449),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1480),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1455),
.A2(n_1411),
.B1(n_1373),
.B2(n_1407),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1453),
.B(n_1478),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1454),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1461),
.B(n_1422),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1459),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1453),
.B(n_1386),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1405),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1481),
.A2(n_1383),
.B(n_1429),
.Y(n_1509)
);

INVx3_ASAP7_75t_SL g1510 ( 
.A(n_1465),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1465),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1482),
.Y(n_1512)
);

AND2x4_ASAP7_75t_SL g1513 ( 
.A(n_1448),
.B(n_1390),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1481),
.B(n_1460),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1461),
.B(n_1390),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1377),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1450),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1456),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1453),
.B(n_1378),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1460),
.A2(n_1411),
.B1(n_1367),
.B2(n_1416),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1473),
.A2(n_1416),
.B1(n_1400),
.B2(n_1445),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1478),
.B(n_1400),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1458),
.B(n_1409),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1514),
.B(n_1462),
.C(n_1473),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1514),
.A2(n_1465),
.B1(n_1462),
.B2(n_1448),
.Y(n_1526)
);

NAND2x1_ASAP7_75t_L g1527 ( 
.A(n_1518),
.B(n_1448),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1502),
.A2(n_1458),
.B1(n_1465),
.B2(n_1464),
.C(n_1448),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1523),
.A2(n_1465),
.B1(n_1448),
.B2(n_1467),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1523),
.A2(n_1467),
.B(n_1464),
.C(n_1491),
.Y(n_1532)
);

AOI33xp33_ASAP7_75t_L g1533 ( 
.A1(n_1520),
.A2(n_1467),
.A3(n_1489),
.B1(n_1469),
.B2(n_1492),
.B3(n_1471),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1521),
.A2(n_1465),
.B1(n_1491),
.B2(n_1457),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1510),
.A2(n_1457),
.B1(n_1483),
.B2(n_1479),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1517),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1500),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1517),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1515),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1502),
.A2(n_1488),
.B1(n_1484),
.B2(n_1475),
.C(n_1489),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1543)
);

AOI222xp33_ASAP7_75t_L g1544 ( 
.A1(n_1521),
.A2(n_1490),
.B1(n_1489),
.B2(n_1492),
.C1(n_1484),
.C2(n_1487),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1508),
.Y(n_1545)
);

AOI222xp33_ASAP7_75t_L g1546 ( 
.A1(n_1520),
.A2(n_1490),
.B1(n_1492),
.B2(n_1487),
.C1(n_1472),
.C2(n_1486),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1511),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1497),
.A2(n_1451),
.B(n_1474),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1504),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1518),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1485),
.C(n_1451),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1493),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1503),
.B(n_1499),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1496),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1509),
.A2(n_1468),
.B(n_1469),
.C(n_1476),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1496),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1506),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1494),
.B(n_1476),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1553),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1553),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1508),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1542),
.B(n_1516),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1551),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1530),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1522),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1549),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1547),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1545),
.Y(n_1571)
);

AOI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1550),
.A2(n_1524),
.B(n_1501),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1508),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1550),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1528),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1577)
);

AND4x1_ASAP7_75t_L g1578 ( 
.A(n_1525),
.B(n_1522),
.C(n_1463),
.D(n_1470),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1548),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1468),
.C(n_1522),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1556),
.A2(n_1466),
.B(n_1512),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

AND2x6_ASAP7_75t_SL g1585 ( 
.A(n_1543),
.B(n_1463),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1511),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1533),
.A2(n_1505),
.B(n_1513),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1559),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1535),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1538),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1547),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1581),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1585),
.B(n_1463),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1554),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1560),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1587),
.A2(n_1529),
.B1(n_1536),
.B2(n_1526),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1586),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1568),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1572),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1568),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1541),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1561),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1562),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1591),
.B(n_1534),
.Y(n_1610)
);

AND2x4_ASAP7_75t_SL g1611 ( 
.A(n_1586),
.B(n_1557),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1577),
.B(n_1541),
.Y(n_1612)
);

NAND2x1_ASAP7_75t_L g1613 ( 
.A(n_1563),
.B(n_1557),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1507),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1565),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1565),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1563),
.B(n_1554),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1564),
.A2(n_1531),
.B1(n_1544),
.B2(n_1552),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1569),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1569),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1566),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1575),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1575),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_1507),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1563),
.B(n_1545),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1507),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1566),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1573),
.B(n_1557),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1589),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1592),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.B(n_1573),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1620),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1573),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1603),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1597),
.A2(n_1546),
.B1(n_1586),
.B2(n_1510),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1626),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1605),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1606),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1614),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1615),
.B(n_1592),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1611),
.B(n_1573),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1610),
.B(n_1598),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1610),
.B(n_1573),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1604),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1610),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1598),
.B(n_1573),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1593),
.B(n_1589),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1612),
.B(n_1585),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1614),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1624),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1602),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1519),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1632),
.B(n_1519),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1608),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1608),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1643),
.B(n_1616),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1640),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1647),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1640),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1654),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1657),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1648),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1617),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1647),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1648),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1654),
.B(n_1598),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1638),
.A2(n_1607),
.B1(n_1602),
.B2(n_1634),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1642),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1641),
.A2(n_1578),
.B1(n_1613),
.B2(n_1598),
.C(n_1570),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1578),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1664),
.A2(n_1613),
.B1(n_1595),
.B2(n_1619),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1635),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1649),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1636),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1644),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1671),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1671),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1687),
.A2(n_1659),
.B(n_1660),
.Y(n_1698)
);

AOI322xp5_ASAP7_75t_L g1699 ( 
.A1(n_1692),
.A2(n_1650),
.A3(n_1609),
.B1(n_1600),
.B2(n_1595),
.C1(n_1619),
.C2(n_1574),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1637),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1678),
.B(n_1659),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1674),
.B(n_1645),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1673),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1670),
.A2(n_1660),
.B1(n_1668),
.B2(n_1667),
.C(n_1645),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1672),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1686),
.A2(n_1607),
.B(n_1602),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1694),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1681),
.A2(n_1651),
.B(n_1639),
.C(n_1602),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1689),
.B(n_1639),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1684),
.A2(n_1681),
.B(n_1690),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1690),
.B(n_1651),
.Y(n_1712)
);

NOR2x1p5_ASAP7_75t_L g1713 ( 
.A(n_1680),
.B(n_1570),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1695),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1711),
.B(n_1689),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1712),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1701),
.B(n_1674),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1712),
.B(n_1696),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1709),
.B(n_1698),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1703),
.B(n_1683),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1700),
.B(n_1683),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1708),
.B(n_1675),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1697),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1718),
.A2(n_1710),
.B1(n_1704),
.B2(n_1713),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1715),
.A2(n_1707),
.B1(n_1705),
.B2(n_1702),
.C(n_1675),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1723),
.A2(n_1685),
.B(n_1677),
.Y(n_1728)
);

OAI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1716),
.A2(n_1699),
.B1(n_1694),
.B2(n_1685),
.C(n_1693),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1693),
.B(n_1677),
.C(n_1679),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1717),
.B(n_1682),
.C(n_1679),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1720),
.A2(n_1691),
.B(n_1682),
.Y(n_1732)
);

AO22x1_ASAP7_75t_L g1733 ( 
.A1(n_1720),
.A2(n_1691),
.B1(n_1607),
.B2(n_1668),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1719),
.A2(n_1570),
.B1(n_1582),
.B2(n_1574),
.Y(n_1734)
);

AOI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1729),
.A2(n_1725),
.B(n_1714),
.C(n_1724),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1726),
.B(n_1722),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1733),
.B(n_1646),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1731),
.Y(n_1738)
);

AOI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1730),
.A2(n_1667),
.B(n_1656),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1738),
.A2(n_1728),
.B(n_1732),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1736),
.B(n_1727),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1737),
.Y(n_1742)
);

NOR2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1735),
.B(n_1646),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1739),
.B(n_1653),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1738),
.A2(n_1734),
.B(n_1656),
.Y(n_1745)
);

AOI322xp5_ASAP7_75t_L g1746 ( 
.A1(n_1741),
.A2(n_1658),
.A3(n_1609),
.B1(n_1600),
.B2(n_1662),
.C1(n_1649),
.C2(n_1607),
.Y(n_1746)
);

OAI322xp33_ASAP7_75t_L g1747 ( 
.A1(n_1740),
.A2(n_1662),
.A3(n_1663),
.B1(n_1669),
.B2(n_1609),
.C1(n_1658),
.C2(n_1596),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1744),
.B(n_1618),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1745),
.A2(n_1742),
.B1(n_1743),
.B2(n_1663),
.C(n_1669),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_R g1750 ( 
.A(n_1742),
.B(n_1571),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1748),
.B(n_1750),
.Y(n_1751)
);

AOI332xp33_ASAP7_75t_L g1752 ( 
.A1(n_1749),
.A2(n_1618),
.A3(n_1621),
.B1(n_1622),
.B2(n_1631),
.B3(n_1625),
.C1(n_1627),
.C2(n_1633),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1747),
.B(n_1537),
.C(n_1621),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1751),
.B(n_1746),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1753),
.B1(n_1752),
.B2(n_1631),
.C(n_1625),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1755),
.Y(n_1756)
);

OAI31xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1756),
.A2(n_1634),
.A3(n_1630),
.B(n_1629),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1757),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1756),
.B(n_1622),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1759),
.B(n_1627),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1633),
.B(n_1630),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1761),
.A2(n_1629),
.B1(n_1623),
.B2(n_1571),
.Y(n_1762)
);

AOI322xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1584),
.A3(n_1583),
.B1(n_1579),
.B2(n_1666),
.C1(n_1665),
.C2(n_1539),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1762),
.A2(n_1596),
.B1(n_1584),
.B2(n_1583),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1763),
.B(n_1584),
.C(n_1583),
.Y(n_1765)
);


endmodule