module real_jpeg_6213_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_1),
.A2(n_39),
.B1(n_72),
.B2(n_196),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_1),
.A2(n_80),
.B1(n_196),
.B2(n_313),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_1),
.A2(n_196),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_91),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_3),
.A2(n_109),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_3),
.A2(n_109),
.B1(n_261),
.B2(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_3),
.A2(n_109),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_4),
.A2(n_240),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_4),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_4),
.A2(n_273),
.B1(n_287),
.B2(n_291),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_4),
.A2(n_102),
.B1(n_273),
.B2(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_4),
.A2(n_111),
.B1(n_208),
.B2(n_273),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_5),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_152),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_5),
.A2(n_152),
.B1(n_198),
.B2(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_5),
.A2(n_152),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_7),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_7),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_7),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_34),
.B1(n_57),
.B2(n_161),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_9),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_9),
.A2(n_89),
.B1(n_183),
.B2(n_187),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_9),
.A2(n_89),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_9),
.A2(n_89),
.B1(n_418),
.B2(n_420),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_76),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_76),
.B1(n_156),
.B2(n_216),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_11),
.A2(n_231),
.B1(n_234),
.B2(n_237),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_11),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_250),
.C(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_11),
.B(n_138),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_11),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_11),
.B(n_83),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_11),
.B(n_188),
.Y(n_323)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_12),
.Y(n_385)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_14),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_14),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_15),
.A2(n_46),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_15),
.A2(n_46),
.B1(n_290),
.B2(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_16),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_221),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_219),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_200),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_20),
.B(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_119),
.C(n_166),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_21),
.A2(n_22),
.B1(n_119),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_84),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_23),
.A2(n_24),
.B(n_86),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B1(n_86),
.B2(n_118),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_24),
.A2(n_44),
.B1(n_118),
.B2(n_430),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_33),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_33),
.B1(n_169),
.B2(n_174),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_25),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_25),
.A2(n_237),
.B(n_257),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_25),
.A2(n_395),
.B1(n_396),
.B2(n_399),
.Y(n_394)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_26),
.B(n_260),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_26),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_26),
.A2(n_334),
.B1(n_364),
.B2(n_370),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_26),
.A2(n_400),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_28),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_29),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_31),
.A2(n_286),
.B(n_294),
.Y(n_285)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_37),
.Y(n_267)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_38),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g293 ( 
.A(n_38),
.Y(n_293)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_44),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_55),
.B1(n_75),
.B2(n_83),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_45),
.A2(n_55),
.B1(n_83),
.B2(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_47),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_48),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_48),
.Y(n_421)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_49),
.Y(n_141)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_49),
.Y(n_242)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_49),
.Y(n_315)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g138 ( 
.A1(n_53),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_55),
.A2(n_75),
.B1(n_83),
.B2(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_55),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_55),
.B(n_239),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_66),
.A2(n_160),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_66),
.A2(n_271),
.B(n_274),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_66),
.A2(n_211),
.B1(n_271),
.B2(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_66),
.A2(n_274),
.B(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_66),
.A2(n_211),
.B1(n_417),
.B2(n_434),
.Y(n_433)
);

AOI22x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_72),
.B(n_281),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_73),
.Y(n_369)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_79),
.Y(n_248)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_81),
.B(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_83),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_107),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g381 ( 
.A1(n_93),
.A2(n_382),
.A3(n_384),
.B1(n_386),
.B2(n_389),
.Y(n_381)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_95),
.B(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_95),
.Y(n_206)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_102),
.B2(n_105),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_106),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_107),
.A2(n_206),
.B(n_441),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_112),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_112),
.A2(n_389),
.B(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_119),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_157),
.B(n_165),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_158),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_138),
.B1(n_145),
.B2(n_153),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_122),
.A2(n_318),
.B(n_324),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_122),
.B(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_122),
.A2(n_138),
.B1(n_360),
.B2(n_443),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_122),
.A2(n_324),
.B(n_459),
.Y(n_458)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_146),
.B1(n_182),
.B2(n_190),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_123),
.A2(n_190),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_123),
.A2(n_190),
.B1(n_356),
.B2(n_411),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_129),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_132),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_132),
.Y(n_330)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_132),
.Y(n_388)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_137),
.Y(n_358)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_137),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_138),
.Y(n_190)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_141),
.Y(n_419)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_143),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_148),
.Y(n_321)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_148),
.Y(n_338)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_164),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_201),
.CI(n_202),
.CON(n_200),
.SN(n_200)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_166),
.B(n_445),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_181),
.C(n_191),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_167),
.B(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_168),
.B(n_177),
.Y(n_453)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_169),
.Y(n_436)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_173),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_174),
.A2(n_294),
.B(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_176),
.Y(n_301)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_178),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_181),
.B(n_191),
.Y(n_428)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_182),
.Y(n_443)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_186),
.Y(n_383)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_190),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_190),
.A2(n_356),
.B(n_359),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B(n_199),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_192),
.A2(n_193),
.B1(n_206),
.B2(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_200),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_209),
.B2(n_218),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_206),
.B(n_237),
.Y(n_362)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_217),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_230),
.B(n_238),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_211),
.A2(n_238),
.B(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI311xp33_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_424),
.A3(n_461),
.B1(n_479),
.C1(n_484),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_375),
.B(n_423),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_347),
.B(n_374),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_306),
.B(n_346),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_277),
.B(n_305),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_254),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_246),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_229),
.A2(n_246),
.B1(n_247),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_237),
.A2(n_319),
.B(n_322),
.Y(n_318)
);

HAxp5_ASAP7_75t_SL g389 ( 
.A(n_237),
.B(n_390),
.CON(n_389),
.SN(n_389)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_268),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_269),
.C(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_297),
.B(n_304),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_284),
.B(n_296),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_295),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_295),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_308),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_331),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_316),
.B2(n_317),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_316),
.C(n_331),
.Y(n_348)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI32xp33_ASAP7_75t_L g337 ( 
.A1(n_323),
.A2(n_338),
.A3(n_339),
.B1(n_342),
.B2(n_344),
.Y(n_337)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_337),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_348),
.B(n_349),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_354),
.B2(n_373),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_353),
.C(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_354),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_361),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_362),
.C(n_363),
.Y(n_402)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_376),
.B(n_377),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_405),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_378)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_393),
.B2(n_394),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_381),
.B(n_393),
.Y(n_457)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_402),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_409),
.B2(n_422),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_410),
.C(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_409),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_447),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_425),
.A2(n_447),
.B(n_480),
.C(n_483),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_444),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_444),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.C(n_431),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_429),
.CI(n_431),
.CON(n_460),
.SN(n_460)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_442),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_435),
.Y(n_469)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_440),
.B1(n_442),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_442),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_460),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_460),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_453),
.C(n_454),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_449),
.A2(n_450),
.B1(n_453),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.C(n_458),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_458),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_481),
.B(n_482),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_471),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_471),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.C(n_470),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_469),
.B1(n_470),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_470),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_476),
.Y(n_481)
);


endmodule