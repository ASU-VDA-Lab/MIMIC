module fake_netlist_5_397_n_1751 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1751);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1751;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_18),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_57),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_40),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_66),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_65),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_93),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_64),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_25),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_44),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx4_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_105),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_106),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_62),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_3),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_95),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_7),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_155),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_49),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_29),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_15),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_21),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_49),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_127),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_72),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_116),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_84),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_47),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_40),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_33),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_161),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_43),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_60),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_88),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_71),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_48),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_56),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_164),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_125),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_115),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_70),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_148),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_109),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_59),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_117),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_114),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_100),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_41),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_119),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_78),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_19),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_41),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_61),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_52),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_81),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_83),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_157),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_124),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_25),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_129),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_143),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_59),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_96),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_24),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_50),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_75),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_63),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_118),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_43),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_32),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_22),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_45),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_145),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_36),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_142),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_123),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_140),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_147),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_135),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_102),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_163),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_89),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_35),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_137),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_55),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_52),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_53),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_113),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_1),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_132),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_21),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_131),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_14),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_12),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_165),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_149),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_0),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_16),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_128),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_154),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_202),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_211),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_202),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_202),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_206),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_212),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_171),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_214),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_208),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_222),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_202),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_202),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_215),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_216),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_240),
.B(n_2),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_240),
.B(n_3),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_280),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_184),
.B(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_289),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_179),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_220),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_175),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_232),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_187),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_252),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_253),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_197),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_254),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_303),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_258),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_179),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_223),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_263),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_279),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_283),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_222),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_236),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_225),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_226),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

BUFx6f_ASAP7_75t_SL g394 ( 
.A(n_200),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_221),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_274),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_228),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_182),
.B(n_5),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_294),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_325),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_182),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_249),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_249),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_234),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_237),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_190),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_219),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_222),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_219),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_291),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_243),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_242),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_243),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_245),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_188),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_256),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_246),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_247),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_251),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_264),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_256),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_266),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_278),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_278),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_200),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_282),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_187),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_346),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_341),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_348),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_345),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_347),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_368),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_191),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_382),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_390),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_392),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_374),
.Y(n_455)
);

BUFx8_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_357),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_358),
.B(n_178),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_398),
.B(n_190),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_397),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_404),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_358),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_360),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_362),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_405),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_409),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_413),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_352),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_354),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_361),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_355),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_178),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_398),
.B(n_191),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_416),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_418),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_427),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_419),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_420),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_421),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_423),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_415),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_414),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_422),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_349),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_363),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_282),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_395),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_477),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_364),
.C(n_377),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_477),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_485),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_361),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_478),
.B(n_396),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_444),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_498),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_460),
.A2(n_483),
.B1(n_446),
.B2(n_455),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_411),
.B1(n_399),
.B2(n_396),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_434),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_426),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_459),
.B(n_426),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_359),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_457),
.B(n_370),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_457),
.B(n_399),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_446),
.Y(n_531)
);

BUFx8_ASAP7_75t_SL g532 ( 
.A(n_430),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_481),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_476),
.B(n_183),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_469),
.B(n_206),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_482),
.B(n_381),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_437),
.B(n_206),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_478),
.B(n_408),
.C(n_388),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_446),
.B(n_268),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_500),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_500),
.B(n_406),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_431),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_431),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_446),
.B(n_370),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_270),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_446),
.B(n_176),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_497),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_432),
.B(n_277),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_482),
.B(n_394),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_471),
.A2(n_394),
.B1(n_386),
.B2(n_393),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_481),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_497),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_438),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_469),
.B(n_206),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_444),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_447),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_497),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_445),
.B(n_206),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_471),
.A2(n_286),
.B1(n_186),
.B2(n_198),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_385),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_436),
.B(n_284),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_469),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_453),
.B(n_401),
.Y(n_570)
);

CKINVDCx6p67_ASAP7_75t_R g571 ( 
.A(n_435),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_495),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_475),
.A2(n_487),
.B1(n_490),
.B2(n_479),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_454),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_461),
.B(n_290),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_475),
.B(n_402),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_462),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_402),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_470),
.B(n_290),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_472),
.B(n_486),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_441),
.B(n_297),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_497),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_488),
.B(n_290),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_489),
.B(n_290),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_504),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_479),
.A2(n_290),
.B1(n_308),
.B2(n_384),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_458),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_473),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_492),
.B(n_403),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_487),
.B(n_308),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_494),
.B(n_403),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_433),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_456),
.B(n_308),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_449),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_450),
.B(n_311),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_474),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_450),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_456),
.A2(n_400),
.B1(n_379),
.B2(n_366),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_301),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_456),
.B(n_308),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_452),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_391),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_456),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_496),
.A2(n_505),
.B1(n_503),
.B2(n_502),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_463),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_502),
.B(n_257),
.Y(n_613)
);

OR2x2_ASAP7_75t_SL g614 ( 
.A(n_503),
.B(n_172),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_504),
.B(n_308),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_504),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_464),
.B(n_173),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_465),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_465),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_504),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_504),
.B(n_261),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_466),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_504),
.B(n_261),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_504),
.B(n_174),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_480),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_499),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_493),
.A2(n_391),
.B1(n_384),
.B2(n_383),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_493),
.B(n_371),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_439),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_439),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_467),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_439),
.B(n_177),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_480),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_440),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_491),
.B(n_331),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_440),
.Y(n_642)
);

INVxp33_ASAP7_75t_SL g643 ( 
.A(n_491),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_491),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_560),
.B(n_371),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_538),
.A2(n_180),
.B(n_192),
.C(n_196),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_499),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_520),
.B(n_523),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_499),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_528),
.B(n_440),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_629),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_519),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_512),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_639),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_567),
.B(n_285),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_506),
.A2(n_526),
.B1(n_538),
.B2(n_548),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_523),
.B(n_261),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_524),
.A2(n_181),
.B1(n_339),
.B2(n_338),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_524),
.B(n_261),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_514),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_529),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_545),
.B(n_285),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_510),
.B(n_181),
.Y(n_665)
);

AO22x1_ASAP7_75t_L g666 ( 
.A1(n_548),
.A2(n_203),
.B1(n_194),
.B2(n_193),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_510),
.B(n_443),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_506),
.A2(n_238),
.B1(n_321),
.B2(n_318),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_509),
.B(n_185),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_532),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_506),
.A2(n_295),
.B1(n_213),
.B2(n_205),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_508),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_544),
.B(n_285),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_555),
.A2(n_185),
.B1(n_189),
.B2(n_195),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_560),
.B(n_372),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_548),
.B(n_261),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_531),
.B(n_261),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_547),
.B(n_201),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_555),
.B(n_261),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_529),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_551),
.A2(n_641),
.B1(n_543),
.B2(n_549),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_574),
.B(n_189),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_593),
.B(n_255),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_612),
.B(n_265),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_534),
.B(n_296),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_506),
.A2(n_199),
.B1(n_339),
.B2(n_338),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_529),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_515),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_582),
.B(n_558),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_591),
.A2(n_224),
.B1(n_293),
.B2(n_235),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_506),
.A2(n_314),
.B1(n_204),
.B2(n_259),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_570),
.B(n_578),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_592),
.B(n_199),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_518),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_620),
.B(n_267),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_596),
.A2(n_530),
.B1(n_551),
.B2(n_507),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_536),
.B(n_269),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_557),
.B(n_204),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_540),
.B(n_259),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_637),
.B(n_271),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_542),
.A2(n_300),
.B1(n_292),
.B2(n_200),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_260),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_540),
.B(n_260),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_613),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_565),
.B(n_312),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_550),
.B(n_313),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_575),
.B(n_313),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_315),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_579),
.B(n_315),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_640),
.B(n_317),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_551),
.A2(n_302),
.B1(n_337),
.B2(n_336),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_579),
.B(n_319),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_589),
.B(n_329),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_585),
.B(n_329),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_595),
.B(n_332),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_610),
.B(n_372),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_609),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_333),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_333),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_600),
.B(n_373),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_551),
.A2(n_281),
.B1(n_210),
.B2(n_217),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_586),
.B(n_218),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_603),
.A2(n_327),
.B1(n_337),
.B2(n_336),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_641),
.B(n_373),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_641),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_640),
.B(n_327),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_566),
.A2(n_328),
.B1(n_335),
.B2(n_326),
.C(n_323),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_632),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_605),
.A2(n_383),
.B(n_380),
.C(n_378),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_580),
.B(n_296),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_580),
.B(n_296),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_608),
.B(n_375),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_586),
.B(n_229),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_617),
.B(n_375),
.Y(n_738)
);

AND2x6_ASAP7_75t_SL g739 ( 
.A(n_530),
.B(n_380),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_618),
.B(n_376),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_535),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_521),
.B(n_327),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_640),
.B(n_230),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_621),
.B(n_376),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_622),
.B(n_378),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_516),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_625),
.B(n_231),
.Y(n_747)
);

AND2x6_ASAP7_75t_SL g748 ( 
.A(n_641),
.B(n_365),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_562),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_633),
.B(n_233),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_614),
.A2(n_288),
.B1(n_239),
.B2(n_244),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_569),
.B(n_248),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_554),
.B(n_250),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_541),
.B(n_365),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_562),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_577),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_568),
.B(n_262),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_563),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_532),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_591),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_619),
.A2(n_369),
.B(n_207),
.C(n_328),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_581),
.B(n_272),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_633),
.B(n_273),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_601),
.B(n_275),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_602),
.B(n_193),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_599),
.B(n_276),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_572),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_599),
.B(n_287),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_513),
.B(n_517),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_572),
.B(n_74),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_584),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_627),
.A2(n_369),
.B(n_335),
.C(n_326),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_513),
.B(n_306),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_587),
.A2(n_310),
.B(n_299),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_522),
.B(n_304),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_513),
.B(n_305),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_606),
.B(n_323),
.Y(n_777)
);

INVx5_ASAP7_75t_L g778 ( 
.A(n_537),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_522),
.B(n_322),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_525),
.B(n_533),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_525),
.B(n_533),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_650),
.A2(n_587),
.B(n_533),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_694),
.B(n_577),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_651),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_653),
.B(n_571),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_669),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_669),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_648),
.A2(n_604),
.B1(n_627),
.B2(n_525),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_656),
.A2(n_648),
.B1(n_665),
.B2(n_698),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_669),
.B(n_630),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_706),
.B(n_194),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_SL g793 ( 
.A1(n_680),
.A2(n_657),
.B(n_660),
.C(n_646),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_651),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_665),
.A2(n_588),
.B1(n_611),
.B2(n_573),
.Y(n_795)
);

OAI321xp33_ASAP7_75t_L g796 ( 
.A1(n_730),
.A2(n_566),
.A3(n_638),
.B1(n_615),
.B2(n_316),
.C(n_203),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_753),
.A2(n_633),
.B1(n_635),
.B2(n_636),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_R g798 ( 
.A(n_671),
.B(n_316),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_667),
.B(n_598),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_616),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_734),
.B(n_633),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_652),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_753),
.A2(n_635),
.B1(n_634),
.B2(n_631),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_598),
.Y(n_804)
);

BUFx8_ASAP7_75t_L g805 ( 
.A(n_756),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_782),
.A2(n_553),
.B(n_556),
.Y(n_806)
);

BUFx4f_ASAP7_75t_L g807 ( 
.A(n_691),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_779),
.B(n_635),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_649),
.B(n_598),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_769),
.A2(n_552),
.B(n_556),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_657),
.A2(n_635),
.B1(n_566),
.B2(n_607),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_658),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_660),
.A2(n_615),
.B(n_624),
.C(n_626),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_682),
.A2(n_624),
.B1(n_626),
.B2(n_552),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_654),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_644),
.B(n_731),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_645),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_654),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_678),
.A2(n_564),
.B(n_623),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_735),
.B(n_616),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_661),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_720),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_779),
.B(n_583),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_677),
.A2(n_559),
.B(n_642),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_663),
.A2(n_689),
.B(n_681),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_673),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_695),
.B(n_594),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_695),
.B(n_594),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_701),
.B(n_594),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_766),
.A2(n_5),
.B(n_6),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_685),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_752),
.A2(n_776),
.B(n_773),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_691),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_759),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_696),
.B(n_561),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_770),
.B(n_561),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_645),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_645),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_676),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_696),
.B(n_561),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_691),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_670),
.B(n_7),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_705),
.A2(n_153),
.B1(n_151),
.B2(n_141),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_658),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_707),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_748),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_766),
.A2(n_112),
.B1(n_110),
.B2(n_108),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_757),
.A2(n_85),
.B(n_82),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_768),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_746),
.B(n_10),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_676),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_762),
.A2(n_12),
.B(n_15),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_768),
.A2(n_65),
.B(n_19),
.C(n_20),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_741),
.A2(n_17),
.B(n_23),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_SL g856 ( 
.A(n_749),
.B(n_17),
.Y(n_856)
);

INVx11_ASAP7_75t_L g857 ( 
.A(n_756),
.Y(n_857)
);

BUFx4f_ASAP7_75t_L g858 ( 
.A(n_719),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_749),
.B(n_23),
.Y(n_859)
);

OAI321xp33_ASAP7_75t_L g860 ( 
.A1(n_714),
.A2(n_24),
.A3(n_26),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_690),
.Y(n_861)
);

OAI21xp33_ASAP7_75t_L g862 ( 
.A1(n_659),
.A2(n_26),
.B(n_27),
.Y(n_862)
);

AOI21xp33_ASAP7_75t_L g863 ( 
.A1(n_725),
.A2(n_28),
.B(n_30),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_699),
.A2(n_31),
.B(n_34),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_775),
.B(n_31),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_764),
.A2(n_34),
.B(n_37),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_755),
.A2(n_37),
.B(n_39),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_725),
.A2(n_39),
.B(n_42),
.C(n_46),
.Y(n_868)
);

O2A1O1Ixp5_ASAP7_75t_L g869 ( 
.A1(n_699),
.A2(n_42),
.B(n_50),
.C(n_51),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_729),
.A2(n_51),
.B(n_53),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_676),
.B(n_54),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_728),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_729),
.A2(n_54),
.B(n_55),
.Y(n_873)
);

NOR2x1_ASAP7_75t_L g874 ( 
.A(n_707),
.B(n_56),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_750),
.A2(n_57),
.B(n_61),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_705),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_737),
.A2(n_715),
.B(n_717),
.C(n_711),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_710),
.A2(n_722),
.B1(n_715),
.B2(n_717),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_662),
.B(n_683),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_664),
.B(n_655),
.Y(n_880)
);

AND2x4_ASAP7_75t_SL g881 ( 
.A(n_767),
.B(n_727),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_737),
.A2(n_722),
.B1(n_710),
.B2(n_711),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_692),
.B(n_742),
.C(n_687),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_750),
.A2(n_763),
.B1(n_743),
.B2(n_697),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_758),
.A2(n_781),
.B(n_771),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_763),
.A2(n_684),
.B(n_686),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_772),
.A2(n_761),
.B(n_675),
.C(n_679),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_668),
.A2(n_672),
.B1(n_688),
.B2(n_693),
.Y(n_889)
);

AOI33xp33_ASAP7_75t_L g890 ( 
.A1(n_726),
.A2(n_733),
.A3(n_674),
.B1(n_703),
.B2(n_732),
.B3(n_666),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_727),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_747),
.A2(n_777),
.B(n_743),
.C(n_721),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_713),
.A2(n_702),
.B(n_744),
.C(n_745),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_723),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_736),
.B(n_738),
.Y(n_895)
);

OA22x2_ASAP7_75t_L g896 ( 
.A1(n_719),
.A2(n_700),
.B1(n_724),
.B2(n_751),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_704),
.A2(n_716),
.B(n_709),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_740),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_778),
.A2(n_718),
.B(n_708),
.Y(n_899)
);

CKINVDCx10_ASAP7_75t_R g900 ( 
.A(n_719),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_754),
.B(n_774),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_739),
.B(n_712),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_778),
.A2(n_650),
.B(n_780),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_778),
.A2(n_650),
.B(n_780),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_650),
.A2(n_782),
.B(n_780),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_648),
.A2(n_646),
.B(n_665),
.C(n_660),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_669),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_669),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_665),
.A2(n_648),
.B(n_768),
.C(n_766),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_678),
.A2(n_650),
.B(n_677),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_760),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_645),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_648),
.A2(n_646),
.B(n_665),
.C(n_660),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_692),
.B(n_478),
.C(n_485),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_678),
.A2(n_650),
.B(n_677),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_648),
.A2(n_656),
.B1(n_694),
.B2(n_523),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_653),
.B(n_512),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_669),
.B(n_512),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_648),
.A2(n_656),
.B1(n_694),
.B2(n_523),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_678),
.A2(n_650),
.B(n_677),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_669),
.B(n_512),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_653),
.B(n_512),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_656),
.A2(n_648),
.B1(n_665),
.B2(n_698),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_651),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_653),
.B(n_512),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_651),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_665),
.B(n_670),
.C(n_695),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_694),
.B(n_512),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_651),
.B(n_650),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_651),
.B(n_650),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_882),
.B(n_909),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_877),
.A2(n_843),
.B(n_927),
.C(n_878),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_815),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_928),
.B(n_917),
.Y(n_934)
);

O2A1O1Ixp5_ASAP7_75t_L g935 ( 
.A1(n_790),
.A2(n_923),
.B(n_887),
.C(n_901),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_906),
.A2(n_913),
.B(n_910),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_880),
.B(n_925),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_915),
.A2(n_920),
.B(n_892),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_894),
.B(n_898),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_929),
.A2(n_930),
.B(n_833),
.Y(n_940)
);

NAND2x1_ASAP7_75t_L g941 ( 
.A(n_787),
.B(n_788),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_799),
.A2(n_904),
.B(n_903),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_916),
.B(n_919),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_793),
.A2(n_783),
.B(n_819),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_802),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_862),
.A2(n_865),
.B(n_867),
.C(n_855),
.Y(n_946)
);

AOI21x1_ASAP7_75t_SL g947 ( 
.A1(n_828),
.A2(n_829),
.B(n_830),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_787),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_922),
.B(n_816),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_812),
.B(n_845),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_812),
.B(n_845),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_863),
.A2(n_860),
.B(n_795),
.C(n_850),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_885),
.B(n_897),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_895),
.B(n_824),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_822),
.B(n_895),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_818),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_821),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_808),
.B(n_785),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_813),
.A2(n_801),
.B(n_804),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_794),
.B(n_924),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_863),
.A2(n_854),
.B(n_868),
.C(n_888),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_809),
.A2(n_791),
.B(n_820),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_871),
.A2(n_796),
.B(n_890),
.C(n_873),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_893),
.A2(n_889),
.B(n_899),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_859),
.A2(n_831),
.B(n_864),
.C(n_837),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_789),
.B(n_883),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_797),
.A2(n_826),
.B(n_814),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_825),
.A2(n_841),
.B(n_836),
.Y(n_968)
);

NOR2x1_ASAP7_75t_SL g969 ( 
.A(n_787),
.B(n_788),
.Y(n_969)
);

NAND2x1_ASAP7_75t_L g970 ( 
.A(n_788),
.B(n_907),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_907),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_870),
.A2(n_851),
.B(n_875),
.C(n_866),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_907),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_811),
.A2(n_803),
.B(n_926),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_823),
.B(n_827),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_812),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_853),
.A2(n_869),
.B(n_902),
.C(n_876),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_832),
.A2(n_861),
.B1(n_896),
.B2(n_908),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_896),
.A2(n_908),
.B1(n_912),
.B2(n_817),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_784),
.B(n_792),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_918),
.A2(n_921),
.B(n_879),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_838),
.B(n_840),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_839),
.B(n_872),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_845),
.B(n_874),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_848),
.B(n_844),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_835),
.B(n_786),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_856),
.A2(n_858),
.A3(n_914),
.B(n_891),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_834),
.A2(n_842),
.B(n_891),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_884),
.B(n_891),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_SL g990 ( 
.A(n_846),
.B(n_807),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_881),
.B(n_911),
.Y(n_991)
);

AO31x2_ASAP7_75t_L g992 ( 
.A1(n_858),
.A2(n_884),
.A3(n_852),
.B(n_807),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_884),
.A2(n_900),
.B(n_857),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_798),
.B(n_847),
.Y(n_994)
);

AOI221x1_ASAP7_75t_L g995 ( 
.A1(n_805),
.A2(n_878),
.B1(n_877),
.B2(n_909),
.C(n_843),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_886),
.B(n_810),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_909),
.A2(n_877),
.B(n_927),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_802),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_894),
.B(n_898),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_894),
.B(n_898),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_928),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_882),
.B(n_909),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_835),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_882),
.B(n_909),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_882),
.A2(n_927),
.B(n_877),
.C(n_909),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_901),
.A2(n_886),
.B(n_905),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_909),
.A2(n_877),
.B(n_927),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_SL g1008 ( 
.A1(n_831),
.A2(n_867),
.B(n_855),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_790),
.A2(n_923),
.A3(n_909),
.B(n_877),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_878),
.A2(n_882),
.B1(n_927),
.B2(n_843),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_928),
.B(n_512),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_898),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_802),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_821),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_882),
.A2(n_877),
.B1(n_927),
.B2(n_909),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_787),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_928),
.B(n_512),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_886),
.A2(n_810),
.B(n_806),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_928),
.B(n_512),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_812),
.B(n_845),
.Y(n_1020)
);

AND3x4_ASAP7_75t_L g1021 ( 
.A(n_914),
.B(n_883),
.C(n_541),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_928),
.B(n_512),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_928),
.B(n_512),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_882),
.A2(n_909),
.B(n_877),
.C(n_843),
.Y(n_1024)
);

AND3x4_ASAP7_75t_L g1025 ( 
.A(n_914),
.B(n_883),
.C(n_541),
.Y(n_1025)
);

AO31x2_ASAP7_75t_L g1026 ( 
.A1(n_790),
.A2(n_923),
.A3(n_909),
.B(n_877),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_894),
.B(n_898),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_878),
.A2(n_877),
.B(n_909),
.C(n_927),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_787),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_894),
.B(n_898),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_787),
.Y(n_1031)
);

AOI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_927),
.A2(n_878),
.B(n_882),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_821),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_802),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_882),
.A2(n_909),
.B(n_877),
.C(n_843),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_787),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_886),
.A2(n_810),
.B(n_806),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_843),
.A2(n_730),
.B1(n_714),
.B2(n_878),
.C(n_796),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_928),
.B(n_512),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_882),
.B(n_909),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_886),
.A2(n_810),
.B(n_806),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_805),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_922),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_927),
.A2(n_878),
.B(n_882),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_802),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_894),
.B(n_898),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_882),
.A2(n_927),
.B(n_877),
.C(n_909),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_882),
.B(n_909),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_894),
.B(n_898),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_802),
.Y(n_1050)
);

INVxp67_ASAP7_75t_SL g1051 ( 
.A(n_800),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_894),
.B(n_898),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_909),
.A2(n_877),
.B(n_927),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_922),
.B(n_512),
.Y(n_1054)
);

AOI21x1_ASAP7_75t_L g1055 ( 
.A1(n_901),
.A2(n_886),
.B(n_905),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_971),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_1014),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1054),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_934),
.B(n_1011),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_1051),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_971),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1010),
.A2(n_954),
.B1(n_1024),
.B2(n_1035),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_945),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_998),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1013),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_SL g1066 ( 
.A(n_1038),
.B(n_1025),
.C(n_1021),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_971),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_934),
.B(n_1017),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_993),
.B(n_1033),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_955),
.B(n_949),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_950),
.B(n_951),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1034),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_950),
.B(n_951),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1032),
.A2(n_1044),
.B1(n_1040),
.B2(n_931),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1045),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_1003),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_1019),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_971),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_973),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1050),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1001),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_955),
.B(n_949),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1043),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1024),
.A2(n_1035),
.B1(n_932),
.B2(n_1047),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1001),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_1020),
.B(n_989),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_1020),
.B(n_984),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_936),
.A2(n_938),
.B(n_935),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_1042),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_973),
.B(n_1029),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1022),
.B(n_1023),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_973),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_937),
.B(n_939),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_976),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_976),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_975),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1021),
.A2(n_1025),
.B(n_980),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_960),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_933),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_956),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1039),
.B(n_999),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_SL g1103 ( 
.A1(n_985),
.A2(n_997),
.B(n_1007),
.C(n_1053),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_973),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1029),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1000),
.B(n_1012),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_L g1107 ( 
.A(n_1005),
.B(n_946),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_957),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1027),
.B(n_1030),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1110)
);

OAI22x1_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_931),
.B1(n_1002),
.B2(n_1004),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_976),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1029),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_983),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1052),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1029),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_1048),
.B1(n_1004),
.B2(n_1040),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_983),
.B(n_990),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_966),
.A2(n_1015),
.B1(n_1048),
.B2(n_986),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_976),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_948),
.B(n_1016),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_992),
.B(n_988),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_982),
.B(n_992),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_987),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_941),
.B(n_970),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_946),
.A2(n_952),
.B(n_1028),
.C(n_977),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_979),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_996),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_992),
.B(n_987),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_948),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1016),
.Y(n_1132)
);

INVx3_ASAP7_75t_SL g1133 ( 
.A(n_1031),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_958),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_943),
.B(n_952),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_982),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_963),
.B(n_1026),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_963),
.B(n_1026),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_1051),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_943),
.A2(n_974),
.B1(n_953),
.B2(n_977),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1031),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1008),
.A2(n_953),
.B1(n_964),
.B2(n_940),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_967),
.A2(n_1028),
.B1(n_981),
.B2(n_995),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_944),
.A2(n_942),
.A3(n_972),
.B(n_959),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_968),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_994),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1036),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_987),
.B(n_1026),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1036),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_969),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

INVx8_ASAP7_75t_L g1152 ( 
.A(n_987),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1009),
.B(n_1026),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_962),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1009),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_961),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_947),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_965),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1006),
.B(n_1055),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1018),
.A2(n_1037),
.B1(n_1041),
.B2(n_947),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_950),
.B(n_951),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_993),
.B(n_1014),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_932),
.A2(n_877),
.B(n_878),
.C(n_1044),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_950),
.B(n_951),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_934),
.B(n_1011),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1014),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1003),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1014),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_957),
.Y(n_1169)
);

OAI22x1_ASAP7_75t_L g1170 ( 
.A1(n_1010),
.A2(n_1025),
.B1(n_1021),
.B2(n_882),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_945),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_945),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_971),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1014),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_936),
.A2(n_938),
.B(n_935),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_945),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_934),
.B(n_1011),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_955),
.B(n_954),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_955),
.B(n_954),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1010),
.A2(n_882),
.B1(n_927),
.B2(n_954),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_971),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_945),
.Y(n_1182)
);

CKINVDCx6p67_ASAP7_75t_R g1183 ( 
.A(n_1042),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_976),
.B(n_787),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_934),
.B(n_1011),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_945),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_945),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_955),
.B(n_954),
.Y(n_1188)
);

INVx5_ASAP7_75t_L g1189 ( 
.A(n_971),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1054),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_945),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_950),
.B(n_951),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_934),
.B(n_927),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1155),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_1083),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1063),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1178),
.B(n_1179),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1077),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1170),
.B(n_1135),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1092),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1066),
.A2(n_1193),
.B1(n_1135),
.B2(n_1180),
.Y(n_1201)
);

BUFx8_ASAP7_75t_L g1202 ( 
.A(n_1168),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_SL g1203 ( 
.A1(n_1163),
.A2(n_1127),
.B(n_1119),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1064),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1077),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1167),
.Y(n_1206)
);

BUFx2_ASAP7_75t_R g1207 ( 
.A(n_1167),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1065),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

BUFx8_ASAP7_75t_SL g1210 ( 
.A(n_1090),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1193),
.A2(n_1107),
.B1(n_1085),
.B2(n_1062),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1076),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1188),
.A2(n_1098),
.B1(n_1190),
.B2(n_1162),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1071),
.B(n_1073),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1081),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1171),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1172),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1183),
.Y(n_1218)
);

AO21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1143),
.A2(n_1074),
.B(n_1117),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1057),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1107),
.A2(n_1074),
.B1(n_1111),
.B2(n_1165),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1176),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1069),
.A2(n_1162),
.B1(n_1090),
.B2(n_1146),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_1177),
.B1(n_1068),
.B2(n_1185),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1153),
.B(n_1137),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1140),
.A2(n_1117),
.B1(n_1156),
.B2(n_1128),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1148),
.B(n_1106),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1102),
.B(n_1110),
.Y(n_1228)
);

BUFx4f_ASAP7_75t_SL g1229 ( 
.A(n_1183),
.Y(n_1229)
);

INVx6_ASAP7_75t_L g1230 ( 
.A(n_1189),
.Y(n_1230)
);

INVx8_ASAP7_75t_L g1231 ( 
.A(n_1091),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1182),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1118),
.A2(n_1078),
.B1(n_1058),
.B2(n_1123),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1186),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1069),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1187),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1134),
.B(n_1099),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1166),
.Y(n_1238)
);

CKINVDCx6p67_ASAP7_75t_R g1239 ( 
.A(n_1169),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1122),
.B(n_1129),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1191),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1071),
.B(n_1073),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1100),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1101),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1097),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1082),
.Y(n_1246)
);

NOR2x1_ASAP7_75t_R g1247 ( 
.A(n_1057),
.B(n_1174),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1082),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1086),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1086),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1115),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1141),
.Y(n_1252)
);

AOI222xp33_ASAP7_75t_L g1253 ( 
.A1(n_1103),
.A2(n_1094),
.B1(n_1114),
.B2(n_1136),
.C1(n_1109),
.C2(n_1124),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1084),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1060),
.Y(n_1255)
);

INVx8_ASAP7_75t_L g1256 ( 
.A(n_1091),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1166),
.Y(n_1257)
);

AO21x1_ASAP7_75t_SL g1258 ( 
.A1(n_1143),
.A2(n_1158),
.B(n_1138),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1139),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1189),
.Y(n_1260)
);

INVx6_ASAP7_75t_L g1261 ( 
.A(n_1189),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1174),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1147),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1073),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1147),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1056),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1069),
.A2(n_1162),
.B1(n_1175),
.B2(n_1089),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1103),
.B(n_1192),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1108),
.A2(n_1075),
.B1(n_1088),
.B2(n_1087),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1160),
.A2(n_1159),
.B(n_1145),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1152),
.A2(n_1089),
.B1(n_1175),
.B2(n_1075),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1144),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1056),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1125),
.B(n_1130),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1144),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1079),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1079),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1159),
.A2(n_1151),
.B(n_1125),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1157),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1189),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1157),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1125),
.Y(n_1283)
);

INVx3_ASAP7_75t_SL g1284 ( 
.A(n_1161),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1080),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1161),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1142),
.A2(n_1126),
.B(n_1150),
.Y(n_1287)
);

AO21x1_ASAP7_75t_L g1288 ( 
.A1(n_1157),
.A2(n_1130),
.B(n_1122),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1161),
.B(n_1192),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1154),
.A2(n_1130),
.B(n_1152),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1126),
.A2(n_1184),
.B(n_1104),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1152),
.A2(n_1088),
.B1(n_1087),
.B2(n_1164),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1184),
.A2(n_1173),
.B(n_1120),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1173),
.A2(n_1120),
.B(n_1121),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1088),
.A2(n_1087),
.B1(n_1133),
.B2(n_1164),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1080),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1112),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1061),
.A2(n_1067),
.B(n_1113),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1113),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1095),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1131),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1091),
.A2(n_1132),
.B1(n_1120),
.B2(n_1095),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1091),
.A2(n_1149),
.B1(n_1131),
.B2(n_1096),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1091),
.Y(n_1304)
);

BUFx2_ASAP7_75t_SL g1305 ( 
.A(n_1113),
.Y(n_1305)
);

INVx8_ASAP7_75t_L g1306 ( 
.A(n_1080),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1093),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1093),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1093),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1194),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_1105),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1225),
.B(n_1116),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1199),
.B(n_1116),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1279),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1246),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1199),
.B(n_1181),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1201),
.A2(n_1211),
.B1(n_1213),
.B2(n_1221),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1235),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1290),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1227),
.B(n_1258),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1278),
.B(n_1274),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1240),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1227),
.B(n_1258),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1290),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1280),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1268),
.B(n_1272),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1275),
.B(n_1219),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1235),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1248),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1203),
.A2(n_1219),
.B1(n_1253),
.B2(n_1200),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1282),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1203),
.A2(n_1226),
.B1(n_1195),
.B2(n_1224),
.Y(n_1332)
);

BUFx8_ASAP7_75t_SL g1333 ( 
.A(n_1210),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1240),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1290),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1240),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1274),
.B(n_1283),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1287),
.B(n_1267),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1288),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1287),
.B(n_1283),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1197),
.A2(n_1228),
.B(n_1237),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1288),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1232),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1233),
.A2(n_1223),
.B1(n_1269),
.B2(n_1237),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1249),
.B(n_1250),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1270),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1270),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1232),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1234),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1239),
.Y(n_1350)
);

INVxp33_ASAP7_75t_L g1351 ( 
.A(n_1254),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1234),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1245),
.A2(n_1251),
.B(n_1259),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1291),
.A2(n_1294),
.B(n_1293),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1289),
.B(n_1198),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1231),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1271),
.B(n_1241),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1196),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1255),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1204),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1304),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1295),
.A2(n_1298),
.B(n_1244),
.Y(n_1363)
);

INVx8_ASAP7_75t_L g1364 ( 
.A(n_1231),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1208),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1209),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1230),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1212),
.A2(n_1215),
.B(n_1216),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1304),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1217),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1222),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1252),
.B(n_1243),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1266),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1263),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1239),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1277),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1214),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1303),
.A2(n_1265),
.B(n_1292),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1310),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1341),
.B(n_1297),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1336),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1317),
.A2(n_1309),
.B1(n_1307),
.B2(n_1302),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1333),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1341),
.B(n_1262),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1340),
.B(n_1308),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1315),
.B(n_1262),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1360),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1355),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1317),
.A2(n_1260),
.B(n_1281),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1324),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1323),
.B(n_1301),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1326),
.B(n_1220),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1358),
.B(n_1301),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1368),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1369),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1368),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1368),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1358),
.B(n_1242),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1358),
.B(n_1242),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1374),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1348),
.B(n_1300),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1311),
.B(n_1242),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1374),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1368),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1325),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1326),
.B(n_1220),
.Y(n_1409)
);

NAND2x1_ASAP7_75t_L g1410 ( 
.A(n_1324),
.B(n_1261),
.Y(n_1410)
);

OAI321xp33_ASAP7_75t_L g1411 ( 
.A1(n_1330),
.A2(n_1332),
.A3(n_1344),
.B1(n_1380),
.B2(n_1363),
.C(n_1353),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1312),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1332),
.A2(n_1286),
.B1(n_1218),
.B2(n_1264),
.C(n_1198),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1354),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1369),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1330),
.A2(n_1286),
.B1(n_1284),
.B2(n_1264),
.C(n_1218),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1345),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1348),
.B(n_1299),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1339),
.A2(n_1305),
.B(n_1256),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1312),
.B(n_1285),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1312),
.B(n_1285),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1314),
.B(n_1284),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1315),
.B(n_1202),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1319),
.B(n_1299),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1337),
.B(n_1313),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1324),
.B(n_1335),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1372),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1337),
.B(n_1285),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1324),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1316),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_1411),
.B(n_1363),
.C(n_1380),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1382),
.B(n_1329),
.Y(n_1432)
);

OA211x2_ASAP7_75t_L g1433 ( 
.A1(n_1410),
.A2(n_1353),
.B(n_1350),
.C(n_1376),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1344),
.C(n_1329),
.D(n_1345),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1391),
.B(n_1318),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1423),
.B(n_1318),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1416),
.A2(n_1328),
.B1(n_1318),
.B2(n_1351),
.C(n_1316),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1430),
.B(n_1370),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1411),
.B(n_1324),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1392),
.A2(n_1328),
.B1(n_1376),
.B2(n_1350),
.C(n_1342),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1417),
.B(n_1370),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1386),
.B(n_1370),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1384),
.A2(n_1338),
.B(n_1327),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1392),
.A2(n_1384),
.B(n_1388),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1390),
.B(n_1425),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1395),
.B(n_1324),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1395),
.B(n_1328),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1396),
.A2(n_1365),
.B1(n_1366),
.B2(n_1359),
.C(n_1361),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1409),
.B(n_1371),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1396),
.A2(n_1365),
.B1(n_1366),
.B2(n_1359),
.C(n_1361),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1409),
.B(n_1371),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1401),
.A2(n_1350),
.B1(n_1376),
.B2(n_1207),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1425),
.B(n_1340),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1371),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1397),
.B(n_1342),
.C(n_1339),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1385),
.A2(n_1205),
.B1(n_1206),
.B2(n_1229),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1381),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1403),
.B(n_1343),
.Y(n_1458)
);

NAND4xp25_ASAP7_75t_L g1459 ( 
.A(n_1404),
.B(n_1372),
.C(n_1313),
.D(n_1343),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1410),
.A2(n_1367),
.B1(n_1379),
.B2(n_1322),
.C(n_1334),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1397),
.B(n_1202),
.C(n_1331),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1420),
.B(n_1352),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1387),
.B(n_1340),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1406),
.A2(n_1372),
.B1(n_1313),
.B2(n_1357),
.C(n_1319),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1421),
.B(n_1357),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1401),
.A2(n_1356),
.B1(n_1379),
.B2(n_1362),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1387),
.B(n_1340),
.Y(n_1467)
);

OAI211xp5_ASAP7_75t_L g1468 ( 
.A1(n_1404),
.A2(n_1346),
.B(n_1378),
.C(n_1377),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1399),
.B(n_1202),
.C(n_1346),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1399),
.B(n_1407),
.C(n_1400),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1393),
.B(n_1324),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1387),
.B(n_1335),
.Y(n_1472)
);

OAI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1422),
.A2(n_1367),
.B1(n_1379),
.B2(n_1322),
.C(n_1334),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1387),
.B(n_1335),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1402),
.A2(n_1356),
.B1(n_1379),
.B2(n_1362),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1402),
.A2(n_1379),
.B1(n_1327),
.B2(n_1338),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1426),
.A2(n_1327),
.B1(n_1362),
.B2(n_1367),
.C(n_1347),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1427),
.B(n_1428),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1427),
.B(n_1335),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1418),
.B(n_1373),
.C(n_1377),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1405),
.B(n_1348),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1393),
.B(n_1335),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1419),
.B(n_1335),
.Y(n_1483)
);

AND2x2_ASAP7_75t_SL g1484 ( 
.A(n_1419),
.B(n_1335),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1405),
.B(n_1349),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1426),
.A2(n_1347),
.B1(n_1378),
.B2(n_1375),
.C(n_1373),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1479),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1457),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1426),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1441),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1431),
.A2(n_1338),
.B1(n_1321),
.B2(n_1394),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1432),
.B(n_1428),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1442),
.B(n_1400),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1445),
.B(n_1426),
.Y(n_1495)
);

BUFx5_ASAP7_75t_L g1496 ( 
.A(n_1483),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1438),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1454),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1470),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1483),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1449),
.B(n_1398),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1451),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1462),
.B(n_1398),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1446),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1453),
.B(n_1472),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1465),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1484),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1393),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1471),
.B(n_1393),
.Y(n_1509)
);

NAND2x1_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1419),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_1429),
.Y(n_1512)
);

AND2x4_ASAP7_75t_SL g1513 ( 
.A(n_1476),
.B(n_1322),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1446),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1481),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1435),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1485),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1463),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1467),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1482),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1447),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1478),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1459),
.B(n_1415),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1455),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1520),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1520),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1488),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1488),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1520),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1407),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1498),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1511),
.B(n_1482),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1429),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1448),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1497),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_1429),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1500),
.B(n_1429),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1496),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1507),
.Y(n_1540)
);

AOI32xp33_ASAP7_75t_L g1541 ( 
.A1(n_1524),
.A2(n_1444),
.A3(n_1439),
.B1(n_1452),
.B2(n_1437),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1494),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1500),
.B(n_1419),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1524),
.B(n_1450),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1507),
.B(n_1496),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1516),
.A2(n_1439),
.B1(n_1434),
.B2(n_1436),
.Y(n_1547)
);

AO22x1_ASAP7_75t_L g1548 ( 
.A1(n_1507),
.A2(n_1356),
.B1(n_1433),
.B2(n_1440),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1494),
.B(n_1486),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1509),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1504),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1424),
.Y(n_1552)
);

AOI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1523),
.A2(n_1443),
.B(n_1469),
.C(n_1461),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1492),
.B(n_1464),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1492),
.B(n_1468),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1490),
.Y(n_1556)
);

NAND2x1_ASAP7_75t_SL g1557 ( 
.A(n_1514),
.B(n_1389),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1496),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1506),
.B(n_1408),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_R g1560 ( 
.A(n_1509),
.B(n_1383),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1501),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1496),
.B(n_1414),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1496),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1522),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1496),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1527),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1528),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1528),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1545),
.B(n_1521),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1525),
.Y(n_1571)
);

INVxp33_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1506),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1541),
.B(n_1496),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1559),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1559),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

CKINVDCx16_ASAP7_75t_R g1578 ( 
.A(n_1560),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1546),
.B(n_1518),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1534),
.B(n_1510),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1546),
.B(n_1518),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1556),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1532),
.B(n_1496),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1502),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1547),
.B(n_1502),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1515),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1554),
.B(n_1515),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1541),
.B(n_1517),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1553),
.A2(n_1513),
.B1(n_1475),
.B2(n_1466),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1531),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1549),
.B(n_1561),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1525),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1531),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1535),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1555),
.B(n_1503),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1519),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_SL g1601 ( 
.A(n_1557),
.B(n_1510),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1540),
.B(n_1460),
.Y(n_1602)
);

NOR2x1p5_ASAP7_75t_L g1603 ( 
.A(n_1540),
.B(n_1205),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1540),
.B(n_1509),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1540),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1550),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1553),
.B(n_1561),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1535),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1594),
.B(n_1530),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1550),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1605),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1606),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1574),
.B(n_1532),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1578),
.A2(n_1491),
.B1(n_1477),
.B2(n_1513),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1599),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1604),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1572),
.B(n_1536),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1572),
.B(n_1536),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1569),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1583),
.B(n_1530),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1607),
.B(n_1542),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_1210),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1574),
.B(n_1532),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1586),
.A2(n_1565),
.B1(n_1539),
.B2(n_1563),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1573),
.B(n_1542),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1602),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1579),
.B(n_1533),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1588),
.B(n_1589),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1580),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1598),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1581),
.B(n_1533),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1604),
.A2(n_1557),
.B(n_1539),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1571),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1613),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1633),
.B(n_1456),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1600),
.Y(n_1650)
);

AOI222xp33_ASAP7_75t_L g1651 ( 
.A1(n_1617),
.A2(n_1601),
.B1(n_1577),
.B2(n_1582),
.C1(n_1548),
.C2(n_1585),
.Y(n_1651)
);

AND4x1_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1591),
.C(n_1581),
.D(n_1585),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1601),
.C(n_1605),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1612),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1614),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1618),
.A2(n_1584),
.B1(n_1548),
.B2(n_1596),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1610),
.B(n_1575),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1610),
.B(n_1625),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1640),
.B(n_1584),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1615),
.Y(n_1664)
);

OAI32xp33_ASAP7_75t_L g1665 ( 
.A1(n_1638),
.A2(n_1560),
.A3(n_1539),
.B1(n_1565),
.B2(n_1563),
.Y(n_1665)
);

AOI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1627),
.A2(n_1576),
.B(n_1563),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1614),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1640),
.B(n_1558),
.Y(n_1668)
);

OAI31xp33_ASAP7_75t_L g1669 ( 
.A1(n_1611),
.A2(n_1637),
.A3(n_1620),
.B(n_1634),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1611),
.A2(n_1558),
.B1(n_1565),
.B2(n_1562),
.Y(n_1670)
);

CKINVDCx14_ASAP7_75t_R g1671 ( 
.A(n_1636),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1661),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1671),
.B(n_1622),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1649),
.B(n_1656),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1648),
.A2(n_1611),
.B1(n_1634),
.B2(n_1620),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1632),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1660),
.A2(n_1651),
.B1(n_1669),
.B2(n_1646),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1664),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1654),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1658),
.A2(n_1620),
.B1(n_1631),
.B2(n_1625),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1664),
.B(n_1609),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1653),
.B(n_1626),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1652),
.A2(n_1624),
.B(n_1558),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1655),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1650),
.A2(n_1626),
.B1(n_1643),
.B2(n_1630),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1655),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1678),
.B(n_1662),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1692),
.B(n_1662),
.Y(n_1695)
);

NAND4xp75_ASAP7_75t_L g1696 ( 
.A(n_1688),
.B(n_1667),
.C(n_1657),
.D(n_1663),
.Y(n_1696)
);

AOI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1684),
.A2(n_1665),
.B(n_1657),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1689),
.A2(n_1670),
.B1(n_1666),
.B2(n_1659),
.C(n_1667),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1680),
.A2(n_1659),
.B(n_1665),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1675),
.B(n_1206),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1680),
.A2(n_1643),
.B1(n_1630),
.B2(n_1639),
.C(n_1642),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1684),
.A2(n_1641),
.B(n_1642),
.C(n_1639),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1679),
.A2(n_1668),
.B1(n_1641),
.B2(n_1644),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1672),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1673),
.Y(n_1705)
);

OAI31xp33_ASAP7_75t_L g1706 ( 
.A1(n_1686),
.A2(n_1668),
.A3(n_1644),
.B(n_1562),
.Y(n_1706)
);

NOR3xp33_ASAP7_75t_L g1707 ( 
.A(n_1700),
.B(n_1676),
.C(n_1682),
.Y(n_1707)
);

NOR3x1_ASAP7_75t_L g1708 ( 
.A(n_1696),
.B(n_1677),
.C(n_1687),
.Y(n_1708)
);

AND2x2_ASAP7_75t_SL g1709 ( 
.A(n_1704),
.B(n_1679),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1697),
.B(n_1691),
.C(n_1681),
.Y(n_1710)
);

OAI322xp33_ASAP7_75t_L g1711 ( 
.A1(n_1701),
.A2(n_1685),
.A3(n_1683),
.B1(n_1674),
.B2(n_1691),
.C1(n_1595),
.C2(n_1571),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1694),
.Y(n_1712)
);

NOR4xp75_ASAP7_75t_L g1713 ( 
.A(n_1693),
.B(n_1533),
.C(n_1562),
.D(n_1537),
.Y(n_1713)
);

OAI322xp33_ASAP7_75t_L g1714 ( 
.A1(n_1698),
.A2(n_1595),
.A3(n_1552),
.B1(n_1529),
.B2(n_1525),
.C1(n_1526),
.C2(n_1543),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_L g1715 ( 
.A(n_1699),
.B(n_1247),
.C(n_1526),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1529),
.C(n_1526),
.Y(n_1716)
);

NOR4xp25_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1529),
.C(n_1552),
.D(n_1544),
.Y(n_1717)
);

NAND4xp25_ASAP7_75t_SL g1718 ( 
.A(n_1710),
.B(n_1702),
.C(n_1706),
.D(n_1703),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1711),
.B(n_1695),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1707),
.A2(n_1552),
.B(n_1544),
.C(n_1538),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1505),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1716),
.B(n_1543),
.C(n_1544),
.Y(n_1722)
);

NOR4xp25_ASAP7_75t_L g1723 ( 
.A(n_1712),
.B(n_1538),
.C(n_1537),
.D(n_1564),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1721),
.Y(n_1724)
);

AO22x2_ASAP7_75t_L g1725 ( 
.A1(n_1718),
.A2(n_1715),
.B1(n_1708),
.B2(n_1713),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_L g1726 ( 
.A(n_1719),
.B(n_1714),
.Y(n_1726)
);

NOR2x2_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1717),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1537),
.B1(n_1538),
.B2(n_1238),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1722),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1721),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1724),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1730),
.B(n_1729),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1726),
.A2(n_1564),
.B(n_1493),
.Y(n_1733)
);

NAND4xp75_ASAP7_75t_L g1734 ( 
.A(n_1728),
.B(n_1489),
.C(n_1495),
.D(n_1238),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1725),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1727),
.A2(n_1257),
.B1(n_1509),
.B2(n_1512),
.Y(n_1736)
);

XNOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1735),
.B(n_1257),
.Y(n_1737)
);

AND4x1_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1489),
.C(n_1495),
.D(n_1508),
.Y(n_1738)
);

XOR2xp5_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1307),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1737),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1740),
.Y(n_1741)
);

OAI22x1_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1731),
.B1(n_1739),
.B2(n_1736),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1733),
.B1(n_1738),
.B2(n_1487),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1487),
.B(n_1503),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1742),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1306),
.B(n_1364),
.Y(n_1746)
);

AO21x2_ASAP7_75t_L g1747 ( 
.A1(n_1744),
.A2(n_1512),
.B(n_1522),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1306),
.B(n_1281),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1747),
.B1(n_1512),
.B2(n_1306),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_R g1750 ( 
.A1(n_1749),
.A2(n_1306),
.B1(n_1309),
.B2(n_1256),
.C(n_1231),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1260),
.B(n_1473),
.C(n_1296),
.Y(n_1751)
);


endmodule