module fake_jpeg_3067_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_20),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AND2x6_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_2),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.C(n_7),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_8),
.A2(n_3),
.B(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_8),
.B1(n_14),
.B2(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_33),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_9),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_34),
.C(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_25),
.C(n_7),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_26),
.C(n_9),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_39),
.B(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_14),
.C(n_16),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.C(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_16),
.C(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_34),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_27),
.B(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_36),
.C(n_38),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_49),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_51),
.B(n_46),
.Y(n_53)
);


endmodule