module real_jpeg_14465_n_16 (n_5, n_4, n_8, n_0, n_12, n_324, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_324;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_31),
.B1(n_35),
.B2(n_48),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_3),
.A2(n_48),
.B1(n_75),
.B2(n_76),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_4),
.A2(n_75),
.B1(n_76),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_136),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_136),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_31),
.B1(n_35),
.B2(n_136),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_75),
.B1(n_76),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_83),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_6),
.A2(n_31),
.B1(n_35),
.B2(n_83),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_75),
.B1(n_76),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_159),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_159),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_7),
.A2(n_31),
.B1(n_35),
.B2(n_159),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_31),
.B1(n_35),
.B2(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_10),
.A2(n_57),
.B1(n_75),
.B2(n_76),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_31),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_39),
.B1(n_75),
.B2(n_76),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_74),
.B(n_75),
.C(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_75),
.B1(n_76),
.B2(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_13),
.B(n_85),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_150),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_103),
.B1(n_104),
.B2(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_13),
.B(n_91),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_14),
.A2(n_34),
.B1(n_75),
.B2(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_14),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_14),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_132)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_316),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_308),
.B(n_315),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_274),
.B(n_305),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_137),
.B(n_273),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_117),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_21),
.B(n_117),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_87),
.B2(n_116),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_22),
.B(n_88),
.C(n_100),
.Y(n_303)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_58),
.C(n_70),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_24),
.A2(n_25),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_28),
.A2(n_103),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_29),
.A2(n_40),
.B1(n_127),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_29),
.A2(n_40),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_30),
.A2(n_40),
.B(n_129),
.Y(n_203)
);

CKINVDCx6p67_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_35),
.B(n_52),
.C(n_150),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_35),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_36),
.A2(n_104),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_38),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_44),
.A2(n_54),
.B(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_45),
.A2(n_60),
.B(n_200),
.C(n_202),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_45),
.B(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_46),
.B(n_61),
.C(n_63),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_49),
.A2(n_56),
.B(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_49),
.A2(n_95),
.B(n_108),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_49),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_49),
.A2(n_55),
.B1(n_207),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_49),
.A2(n_55),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_49),
.A2(n_55),
.B1(n_215),
.B2(n_225),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_49),
.A2(n_55),
.B(n_95),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_54),
.B(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_70),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_65),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_59),
.A2(n_154),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_64),
.B1(n_74),
.B2(n_79),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_79),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_64),
.B(n_150),
.CON(n_201),
.SN(n_201)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_65),
.B(n_155),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_66),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_66),
.A2(n_91),
.B1(n_153),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_66),
.A2(n_91),
.B1(n_188),
.B2(n_201),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_66),
.A2(n_91),
.B(n_132),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_81),
.B(n_84),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_71),
.A2(n_80),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_71),
.A2(n_114),
.B(n_312),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_82),
.B1(n_85),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_85),
.B1(n_158),
.B2(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_72),
.B(n_115),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_72),
.A2(n_85),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_73)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_80),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_84),
.B(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_100),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_99),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_92),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_94),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_99),
.B(n_277),
.C(n_290),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_99),
.B(n_277),
.CI(n_290),
.CON(n_304),
.SN(n_304)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_101),
.A2(n_102),
.B(n_111),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_103),
.A2(n_104),
.B1(n_230),
.B2(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_104),
.B(n_150),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_123),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_122),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_123),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_134),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_130),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_133),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_267),
.B(n_272),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_176),
.B1(n_192),
.B2(n_266),
.C(n_324),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_140),
.B(n_165),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_161),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_141),
.B(n_162),
.C(n_163),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_151),
.C(n_156),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_143),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_154),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_175),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_175),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_177),
.B(n_190),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_178),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_182),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_265),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_260),
.B(n_264),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_216),
.B(n_259),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_211),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_211),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_204),
.C(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_203),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_214),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_254),
.B(n_258),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_244),
.B(n_253),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_233),
.B(n_243),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_226),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_242),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_249),
.C(n_252),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_302),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_291),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_291),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_289),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_285),
.C(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_285),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_295),
.C(n_300),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_289),
.B1(n_294),
.B2(n_301),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_292),
.C(n_301),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_297),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_314),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_319),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.CI(n_313),
.CON(n_309),
.SN(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);


endmodule