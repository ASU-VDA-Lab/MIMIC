module real_aes_2119_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_830, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_830;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g216 ( .A(n_0), .B(n_153), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_1), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_3), .B(n_129), .Y(n_174) );
NAND2xp33_ASAP7_75t_SL g236 ( .A(n_4), .B(n_135), .Y(n_236) );
INVx1_ASAP7_75t_L g228 ( .A(n_5), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_6), .B(n_179), .Y(n_452) );
INVx1_ASAP7_75t_L g496 ( .A(n_7), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_8), .Y(n_827) );
AND2x2_ASAP7_75t_L g172 ( .A(n_9), .B(n_158), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_10), .Y(n_488) );
INVx2_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_12), .Y(n_437) );
INVx1_ASAP7_75t_L g461 ( .A(n_13), .Y(n_461) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_14), .A2(n_137), .B1(n_232), .B2(n_234), .C(n_235), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_15), .B(n_129), .Y(n_196) );
INVx1_ASAP7_75t_L g441 ( .A(n_16), .Y(n_441) );
NOR2xp33_ASAP7_75t_SL g824 ( .A(n_16), .B(n_442), .Y(n_824) );
INVx1_ASAP7_75t_L g459 ( .A(n_17), .Y(n_459) );
INVx1_ASAP7_75t_SL g555 ( .A(n_18), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_19), .B(n_130), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_20), .A2(n_137), .B(n_176), .Y(n_175) );
AOI221xp5_ASAP7_75t_SL g205 ( .A1(n_21), .A2(n_38), .B1(n_129), .B2(n_137), .C(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_22), .B(n_153), .Y(n_177) );
AOI33xp33_ASAP7_75t_L g505 ( .A1(n_23), .A2(n_50), .A3(n_122), .B1(n_142), .B2(n_506), .B3(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g482 ( .A(n_24), .Y(n_482) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_26), .A2(n_89), .B(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g159 ( .A(n_26), .B(n_89), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_27), .B(n_151), .Y(n_200) );
INVxp67_ASAP7_75t_L g230 ( .A(n_28), .Y(n_230) );
AND2x2_ASAP7_75t_L g169 ( .A(n_29), .B(n_157), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_30), .B(n_120), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_31), .A2(n_137), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_32), .B(n_151), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_33), .A2(n_49), .B1(n_641), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_33), .Y(n_816) );
AND2x2_ASAP7_75t_L g127 ( .A(n_34), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g135 ( .A(n_34), .B(n_125), .Y(n_135) );
INVx1_ASAP7_75t_L g141 ( .A(n_34), .Y(n_141) );
OR2x6_ASAP7_75t_L g439 ( .A(n_35), .B(n_440), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g825 ( .A(n_35), .B(n_437), .C(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_36), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_37), .B(n_120), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_39), .A2(n_179), .B1(n_212), .B2(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_40), .B(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_41), .A2(n_80), .B1(n_137), .B2(n_139), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_42), .B(n_130), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_43), .B(n_153), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_44), .B(n_115), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_45), .B(n_130), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_46), .Y(n_526) );
AND2x2_ASAP7_75t_L g219 ( .A(n_47), .B(n_157), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_48), .B(n_157), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_49), .Y(n_641) );
HB1xp67_ASAP7_75t_SL g712 ( .A(n_49), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_51), .B(n_130), .Y(n_474) );
INVx1_ASAP7_75t_L g123 ( .A(n_52), .Y(n_123) );
INVx1_ASAP7_75t_L g132 ( .A(n_52), .Y(n_132) );
AND2x2_ASAP7_75t_L g475 ( .A(n_53), .B(n_157), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_54), .A2(n_73), .B1(n_120), .B2(n_139), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_55), .B(n_120), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_56), .B(n_129), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_57), .B(n_212), .Y(n_490) );
AOI21xp5_ASAP7_75t_SL g515 ( .A1(n_58), .A2(n_139), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g160 ( .A(n_59), .B(n_157), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_60), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_61), .B(n_151), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_62), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_63), .B(n_158), .Y(n_201) );
INVx1_ASAP7_75t_L g455 ( .A(n_64), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_65), .A2(n_137), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g473 ( .A(n_66), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_67), .B(n_151), .Y(n_178) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_68), .B(n_115), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_69), .A2(n_139), .B(n_472), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_70), .A2(n_101), .B1(n_821), .B2(n_828), .Y(n_100) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_71), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_72), .B(n_120), .Y(n_508) );
AND2x2_ASAP7_75t_L g557 ( .A(n_74), .B(n_234), .Y(n_557) );
INVx1_ASAP7_75t_L g457 ( .A(n_75), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_76), .A2(n_139), .B(n_554), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_77), .A2(n_114), .B(n_139), .C(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_78), .A2(n_83), .B1(n_120), .B2(n_129), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_79), .B(n_129), .Y(n_155) );
INVx1_ASAP7_75t_L g442 ( .A(n_81), .Y(n_442) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_82), .B(n_234), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_84), .A2(n_139), .B1(n_503), .B2(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_85), .B(n_153), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_86), .B(n_153), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_87), .A2(n_103), .B1(n_790), .B2(n_794), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_88), .A2(n_137), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g517 ( .A(n_90), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_91), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g509 ( .A(n_92), .B(n_234), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_93), .A2(n_480), .B(n_481), .C(n_483), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_94), .B(n_129), .Y(n_218) );
INVxp67_ASAP7_75t_L g233 ( .A(n_95), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_96), .B(n_151), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_97), .A2(n_137), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_98), .B(n_799), .Y(n_798) );
BUFx2_ASAP7_75t_SL g808 ( .A(n_98), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_99), .B(n_130), .Y(n_518) );
OA21x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_798), .B(n_804), .Y(n_101) );
OAI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_104), .B(n_789), .Y(n_102) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_436), .B1(n_443), .B2(n_785), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_107), .A2(n_444), .B1(n_791), .B2(n_792), .Y(n_790) );
AND3x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_307), .C(n_381), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_249), .C(n_280), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_182), .B(n_191), .C(n_220), .Y(n_109) );
AOI21x1_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_161), .B(n_180), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_111), .A2(n_283), .B1(n_289), .B2(n_292), .Y(n_282) );
AND2x2_ASAP7_75t_L g416 ( .A(n_111), .B(n_184), .Y(n_416) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_145), .Y(n_111) );
BUFx2_ASAP7_75t_L g187 ( .A(n_112), .Y(n_187) );
AND2x2_ASAP7_75t_L g275 ( .A(n_112), .B(n_146), .Y(n_275) );
AND2x2_ASAP7_75t_L g346 ( .A(n_112), .B(n_190), .Y(n_346) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_113), .Y(n_240) );
AOI21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_144), .Y(n_113) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_114), .A2(n_501), .B(n_509), .Y(n_500) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_114), .A2(n_501), .B(n_509), .Y(n_572) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_115), .A2(n_196), .B(n_197), .Y(n_195) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_115), .A2(n_494), .B(n_498), .Y(n_493) );
BUFx4f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx3_ASAP7_75t_L g212 ( .A(n_116), .Y(n_212) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_117), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g179 ( .A(n_117), .B(n_159), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_136), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_120), .A2(n_139), .B1(n_227), .B2(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g491 ( .A(n_120), .Y(n_491) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g524 ( .A(n_121), .Y(n_524) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
OR2x6_ASAP7_75t_L g456 ( .A(n_122), .B(n_143), .Y(n_456) );
INVxp33_ASAP7_75t_L g506 ( .A(n_122), .Y(n_506) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g138 ( .A(n_123), .B(n_125), .Y(n_138) );
AND2x4_ASAP7_75t_L g151 ( .A(n_123), .B(n_133), .Y(n_151) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g525 ( .A(n_126), .Y(n_525) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_L g137 ( .A(n_127), .B(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g143 ( .A(n_128), .Y(n_143) );
AND2x6_ASAP7_75t_L g153 ( .A(n_128), .B(n_131), .Y(n_153) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
INVx1_ASAP7_75t_L g237 ( .A(n_130), .Y(n_237) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g154 ( .A(n_135), .Y(n_154) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_135), .Y(n_483) );
AND2x4_ASAP7_75t_L g139 ( .A(n_138), .B(n_140), .Y(n_139) );
INVxp67_ASAP7_75t_L g489 ( .A(n_139), .Y(n_489) );
NOR2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
INVx1_ASAP7_75t_L g507 ( .A(n_142), .Y(n_507) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g239 ( .A(n_145), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g181 ( .A(n_146), .B(n_171), .Y(n_181) );
OR2x2_ASAP7_75t_L g189 ( .A(n_146), .B(n_190), .Y(n_189) );
AND2x4_ASAP7_75t_L g244 ( .A(n_146), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g291 ( .A(n_146), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_146), .B(n_190), .Y(n_299) );
AND2x2_ASAP7_75t_L g336 ( .A(n_146), .B(n_240), .Y(n_336) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_146), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_146), .B(n_170), .Y(n_377) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_156), .B(n_160), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_155), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_154), .Y(n_149) );
INVxp67_ASAP7_75t_L g462 ( .A(n_151), .Y(n_462) );
INVxp67_ASAP7_75t_L g460 ( .A(n_153), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_154), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_154), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_154), .A2(n_216), .B(n_217), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_154), .B(n_179), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_154), .A2(n_456), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_154), .A2(n_456), .B(n_496), .C(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g503 ( .A(n_154), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_154), .A2(n_456), .B(n_517), .C(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_154), .A2(n_529), .B(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g554 ( .A1(n_154), .A2(n_456), .B(n_555), .C(n_556), .Y(n_554) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_156), .A2(n_163), .B(n_169), .Y(n_162) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_163), .B(n_169), .Y(n_190) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_156), .A2(n_551), .B(n_557), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_157), .A2(n_205), .B(n_209), .Y(n_204) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g278 ( .A(n_161), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_161), .B(n_239), .Y(n_334) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_161), .Y(n_435) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_170), .Y(n_161) );
AND2x2_ASAP7_75t_L g180 ( .A(n_162), .B(n_181), .Y(n_180) );
OR2x2_ASAP7_75t_L g260 ( .A(n_162), .B(n_171), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_162), .B(n_291), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
AND2x2_ASAP7_75t_L g327 ( .A(n_170), .B(n_244), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_170), .B(n_239), .Y(n_383) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g185 ( .A(n_171), .Y(n_185) );
AND2x2_ASAP7_75t_L g254 ( .A(n_171), .B(n_245), .Y(n_254) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
AND2x4_ASAP7_75t_L g281 ( .A(n_171), .B(n_190), .Y(n_281) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_171), .B(n_240), .Y(n_428) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_179), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_179), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_179), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_179), .B(n_233), .Y(n_232) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_179), .B(n_236), .C(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_179), .A2(n_515), .B(n_519), .Y(n_514) );
INVx1_ASAP7_75t_L g407 ( .A(n_180), .Y(n_407) );
INVx1_ASAP7_75t_L g349 ( .A(n_181), .Y(n_349) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_186), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g271 ( .A(n_185), .B(n_189), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_185), .B(n_240), .Y(n_364) );
AND2x2_ASAP7_75t_L g366 ( .A(n_185), .B(n_188), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_185), .A2(n_248), .A3(n_403), .B1(n_433), .B2(n_435), .Y(n_432) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
AND2x2_ASAP7_75t_L g258 ( .A(n_187), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g376 ( .A(n_187), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g399 ( .A(n_187), .B(n_260), .Y(n_399) );
AND2x2_ASAP7_75t_L g426 ( .A(n_187), .B(n_327), .Y(n_426) );
AND2x2_ASAP7_75t_L g352 ( .A(n_188), .B(n_240), .Y(n_352) );
AND2x2_ASAP7_75t_L g427 ( .A(n_188), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g245 ( .A(n_190), .Y(n_245) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NOR2x1p5_ASAP7_75t_L g285 ( .A(n_193), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g303 ( .A(n_193), .Y(n_303) );
OR2x2_ASAP7_75t_L g331 ( .A(n_193), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_SL g248 ( .A(n_194), .B(n_225), .Y(n_248) );
AND2x4_ASAP7_75t_L g264 ( .A(n_194), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g267 ( .A(n_194), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g295 ( .A(n_194), .B(n_204), .Y(n_295) );
OR2x2_ASAP7_75t_L g320 ( .A(n_194), .B(n_269), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_194), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_194), .B(n_204), .Y(n_355) );
INVx2_ASAP7_75t_L g371 ( .A(n_194), .Y(n_371) );
AND2x2_ASAP7_75t_L g386 ( .A(n_194), .B(n_224), .Y(n_386) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_194), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_194), .Y(n_415) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_201), .Y(n_194) );
AND2x2_ASAP7_75t_L g279 ( .A(n_202), .B(n_264), .Y(n_279) );
AND2x2_ASAP7_75t_L g300 ( .A(n_202), .B(n_248), .Y(n_300) );
INVx1_ASAP7_75t_L g332 ( .A(n_202), .Y(n_332) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_210), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g223 ( .A(n_204), .Y(n_223) );
INVx2_ASAP7_75t_L g269 ( .A(n_204), .Y(n_269) );
BUFx3_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
AND2x2_ASAP7_75t_L g325 ( .A(n_204), .B(n_210), .Y(n_325) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_204), .Y(n_423) );
INVx2_ASAP7_75t_L g238 ( .A(n_210), .Y(n_238) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
INVx1_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
OR2x2_ASAP7_75t_L g268 ( .A(n_210), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g288 ( .A(n_210), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_210), .B(n_265), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_210), .B(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_219), .Y(n_211) );
INVx4_ASAP7_75t_L g234 ( .A(n_212), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_212), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_239), .B(n_241), .Y(n_220) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_222), .B(n_224), .Y(n_221) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_222), .Y(n_431) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_SL g257 ( .A(n_223), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_223), .B(n_263), .Y(n_305) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_223), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_224), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g310 ( .A(n_224), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g361 ( .A(n_224), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_224), .A2(n_366), .B1(n_367), .B2(n_372), .C(n_375), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_224), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
INVx3_ASAP7_75t_L g265 ( .A(n_225), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_225), .B(n_269), .Y(n_369) );
AND2x2_ASAP7_75t_L g398 ( .A(n_225), .B(n_371), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_225), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
INVx3_ASAP7_75t_L g468 ( .A(n_234), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_234), .A2(n_468), .B1(n_479), .B2(n_484), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_237), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_237), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g306 ( .A(n_239), .B(n_281), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_239), .A2(n_259), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g243 ( .A(n_240), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
OR2x2_ASAP7_75t_L g298 ( .A(n_240), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_240), .B(n_281), .Y(n_390) );
OR2x2_ASAP7_75t_L g422 ( .A(n_240), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g434 ( .A(n_240), .B(n_340), .Y(n_434) );
INVxp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g312 ( .A(n_243), .Y(n_312) );
INVx3_ASAP7_75t_SL g378 ( .A(n_244), .Y(n_378) );
INVxp67_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AOI322xp5_ASAP7_75t_L g250 ( .A1(n_248), .A2(n_251), .A3(n_255), .B1(n_258), .B2(n_261), .C1(n_266), .C2(n_270), .Y(n_250) );
INVx1_ASAP7_75t_SL g339 ( .A(n_248), .Y(n_339) );
AND2x4_ASAP7_75t_L g424 ( .A(n_248), .B(n_311), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_272), .Y(n_249) );
NOR2x1_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OR2x2_ASAP7_75t_L g277 ( .A(n_252), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g373 ( .A(n_252), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g401 ( .A(n_252), .B(n_254), .Y(n_401) );
AOI32xp33_ASAP7_75t_L g402 ( .A1(n_252), .A2(n_253), .A3(n_403), .B1(n_405), .B2(n_408), .Y(n_402) );
OR2x2_ASAP7_75t_L g406 ( .A(n_252), .B(n_299), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_253), .B(n_278), .C(n_363), .Y(n_362) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_253), .A2(n_319), .B1(n_383), .B2(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g385 ( .A(n_256), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_260), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OAI322xp33_ASAP7_75t_L g308 ( .A1(n_264), .A2(n_268), .A3(n_277), .B1(n_309), .B2(n_312), .C1(n_313), .C2(n_314), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_264), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_264), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g287 ( .A(n_265), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g319 ( .A(n_265), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_265), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g380 ( .A(n_268), .Y(n_380) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_269), .Y(n_311) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_279), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_275), .B(n_323), .Y(n_322) );
AOI322xp5_ASAP7_75t_SL g417 ( .A1(n_275), .A2(n_281), .A3(n_398), .B1(n_416), .B2(n_418), .C1(n_421), .C2(n_424), .Y(n_417) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_296), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_281), .B(n_291), .Y(n_313) );
INVx2_ASAP7_75t_SL g323 ( .A(n_281), .Y(n_323) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g348 ( .A(n_287), .Y(n_348) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g393 ( .A(n_294), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g347 ( .A(n_295), .B(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_301), .B2(n_306), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR4xp75_ASAP7_75t_L g307 ( .A(n_308), .B(n_321), .C(n_341), .D(n_357), .Y(n_307) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_319), .A2(n_396), .B1(n_399), .B2(n_400), .Y(n_395) );
OR2x2_ASAP7_75t_L g360 ( .A(n_320), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g404 ( .A(n_320), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B1(n_326), .B2(n_328), .C(n_329), .Y(n_321) );
INVx2_ASAP7_75t_L g340 ( .A(n_325), .Y(n_340) );
AND2x2_ASAP7_75t_L g397 ( .A(n_325), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_335), .B2(n_337), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_343), .B1(n_359), .B2(n_362), .Y(n_358) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_830), .Y(n_341) );
AND2x2_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g409 ( .A(n_348), .B(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_365), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_379), .Y(n_375) );
NOR3xp33_ASAP7_75t_SL g381 ( .A(n_382), .B(n_387), .C(n_411), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_402), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_393), .C(n_395), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g403 ( .A(n_394), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NAND4xp25_ASAP7_75t_SL g411 ( .A(n_412), .B(n_417), .C(n_425), .D(n_432), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_427), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_436), .Y(n_793) );
OR2x6_ASAP7_75t_SL g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x6_ASAP7_75t_SL g788 ( .A(n_437), .B(n_439), .Y(n_788) );
OR2x2_ASAP7_75t_L g797 ( .A(n_437), .B(n_439), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_437), .B(n_438), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI211x1_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_641), .B(n_642), .C(n_782), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND4x1_ASAP7_75t_L g782 ( .A(n_446), .B(n_643), .C(n_783), .D(n_784), .Y(n_782) );
NAND3x1_ASAP7_75t_L g813 ( .A(n_446), .B(n_643), .C(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_609), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_532), .B(n_544), .C(n_585), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_464), .B(n_510), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_450), .A2(n_533), .B(n_538), .C(n_543), .Y(n_532) );
NAND2x1_ASAP7_75t_L g662 ( .A(n_450), .B(n_663), .Y(n_662) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_450), .B(n_682), .Y(n_753) );
AND2x2_ASAP7_75t_L g772 ( .A(n_450), .B(n_512), .Y(n_772) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g549 ( .A(n_451), .Y(n_549) );
AND2x2_ASAP7_75t_L g620 ( .A(n_451), .B(n_550), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_451), .B(n_521), .Y(n_625) );
NOR2x1_ASAP7_75t_SL g741 ( .A(n_451), .B(n_512), .Y(n_741) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_458), .B(n_463), .Y(n_453) );
INVxp67_ASAP7_75t_L g480 ( .A(n_456), .Y(n_480) );
INVx2_ASAP7_75t_L g531 ( .A(n_456), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_458) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_492), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_466), .B(n_590), .Y(n_656) );
AND2x2_ASAP7_75t_L g773 ( .A(n_466), .B(n_614), .Y(n_773) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_467), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g562 ( .A(n_467), .Y(n_562) );
AND2x2_ASAP7_75t_L g570 ( .A(n_467), .B(n_571), .Y(n_570) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_467), .B(n_476), .Y(n_708) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_475), .Y(n_467) );
AO21x2_ASAP7_75t_L g593 ( .A1(n_468), .A2(n_469), .B(n_475), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g660 ( .A(n_476), .B(n_500), .Y(n_660) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g536 ( .A(n_477), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
INVx1_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_477), .B(n_593), .Y(n_617) );
AND2x2_ASAP7_75t_L g666 ( .A(n_477), .B(n_493), .Y(n_666) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g621 ( .A(n_492), .B(n_616), .Y(n_621) );
AND2x2_ASAP7_75t_L g677 ( .A(n_492), .B(n_560), .Y(n_677) );
AND2x2_ASAP7_75t_L g692 ( .A(n_492), .B(n_606), .Y(n_692) );
AND2x2_ASAP7_75t_L g729 ( .A(n_492), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g745 ( .A(n_492), .Y(n_745) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
INVx1_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_493), .B(n_572), .Y(n_575) );
INVx1_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
INVxp67_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g534 ( .A(n_500), .Y(n_534) );
AND2x4_ASAP7_75t_L g561 ( .A(n_500), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_502), .B(n_508), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g543 ( .A(n_510), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_510), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_511), .B(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_511), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_511), .B(n_578), .Y(n_721) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_511), .Y(n_759) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
INVx2_ASAP7_75t_L g584 ( .A(n_512), .Y(n_584) );
AND2x2_ASAP7_75t_L g595 ( .A(n_512), .B(n_521), .Y(n_595) );
INVx4_ASAP7_75t_L g603 ( .A(n_512), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_512), .B(n_579), .Y(n_639) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_512), .Y(n_652) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x4_ASAP7_75t_L g630 ( .A(n_520), .B(n_603), .Y(n_630) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g581 ( .A(n_521), .B(n_549), .Y(n_581) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_521), .Y(n_602) );
INVx2_ASAP7_75t_L g651 ( .A(n_521), .Y(n_651) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .C(n_526), .Y(n_523) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_534), .B(n_539), .Y(n_640) );
NAND2x1_ASAP7_75t_SL g754 ( .A(n_534), .B(n_536), .Y(n_754) );
OR2x2_ASAP7_75t_L g633 ( .A(n_535), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g736 ( .A(n_535), .Y(n_736) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g626 ( .A(n_536), .B(n_561), .Y(n_626) );
AND2x2_ASAP7_75t_L g742 ( .A(n_536), .B(n_735), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_538), .A2(n_751), .B1(n_754), .B2(n_755), .C(n_757), .Y(n_750) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_539), .A2(n_695), .B1(n_697), .B2(n_699), .Y(n_694) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_540), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g608 ( .A(n_540), .Y(n_608) );
BUFx2_ASAP7_75t_L g689 ( .A(n_540), .Y(n_689) );
AND2x2_ASAP7_75t_L g659 ( .A(n_541), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_563), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g632 ( .A(n_548), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_548), .B(n_758), .C(n_759), .D(n_760), .Y(n_757) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g567 ( .A(n_549), .Y(n_567) );
AND2x2_ASAP7_75t_L g650 ( .A(n_549), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g566 ( .A(n_550), .Y(n_566) );
INVx2_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_550), .Y(n_607) );
INVx1_ASAP7_75t_L g624 ( .A(n_550), .Y(n_624) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_550), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g771 ( .A(n_559), .Y(n_771) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g569 ( .A(n_560), .Y(n_569) );
AND2x2_ASAP7_75t_L g665 ( .A(n_561), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g765 ( .A(n_561), .B(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_568), .B1(n_573), .B2(n_576), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_565), .B(n_630), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_565), .B(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g746 ( .A(n_565), .B(n_724), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_565), .A2(n_601), .B(n_723), .Y(n_776) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_566), .B(n_650), .Y(n_687) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_566), .Y(n_703) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g573 ( .A(n_569), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g590 ( .A(n_571), .Y(n_590) );
AND2x2_ASAP7_75t_L g614 ( .A(n_571), .B(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g735 ( .A(n_571), .B(n_592), .Y(n_735) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_572), .B(n_593), .Y(n_634) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g710 ( .A(n_575), .B(n_617), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g691 ( .A(n_577), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_578), .B(n_587), .C(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g658 ( .A(n_578), .B(n_601), .Y(n_658) );
AND2x2_ASAP7_75t_L g740 ( .A(n_578), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g766 ( .A(n_578), .Y(n_766) );
INVx1_ASAP7_75t_L g780 ( .A(n_578), .Y(n_780) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g583 ( .A(n_581), .B(n_584), .Y(n_583) );
INVx4_ASAP7_75t_L g739 ( .A(n_581), .Y(n_739) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g779 ( .A(n_583), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g682 ( .A(n_584), .Y(n_682) );
AO22x1_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_594), .B1(n_596), .B2(n_604), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_588), .B(n_592), .Y(n_672) );
INVx3_ASAP7_75t_L g706 ( .A(n_588), .Y(n_706) );
BUFx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g606 ( .A(n_592), .Y(n_606) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g684 ( .A(n_593), .B(n_599), .Y(n_684) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_593), .Y(n_731) );
AOI31xp33_ASAP7_75t_L g635 ( .A1(n_594), .A2(n_636), .A3(n_638), .B(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_595), .A2(n_612), .B1(n_618), .B2(n_621), .Y(n_611) );
AND2x2_ASAP7_75t_L g695 ( .A(n_595), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g702 ( .A(n_595), .B(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_601), .B(n_756), .Y(n_755) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OR2x2_ASAP7_75t_L g631 ( .A(n_603), .B(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_603), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g726 ( .A(n_606), .B(n_666), .Y(n_726) );
INVx1_ASAP7_75t_L g761 ( .A(n_606), .Y(n_761) );
AND2x2_ASAP7_75t_L g711 ( .A(n_607), .B(n_650), .Y(n_711) );
BUFx2_ASAP7_75t_L g756 ( .A(n_607), .Y(n_756) );
AND2x2_ASAP7_75t_L g699 ( .A(n_608), .B(n_700), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_627), .C(n_635), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_622), .Y(n_610) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AND2x2_ASAP7_75t_L g688 ( .A(n_614), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_620), .B(n_630), .Y(n_653) );
AND2x2_ASAP7_75t_L g675 ( .A(n_620), .B(n_652), .Y(n_675) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_620), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
AND2x2_ASAP7_75t_L g778 ( .A(n_623), .B(n_652), .Y(n_778) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g752 ( .A(n_624), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g669 ( .A(n_625), .Y(n_669) );
AND2x2_ASAP7_75t_L g769 ( .A(n_625), .B(n_652), .Y(n_769) );
AOI21xp33_ASAP7_75t_R g627 ( .A1(n_628), .A2(n_631), .B(n_633), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_629), .B(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_630), .Y(n_637) );
INVx1_ASAP7_75t_L g700 ( .A(n_634), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_636), .A2(n_654), .B1(n_668), .B2(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g668 ( .A(n_639), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_641), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_641), .B(n_748), .Y(n_747) );
NOR2xp67_ASAP7_75t_SL g783 ( .A(n_641), .B(n_714), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_712), .B(n_713), .C(n_747), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_678), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_667), .C(n_673), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_654), .B(n_657), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_653), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_649), .A2(n_688), .B1(n_691), .B2(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g725 ( .A(n_651), .Y(n_725) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g717 ( .A(n_656), .B(n_706), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_661), .B2(n_665), .Y(n_657) );
INVx1_ASAP7_75t_L g671 ( .A(n_660), .Y(n_671) );
AND2x4_ASAP7_75t_L g683 ( .A(n_660), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g719 ( .A(n_662), .Y(n_719) );
INVx1_ASAP7_75t_L g696 ( .A(n_663), .Y(n_696) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_665), .A2(n_675), .B1(n_723), .B2(n_726), .Y(n_722) );
INVxp67_ASAP7_75t_L g767 ( .A(n_666), .Y(n_767) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_669), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVxp33_ASAP7_75t_L g781 ( .A(n_672), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_693), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_680), .B(n_690), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_685), .B2(n_688), .Y(n_680) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_701), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_709), .B2(n_711), .Y(n_701) );
NOR2xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g758 ( .A(n_706), .Y(n_758) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g814 ( .A(n_715), .B(n_749), .Y(n_814) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_727), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_722), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND4xp25_ASAP7_75t_SL g727 ( .A(n_728), .B(n_732), .C(n_737), .D(n_743), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g770 ( .A(n_735), .B(n_771), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B(n_742), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g784 ( .A(n_748), .Y(n_784) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR3x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_762), .C(n_774), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_767), .B(n_768), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_768) );
INVx1_ASAP7_75t_L g775 ( .A(n_773), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_777), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B(n_781), .Y(n_777) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx6p67_ASAP7_75t_R g791 ( .A(n_786), .Y(n_791) );
INVx3_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_800), .A2(n_810), .B(n_819), .Y(n_809) );
NOR2xp33_ASAP7_75t_SL g800 ( .A(n_801), .B(n_803), .Y(n_800) );
INVx1_ASAP7_75t_SL g820 ( .A(n_801), .Y(n_820) );
BUFx2_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
CKINVDCx8_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
OAI22xp5_ASAP7_75t_SL g810 ( .A1(n_811), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_813), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_815), .Y(n_818) );
INVx1_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_SL g828 ( .A(n_821), .Y(n_828) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_SL g823 ( .A(n_824), .B(n_825), .Y(n_823) );
endmodule