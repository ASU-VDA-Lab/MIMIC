module real_jpeg_31188_n_8 (n_5, n_4, n_68, n_0, n_70, n_1, n_2, n_71, n_66, n_6, n_72, n_7, n_3, n_69, n_67, n_8);

input n_5;
input n_4;
input n_68;
input n_0;
input n_70;
input n_1;
input n_2;
input n_71;
input n_66;
input n_6;
input n_72;
input n_7;
input n_3;
input n_69;
input n_67;

output n_8;

wire n_17;
wire n_57;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

AOI221xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_3),
.B1(n_30),
.B2(n_34),
.C(n_36),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_30),
.C(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g9 ( 
.A(n_5),
.B(n_10),
.CON(n_9),
.SN(n_9)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_16),
.Y(n_8)
);

BUFx24_ASAP7_75t_SL g64 ( 
.A(n_9),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_55),
.B(n_62),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.C(n_51),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_40),
.B(n_49),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_69),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_66),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_67),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_68),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_70),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_71),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_72),
.Y(n_58)
);


endmodule